module pci_bridge32_slow (
ispd_clk,
pci_ad_i_0_,
pci_ad_i_10_,
pci_ad_i_11_,
pci_ad_i_12_,
pci_ad_i_13_,
pci_ad_i_14_,
pci_ad_i_15_,
pci_ad_i_16_,
pci_ad_i_17_,
pci_ad_i_18_,
pci_ad_i_19_,
pci_ad_i_1_,
pci_ad_i_20_,
pci_ad_i_21_,
pci_ad_i_22_,
pci_ad_i_23_,
pci_ad_i_24_,
pci_ad_i_25_,
pci_ad_i_26_,
pci_ad_i_27_,
pci_ad_i_28_,
pci_ad_i_29_,
pci_ad_i_2_,
pci_ad_i_30_,
pci_ad_i_31_,
pci_ad_i_3_,
pci_ad_i_4_,
pci_ad_i_5_,
pci_ad_i_6_,
pci_ad_i_7_,
pci_ad_i_8_,
pci_ad_i_9_,
pci_cbe_i_0_,
pci_cbe_i_1_,
pci_cbe_i_2_,
pci_cbe_i_3_,
pci_devsel_i,
pci_frame_i,
pci_gnt_i,
pci_idsel_i,
pci_irdy_i,
pci_par_i,
pci_perr_i,
pci_rst_i,
pci_rst_oe_o,
pci_stop_i,
pci_trdy_i,
wb_int_i,
wbm_ack_i,
wbm_dat_i_0_,
wbm_dat_i_10_,
wbm_dat_i_11_,
wbm_dat_i_12_,
wbm_dat_i_13_,
wbm_dat_i_14_,
wbm_dat_i_15_,
wbm_dat_i_16_,
wbm_dat_i_17_,
wbm_dat_i_18_,
wbm_dat_i_19_,
wbm_dat_i_1_,
wbm_dat_i_20_,
wbm_dat_i_21_,
wbm_dat_i_22_,
wbm_dat_i_23_,
wbm_dat_i_24_,
wbm_dat_i_25_,
wbm_dat_i_26_,
wbm_dat_i_27_,
wbm_dat_i_28_,
wbm_dat_i_29_,
wbm_dat_i_2_,
wbm_dat_i_30_,
wbm_dat_i_31_,
wbm_dat_i_3_,
wbm_dat_i_4_,
wbm_dat_i_5_,
wbm_dat_i_6_,
wbm_dat_i_7_,
wbm_dat_i_8_,
wbm_dat_i_9_,
wbm_err_i,
wbm_rty_i,
wbs_adr_i_0_,
wbs_adr_i_10_,
wbs_adr_i_11_,
wbs_adr_i_12_,
wbs_adr_i_13_,
wbs_adr_i_14_,
wbs_adr_i_15_,
wbs_adr_i_16_,
wbs_adr_i_17_,
wbs_adr_i_18_,
wbs_adr_i_19_,
wbs_adr_i_1_,
wbs_adr_i_20_,
wbs_adr_i_21_,
wbs_adr_i_22_,
wbs_adr_i_23_,
wbs_adr_i_24_,
wbs_adr_i_25_,
wbs_adr_i_26_,
wbs_adr_i_27_,
wbs_adr_i_28_,
wbs_adr_i_29_,
wbs_adr_i_2_,
wbs_adr_i_30_,
wbs_adr_i_31_,
wbs_adr_i_3_,
wbs_adr_i_4_,
wbs_adr_i_5_,
wbs_adr_i_6_,
wbs_adr_i_7_,
wbs_adr_i_8_,
wbs_adr_i_9_,
wbs_bte_i_0_,
wbs_bte_i_1_,
wbs_cti_i_0_,
wbs_cti_i_1_,
wbs_cti_i_2_,
wbs_cyc_i,
wbs_dat_i_0_,
wbs_dat_i_10_,
wbs_dat_i_11_,
wbs_dat_i_12_,
wbs_dat_i_13_,
wbs_dat_i_14_,
wbs_dat_i_15_,
wbs_dat_i_16_,
wbs_dat_i_17_,
wbs_dat_i_18_,
wbs_dat_i_19_,
wbs_dat_i_1_,
wbs_dat_i_20_,
wbs_dat_i_21_,
wbs_dat_i_22_,
wbs_dat_i_23_,
wbs_dat_i_24_,
wbs_dat_i_25_,
wbs_dat_i_26_,
wbs_dat_i_27_,
wbs_dat_i_28_,
wbs_dat_i_29_,
wbs_dat_i_2_,
wbs_dat_i_30_,
wbs_dat_i_31_,
wbs_dat_i_3_,
wbs_dat_i_4_,
wbs_dat_i_5_,
wbs_dat_i_6_,
wbs_dat_i_7_,
wbs_dat_i_8_,
wbs_dat_i_9_,
wbs_sel_i_0_,
wbs_sel_i_1_,
wbs_sel_i_2_,
wbs_sel_i_3_,
wbs_stb_i,
wbs_we_i,
pci_ad_o_0_,
pci_ad_o_10_,
pci_ad_o_11_,
pci_ad_o_12_,
pci_ad_o_13_,
pci_ad_o_14_,
pci_ad_o_15_,
pci_ad_o_16_,
pci_ad_o_17_,
pci_ad_o_18_,
pci_ad_o_19_,
pci_ad_o_1_,
pci_ad_o_20_,
pci_ad_o_21_,
pci_ad_o_22_,
pci_ad_o_23_,
pci_ad_o_24_,
pci_ad_o_25_,
pci_ad_o_26_,
pci_ad_o_27_,
pci_ad_o_28_,
pci_ad_o_29_,
pci_ad_o_2_,
pci_ad_o_30_,
pci_ad_o_31_,
pci_ad_o_3_,
pci_ad_o_4_,
pci_ad_o_5_,
pci_ad_o_6_,
pci_ad_o_7_,
pci_ad_o_8_,
pci_ad_o_9_,
pci_ad_oe_o_0_,
pci_ad_oe_o_10_,
pci_ad_oe_o_11_,
pci_ad_oe_o_12_,
pci_ad_oe_o_13_,
pci_ad_oe_o_14_,
pci_ad_oe_o_15_,
pci_ad_oe_o_16_,
pci_ad_oe_o_17_,
pci_ad_oe_o_18_,
pci_ad_oe_o_19_,
pci_ad_oe_o_1_,
pci_ad_oe_o_20_,
pci_ad_oe_o_21_,
pci_ad_oe_o_22_,
pci_ad_oe_o_23_,
pci_ad_oe_o_24_,
pci_ad_oe_o_25_,
pci_ad_oe_o_26_,
pci_ad_oe_o_27_,
pci_ad_oe_o_28_,
pci_ad_oe_o_29_,
pci_ad_oe_o_2_,
pci_ad_oe_o_30_,
pci_ad_oe_o_31_,
pci_ad_oe_o_3_,
pci_ad_oe_o_4_,
pci_ad_oe_o_5_,
pci_ad_oe_o_6_,
pci_ad_oe_o_7_,
pci_ad_oe_o_8_,
pci_ad_oe_o_9_,
pci_cbe_o_0_,
pci_cbe_o_1_,
pci_cbe_o_2_,
pci_cbe_o_3_,
pci_cbe_oe_o_0_,
pci_cbe_oe_o_1_,
pci_cbe_oe_o_2_,
pci_cbe_oe_o_3_,
pci_devsel_o,
pci_devsel_oe_o,
pci_frame_o,
pci_frame_oe_o,
pci_inta_oe_o,
pci_irdy_o,
pci_irdy_oe_o,
pci_par_o,
pci_par_oe_o,
pci_perr_o,
pci_perr_oe_o,
pci_req_o,
pci_req_oe_o,
pci_serr_o,
pci_serr_oe_o,
pci_stop_o,
pci_stop_oe_o,
pci_trdy_o,
pci_trdy_oe_o,
wb_rst_o,
wbm_adr_o_0_,
wbm_adr_o_10_,
wbm_adr_o_11_,
wbm_adr_o_12_,
wbm_adr_o_13_,
wbm_adr_o_14_,
wbm_adr_o_15_,
wbm_adr_o_16_,
wbm_adr_o_17_,
wbm_adr_o_18_,
wbm_adr_o_19_,
wbm_adr_o_1_,
wbm_adr_o_20_,
wbm_adr_o_21_,
wbm_adr_o_22_,
wbm_adr_o_23_,
wbm_adr_o_24_,
wbm_adr_o_25_,
wbm_adr_o_26_,
wbm_adr_o_27_,
wbm_adr_o_28_,
wbm_adr_o_29_,
wbm_adr_o_2_,
wbm_adr_o_30_,
wbm_adr_o_31_,
wbm_adr_o_3_,
wbm_adr_o_4_,
wbm_adr_o_5_,
wbm_adr_o_6_,
wbm_adr_o_7_,
wbm_adr_o_8_,
wbm_adr_o_9_,
wbm_cti_o_0_,
wbm_cti_o_1_,
wbm_cti_o_2_,
wbm_cyc_o,
wbm_dat_o_0_,
wbm_dat_o_10_,
wbm_dat_o_11_,
wbm_dat_o_12_,
wbm_dat_o_13_,
wbm_dat_o_14_,
wbm_dat_o_15_,
wbm_dat_o_16_,
wbm_dat_o_17_,
wbm_dat_o_18_,
wbm_dat_o_19_,
wbm_dat_o_1_,
wbm_dat_o_20_,
wbm_dat_o_21_,
wbm_dat_o_22_,
wbm_dat_o_23_,
wbm_dat_o_24_,
wbm_dat_o_25_,
wbm_dat_o_26_,
wbm_dat_o_27_,
wbm_dat_o_28_,
wbm_dat_o_29_,
wbm_dat_o_2_,
wbm_dat_o_30_,
wbm_dat_o_31_,
wbm_dat_o_3_,
wbm_dat_o_4_,
wbm_dat_o_5_,
wbm_dat_o_6_,
wbm_dat_o_7_,
wbm_dat_o_8_,
wbm_dat_o_9_,
wbm_sel_o_0_,
wbm_sel_o_1_,
wbm_sel_o_2_,
wbm_sel_o_3_,
wbm_stb_o,
wbm_we_o,
wbs_ack_o,
wbs_dat_o_0_,
wbs_dat_o_10_,
wbs_dat_o_11_,
wbs_dat_o_12_,
wbs_dat_o_13_,
wbs_dat_o_14_,
wbs_dat_o_15_,
wbs_dat_o_16_,
wbs_dat_o_17_,
wbs_dat_o_18_,
wbs_dat_o_19_,
wbs_dat_o_1_,
wbs_dat_o_20_,
wbs_dat_o_21_,
wbs_dat_o_22_,
wbs_dat_o_23_,
wbs_dat_o_24_,
wbs_dat_o_25_,
wbs_dat_o_26_,
wbs_dat_o_27_,
wbs_dat_o_28_,
wbs_dat_o_29_,
wbs_dat_o_2_,
wbs_dat_o_30_,
wbs_dat_o_31_,
wbs_dat_o_3_,
wbs_dat_o_4_,
wbs_dat_o_5_,
wbs_dat_o_6_,
wbs_dat_o_7_,
wbs_dat_o_8_,
wbs_dat_o_9_,
wbs_err_o,
wbs_rty_o
);

// Start PIs
input ispd_clk;
input pci_ad_i_0_;
input pci_ad_i_10_;
input pci_ad_i_11_;
input pci_ad_i_12_;
input pci_ad_i_13_;
input pci_ad_i_14_;
input pci_ad_i_15_;
input pci_ad_i_16_;
input pci_ad_i_17_;
input pci_ad_i_18_;
input pci_ad_i_19_;
input pci_ad_i_1_;
input pci_ad_i_20_;
input pci_ad_i_21_;
input pci_ad_i_22_;
input pci_ad_i_23_;
input pci_ad_i_24_;
input pci_ad_i_25_;
input pci_ad_i_26_;
input pci_ad_i_27_;
input pci_ad_i_28_;
input pci_ad_i_29_;
input pci_ad_i_2_;
input pci_ad_i_30_;
input pci_ad_i_31_;
input pci_ad_i_3_;
input pci_ad_i_4_;
input pci_ad_i_5_;
input pci_ad_i_6_;
input pci_ad_i_7_;
input pci_ad_i_8_;
input pci_ad_i_9_;
input pci_cbe_i_0_;
input pci_cbe_i_1_;
input pci_cbe_i_2_;
input pci_cbe_i_3_;
input pci_devsel_i;
input pci_frame_i;
input pci_gnt_i;
input pci_idsel_i;
input pci_irdy_i;
input pci_par_i;
input pci_perr_i;
input pci_rst_i;
input pci_rst_oe_o;
input pci_stop_i;
input pci_trdy_i;
input wb_int_i;
input wbm_ack_i;
input wbm_dat_i_0_;
input wbm_dat_i_10_;
input wbm_dat_i_11_;
input wbm_dat_i_12_;
input wbm_dat_i_13_;
input wbm_dat_i_14_;
input wbm_dat_i_15_;
input wbm_dat_i_16_;
input wbm_dat_i_17_;
input wbm_dat_i_18_;
input wbm_dat_i_19_;
input wbm_dat_i_1_;
input wbm_dat_i_20_;
input wbm_dat_i_21_;
input wbm_dat_i_22_;
input wbm_dat_i_23_;
input wbm_dat_i_24_;
input wbm_dat_i_25_;
input wbm_dat_i_26_;
input wbm_dat_i_27_;
input wbm_dat_i_28_;
input wbm_dat_i_29_;
input wbm_dat_i_2_;
input wbm_dat_i_30_;
input wbm_dat_i_31_;
input wbm_dat_i_3_;
input wbm_dat_i_4_;
input wbm_dat_i_5_;
input wbm_dat_i_6_;
input wbm_dat_i_7_;
input wbm_dat_i_8_;
input wbm_dat_i_9_;
input wbm_err_i;
input wbm_rty_i;
input wbs_adr_i_0_;
input wbs_adr_i_10_;
input wbs_adr_i_11_;
input wbs_adr_i_12_;
input wbs_adr_i_13_;
input wbs_adr_i_14_;
input wbs_adr_i_15_;
input wbs_adr_i_16_;
input wbs_adr_i_17_;
input wbs_adr_i_18_;
input wbs_adr_i_19_;
input wbs_adr_i_1_;
input wbs_adr_i_20_;
input wbs_adr_i_21_;
input wbs_adr_i_22_;
input wbs_adr_i_23_;
input wbs_adr_i_24_;
input wbs_adr_i_25_;
input wbs_adr_i_26_;
input wbs_adr_i_27_;
input wbs_adr_i_28_;
input wbs_adr_i_29_;
input wbs_adr_i_2_;
input wbs_adr_i_30_;
input wbs_adr_i_31_;
input wbs_adr_i_3_;
input wbs_adr_i_4_;
input wbs_adr_i_5_;
input wbs_adr_i_6_;
input wbs_adr_i_7_;
input wbs_adr_i_8_;
input wbs_adr_i_9_;
input wbs_bte_i_0_;
input wbs_bte_i_1_;
input wbs_cti_i_0_;
input wbs_cti_i_1_;
input wbs_cti_i_2_;
input wbs_cyc_i;
input wbs_dat_i_0_;
input wbs_dat_i_10_;
input wbs_dat_i_11_;
input wbs_dat_i_12_;
input wbs_dat_i_13_;
input wbs_dat_i_14_;
input wbs_dat_i_15_;
input wbs_dat_i_16_;
input wbs_dat_i_17_;
input wbs_dat_i_18_;
input wbs_dat_i_19_;
input wbs_dat_i_1_;
input wbs_dat_i_20_;
input wbs_dat_i_21_;
input wbs_dat_i_22_;
input wbs_dat_i_23_;
input wbs_dat_i_24_;
input wbs_dat_i_25_;
input wbs_dat_i_26_;
input wbs_dat_i_27_;
input wbs_dat_i_28_;
input wbs_dat_i_29_;
input wbs_dat_i_2_;
input wbs_dat_i_30_;
input wbs_dat_i_31_;
input wbs_dat_i_3_;
input wbs_dat_i_4_;
input wbs_dat_i_5_;
input wbs_dat_i_6_;
input wbs_dat_i_7_;
input wbs_dat_i_8_;
input wbs_dat_i_9_;
input wbs_sel_i_0_;
input wbs_sel_i_1_;
input wbs_sel_i_2_;
input wbs_sel_i_3_;
input wbs_stb_i;
input wbs_we_i;

// Start POs
output pci_ad_o_0_;
output pci_ad_o_10_;
output pci_ad_o_11_;
output pci_ad_o_12_;
output pci_ad_o_13_;
output pci_ad_o_14_;
output pci_ad_o_15_;
output pci_ad_o_16_;
output pci_ad_o_17_;
output pci_ad_o_18_;
output pci_ad_o_19_;
output pci_ad_o_1_;
output pci_ad_o_20_;
output pci_ad_o_21_;
output pci_ad_o_22_;
output pci_ad_o_23_;
output pci_ad_o_24_;
output pci_ad_o_25_;
output pci_ad_o_26_;
output pci_ad_o_27_;
output pci_ad_o_28_;
output pci_ad_o_29_;
output pci_ad_o_2_;
output pci_ad_o_30_;
output pci_ad_o_31_;
output pci_ad_o_3_;
output pci_ad_o_4_;
output pci_ad_o_5_;
output pci_ad_o_6_;
output pci_ad_o_7_;
output pci_ad_o_8_;
output pci_ad_o_9_;
output pci_ad_oe_o_0_;
output pci_ad_oe_o_10_;
output pci_ad_oe_o_11_;
output pci_ad_oe_o_12_;
output pci_ad_oe_o_13_;
output pci_ad_oe_o_14_;
output pci_ad_oe_o_15_;
output pci_ad_oe_o_16_;
output pci_ad_oe_o_17_;
output pci_ad_oe_o_18_;
output pci_ad_oe_o_19_;
output pci_ad_oe_o_1_;
output pci_ad_oe_o_20_;
output pci_ad_oe_o_21_;
output pci_ad_oe_o_22_;
output pci_ad_oe_o_23_;
output pci_ad_oe_o_24_;
output pci_ad_oe_o_25_;
output pci_ad_oe_o_26_;
output pci_ad_oe_o_27_;
output pci_ad_oe_o_28_;
output pci_ad_oe_o_29_;
output pci_ad_oe_o_2_;
output pci_ad_oe_o_30_;
output pci_ad_oe_o_31_;
output pci_ad_oe_o_3_;
output pci_ad_oe_o_4_;
output pci_ad_oe_o_5_;
output pci_ad_oe_o_6_;
output pci_ad_oe_o_7_;
output pci_ad_oe_o_8_;
output pci_ad_oe_o_9_;
output pci_cbe_o_0_;
output pci_cbe_o_1_;
output pci_cbe_o_2_;
output pci_cbe_o_3_;
output pci_cbe_oe_o_0_;
output pci_cbe_oe_o_1_;
output pci_cbe_oe_o_2_;
output pci_cbe_oe_o_3_;
output pci_devsel_o;
output pci_devsel_oe_o;
output pci_frame_o;
output pci_frame_oe_o;
output pci_inta_oe_o;
output pci_irdy_o;
output pci_irdy_oe_o;
output pci_par_o;
output pci_par_oe_o;
output pci_perr_o;
output pci_perr_oe_o;
output pci_req_o;
output pci_req_oe_o;
output pci_serr_o;
output pci_serr_oe_o;
output pci_stop_o;
output pci_stop_oe_o;
output pci_trdy_o;
output pci_trdy_oe_o;
output wb_rst_o;
output wbm_adr_o_0_;
output wbm_adr_o_10_;
output wbm_adr_o_11_;
output wbm_adr_o_12_;
output wbm_adr_o_13_;
output wbm_adr_o_14_;
output wbm_adr_o_15_;
output wbm_adr_o_16_;
output wbm_adr_o_17_;
output wbm_adr_o_18_;
output wbm_adr_o_19_;
output wbm_adr_o_1_;
output wbm_adr_o_20_;
output wbm_adr_o_21_;
output wbm_adr_o_22_;
output wbm_adr_o_23_;
output wbm_adr_o_24_;
output wbm_adr_o_25_;
output wbm_adr_o_26_;
output wbm_adr_o_27_;
output wbm_adr_o_28_;
output wbm_adr_o_29_;
output wbm_adr_o_2_;
output wbm_adr_o_30_;
output wbm_adr_o_31_;
output wbm_adr_o_3_;
output wbm_adr_o_4_;
output wbm_adr_o_5_;
output wbm_adr_o_6_;
output wbm_adr_o_7_;
output wbm_adr_o_8_;
output wbm_adr_o_9_;
output wbm_cti_o_0_;
output wbm_cti_o_1_;
output wbm_cti_o_2_;
output wbm_cyc_o;
output wbm_dat_o_0_;
output wbm_dat_o_10_;
output wbm_dat_o_11_;
output wbm_dat_o_12_;
output wbm_dat_o_13_;
output wbm_dat_o_14_;
output wbm_dat_o_15_;
output wbm_dat_o_16_;
output wbm_dat_o_17_;
output wbm_dat_o_18_;
output wbm_dat_o_19_;
output wbm_dat_o_1_;
output wbm_dat_o_20_;
output wbm_dat_o_21_;
output wbm_dat_o_22_;
output wbm_dat_o_23_;
output wbm_dat_o_24_;
output wbm_dat_o_25_;
output wbm_dat_o_26_;
output wbm_dat_o_27_;
output wbm_dat_o_28_;
output wbm_dat_o_29_;
output wbm_dat_o_2_;
output wbm_dat_o_30_;
output wbm_dat_o_31_;
output wbm_dat_o_3_;
output wbm_dat_o_4_;
output wbm_dat_o_5_;
output wbm_dat_o_6_;
output wbm_dat_o_7_;
output wbm_dat_o_8_;
output wbm_dat_o_9_;
output wbm_sel_o_0_;
output wbm_sel_o_1_;
output wbm_sel_o_2_;
output wbm_sel_o_3_;
output wbm_stb_o;
output wbm_we_o;
output wbs_ack_o;
output wbs_dat_o_0_;
output wbs_dat_o_10_;
output wbs_dat_o_11_;
output wbs_dat_o_12_;
output wbs_dat_o_13_;
output wbs_dat_o_14_;
output wbs_dat_o_15_;
output wbs_dat_o_16_;
output wbs_dat_o_17_;
output wbs_dat_o_18_;
output wbs_dat_o_19_;
output wbs_dat_o_1_;
output wbs_dat_o_20_;
output wbs_dat_o_21_;
output wbs_dat_o_22_;
output wbs_dat_o_23_;
output wbs_dat_o_24_;
output wbs_dat_o_25_;
output wbs_dat_o_26_;
output wbs_dat_o_27_;
output wbs_dat_o_28_;
output wbs_dat_o_29_;
output wbs_dat_o_2_;
output wbs_dat_o_30_;
output wbs_dat_o_31_;
output wbs_dat_o_3_;
output wbs_dat_o_4_;
output wbs_dat_o_5_;
output wbs_dat_o_6_;
output wbs_dat_o_7_;
output wbs_dat_o_8_;
output wbs_dat_o_9_;
output wbs_err_o;
output wbs_rty_o;

// Start wires
wire ispd_clk;
wire pci_ad_i_0_;
wire pci_ad_i_10_;
wire pci_ad_i_11_;
wire pci_ad_i_12_;
wire pci_ad_i_13_;
wire pci_ad_i_14_;
wire pci_ad_i_15_;
wire pci_ad_i_16_;
wire pci_ad_i_17_;
wire pci_ad_i_18_;
wire pci_ad_i_19_;
wire pci_ad_i_1_;
wire pci_ad_i_20_;
wire pci_ad_i_21_;
wire pci_ad_i_22_;
wire pci_ad_i_23_;
wire pci_ad_i_24_;
wire pci_ad_i_25_;
wire pci_ad_i_26_;
wire pci_ad_i_27_;
wire pci_ad_i_28_;
wire pci_ad_i_29_;
wire pci_ad_i_2_;
wire pci_ad_i_30_;
wire pci_ad_i_31_;
wire pci_ad_i_3_;
wire pci_ad_i_4_;
wire pci_ad_i_5_;
wire pci_ad_i_6_;
wire pci_ad_i_7_;
wire pci_ad_i_8_;
wire pci_ad_i_9_;
wire pci_cbe_i_0_;
wire pci_cbe_i_1_;
wire pci_cbe_i_2_;
wire pci_cbe_i_3_;
wire pci_devsel_i;
wire pci_frame_i;
wire pci_gnt_i;
wire pci_idsel_i;
wire pci_irdy_i;
wire pci_par_i;
wire pci_perr_i;
wire pci_rst_i;
wire pci_rst_oe_o;
wire pci_stop_i;
wire pci_trdy_i;
wire wb_int_i;
wire wbm_ack_i;
wire wbm_dat_i_0_;
wire wbm_dat_i_10_;
wire wbm_dat_i_11_;
wire wbm_dat_i_12_;
wire wbm_dat_i_13_;
wire wbm_dat_i_14_;
wire wbm_dat_i_15_;
wire wbm_dat_i_16_;
wire wbm_dat_i_17_;
wire wbm_dat_i_18_;
wire wbm_dat_i_19_;
wire wbm_dat_i_1_;
wire wbm_dat_i_20_;
wire wbm_dat_i_21_;
wire wbm_dat_i_22_;
wire wbm_dat_i_23_;
wire wbm_dat_i_24_;
wire wbm_dat_i_25_;
wire wbm_dat_i_26_;
wire wbm_dat_i_27_;
wire wbm_dat_i_28_;
wire wbm_dat_i_29_;
wire wbm_dat_i_2_;
wire wbm_dat_i_30_;
wire wbm_dat_i_31_;
wire wbm_dat_i_3_;
wire wbm_dat_i_4_;
wire wbm_dat_i_5_;
wire wbm_dat_i_6_;
wire wbm_dat_i_7_;
wire wbm_dat_i_8_;
wire wbm_dat_i_9_;
wire wbm_err_i;
wire wbm_rty_i;
wire wbs_adr_i_0_;
wire wbs_adr_i_10_;
wire wbs_adr_i_11_;
wire wbs_adr_i_12_;
wire wbs_adr_i_13_;
wire wbs_adr_i_14_;
wire wbs_adr_i_15_;
wire wbs_adr_i_16_;
wire wbs_adr_i_17_;
wire wbs_adr_i_18_;
wire wbs_adr_i_19_;
wire wbs_adr_i_1_;
wire wbs_adr_i_20_;
wire wbs_adr_i_21_;
wire wbs_adr_i_22_;
wire wbs_adr_i_23_;
wire wbs_adr_i_24_;
wire wbs_adr_i_25_;
wire wbs_adr_i_26_;
wire wbs_adr_i_27_;
wire wbs_adr_i_28_;
wire wbs_adr_i_29_;
wire wbs_adr_i_2_;
wire wbs_adr_i_30_;
wire wbs_adr_i_31_;
wire wbs_adr_i_3_;
wire wbs_adr_i_4_;
wire wbs_adr_i_5_;
wire wbs_adr_i_6_;
wire wbs_adr_i_7_;
wire wbs_adr_i_8_;
wire wbs_adr_i_9_;
wire wbs_bte_i_0_;
wire wbs_bte_i_1_;
wire wbs_cti_i_0_;
wire wbs_cti_i_1_;
wire wbs_cti_i_2_;
wire wbs_cyc_i;
wire wbs_dat_i_0_;
wire wbs_dat_i_10_;
wire wbs_dat_i_11_;
wire wbs_dat_i_12_;
wire wbs_dat_i_13_;
wire wbs_dat_i_14_;
wire wbs_dat_i_15_;
wire wbs_dat_i_16_;
wire wbs_dat_i_17_;
wire wbs_dat_i_18_;
wire wbs_dat_i_19_;
wire wbs_dat_i_1_;
wire wbs_dat_i_20_;
wire wbs_dat_i_21_;
wire wbs_dat_i_22_;
wire wbs_dat_i_23_;
wire wbs_dat_i_24_;
wire wbs_dat_i_25_;
wire wbs_dat_i_26_;
wire wbs_dat_i_27_;
wire wbs_dat_i_28_;
wire wbs_dat_i_29_;
wire wbs_dat_i_2_;
wire wbs_dat_i_30_;
wire wbs_dat_i_31_;
wire wbs_dat_i_3_;
wire wbs_dat_i_4_;
wire wbs_dat_i_5_;
wire wbs_dat_i_6_;
wire wbs_dat_i_7_;
wire wbs_dat_i_8_;
wire wbs_dat_i_9_;
wire wbs_sel_i_0_;
wire wbs_sel_i_1_;
wire wbs_sel_i_2_;
wire wbs_sel_i_3_;
wire wbs_stb_i;
wire wbs_we_i;
wire pci_ad_o_0_;
wire pci_ad_o_10_;
wire pci_ad_o_11_;
wire pci_ad_o_12_;
wire pci_ad_o_13_;
wire pci_ad_o_14_;
wire pci_ad_o_15_;
wire pci_ad_o_16_;
wire pci_ad_o_17_;
wire pci_ad_o_18_;
wire pci_ad_o_19_;
wire pci_ad_o_1_;
wire pci_ad_o_20_;
wire pci_ad_o_21_;
wire pci_ad_o_22_;
wire pci_ad_o_23_;
wire pci_ad_o_24_;
wire pci_ad_o_25_;
wire pci_ad_o_26_;
wire pci_ad_o_27_;
wire pci_ad_o_28_;
wire pci_ad_o_29_;
wire pci_ad_o_2_;
wire pci_ad_o_30_;
wire pci_ad_o_31_;
wire pci_ad_o_3_;
wire pci_ad_o_4_;
wire pci_ad_o_5_;
wire pci_ad_o_6_;
wire pci_ad_o_7_;
wire pci_ad_o_8_;
wire pci_ad_o_9_;
wire pci_ad_oe_o_0_;
wire pci_ad_oe_o_10_;
wire pci_ad_oe_o_11_;
wire pci_ad_oe_o_12_;
wire pci_ad_oe_o_13_;
wire pci_ad_oe_o_14_;
wire pci_ad_oe_o_15_;
wire pci_ad_oe_o_16_;
wire pci_ad_oe_o_17_;
wire pci_ad_oe_o_18_;
wire pci_ad_oe_o_19_;
wire pci_ad_oe_o_1_;
wire pci_ad_oe_o_20_;
wire pci_ad_oe_o_21_;
wire pci_ad_oe_o_22_;
wire pci_ad_oe_o_23_;
wire pci_ad_oe_o_24_;
wire pci_ad_oe_o_25_;
wire pci_ad_oe_o_26_;
wire pci_ad_oe_o_27_;
wire pci_ad_oe_o_28_;
wire pci_ad_oe_o_29_;
wire pci_ad_oe_o_2_;
wire pci_ad_oe_o_30_;
wire pci_ad_oe_o_31_;
wire pci_ad_oe_o_3_;
wire pci_ad_oe_o_4_;
wire pci_ad_oe_o_5_;
wire pci_ad_oe_o_6_;
wire pci_ad_oe_o_7_;
wire pci_ad_oe_o_8_;
wire pci_ad_oe_o_9_;
wire pci_cbe_o_0_;
wire pci_cbe_o_1_;
wire pci_cbe_o_2_;
wire pci_cbe_o_3_;
wire pci_cbe_oe_o_0_;
wire pci_cbe_oe_o_1_;
wire pci_cbe_oe_o_2_;
wire pci_cbe_oe_o_3_;
wire pci_devsel_o;
wire pci_devsel_oe_o;
wire pci_frame_o;
wire pci_frame_oe_o;
wire pci_inta_oe_o;
wire pci_irdy_o;
wire pci_irdy_oe_o;
wire pci_par_o;
wire pci_par_oe_o;
wire pci_perr_o;
wire pci_perr_oe_o;
wire pci_req_o;
wire pci_req_oe_o;
wire pci_serr_o;
wire pci_serr_oe_o;
wire pci_stop_o;
wire pci_stop_oe_o;
wire pci_trdy_o;
wire pci_trdy_oe_o;
wire wb_rst_o;
wire wbm_adr_o_0_;
wire wbm_adr_o_10_;
wire wbm_adr_o_11_;
wire wbm_adr_o_12_;
wire wbm_adr_o_13_;
wire wbm_adr_o_14_;
wire wbm_adr_o_15_;
wire wbm_adr_o_16_;
wire wbm_adr_o_17_;
wire wbm_adr_o_18_;
wire wbm_adr_o_19_;
wire wbm_adr_o_1_;
wire wbm_adr_o_20_;
wire wbm_adr_o_21_;
wire wbm_adr_o_22_;
wire wbm_adr_o_23_;
wire wbm_adr_o_24_;
wire wbm_adr_o_25_;
wire wbm_adr_o_26_;
wire wbm_adr_o_27_;
wire wbm_adr_o_28_;
wire wbm_adr_o_29_;
wire wbm_adr_o_2_;
wire wbm_adr_o_30_;
wire wbm_adr_o_31_;
wire wbm_adr_o_3_;
wire wbm_adr_o_4_;
wire wbm_adr_o_5_;
wire wbm_adr_o_6_;
wire wbm_adr_o_7_;
wire wbm_adr_o_8_;
wire wbm_adr_o_9_;
wire wbm_cti_o_0_;
wire wbm_cti_o_1_;
wire wbm_cti_o_2_;
wire wbm_cyc_o;
wire wbm_dat_o_0_;
wire wbm_dat_o_10_;
wire wbm_dat_o_11_;
wire wbm_dat_o_12_;
wire wbm_dat_o_13_;
wire wbm_dat_o_14_;
wire wbm_dat_o_15_;
wire wbm_dat_o_16_;
wire wbm_dat_o_17_;
wire wbm_dat_o_18_;
wire wbm_dat_o_19_;
wire wbm_dat_o_1_;
wire wbm_dat_o_20_;
wire wbm_dat_o_21_;
wire wbm_dat_o_22_;
wire wbm_dat_o_23_;
wire wbm_dat_o_24_;
wire wbm_dat_o_25_;
wire wbm_dat_o_26_;
wire wbm_dat_o_27_;
wire wbm_dat_o_28_;
wire wbm_dat_o_29_;
wire wbm_dat_o_2_;
wire wbm_dat_o_30_;
wire wbm_dat_o_31_;
wire wbm_dat_o_3_;
wire wbm_dat_o_4_;
wire wbm_dat_o_5_;
wire wbm_dat_o_6_;
wire wbm_dat_o_7_;
wire wbm_dat_o_8_;
wire wbm_dat_o_9_;
wire wbm_sel_o_0_;
wire wbm_sel_o_1_;
wire wbm_sel_o_2_;
wire wbm_sel_o_3_;
wire wbm_stb_o;
wire wbm_we_o;
wire wbs_ack_o;
wire wbs_dat_o_0_;
wire wbs_dat_o_10_;
wire wbs_dat_o_11_;
wire wbs_dat_o_12_;
wire wbs_dat_o_13_;
wire wbs_dat_o_14_;
wire wbs_dat_o_15_;
wire wbs_dat_o_16_;
wire wbs_dat_o_17_;
wire wbs_dat_o_18_;
wire wbs_dat_o_19_;
wire wbs_dat_o_1_;
wire wbs_dat_o_20_;
wire wbs_dat_o_21_;
wire wbs_dat_o_22_;
wire wbs_dat_o_23_;
wire wbs_dat_o_24_;
wire wbs_dat_o_25_;
wire wbs_dat_o_26_;
wire wbs_dat_o_27_;
wire wbs_dat_o_28_;
wire wbs_dat_o_29_;
wire wbs_dat_o_2_;
wire wbs_dat_o_30_;
wire wbs_dat_o_31_;
wire wbs_dat_o_3_;
wire wbs_dat_o_4_;
wire wbs_dat_o_5_;
wire wbs_dat_o_6_;
wire wbs_dat_o_7_;
wire wbs_dat_o_8_;
wire wbs_dat_o_9_;
wire wbs_err_o;
wire wbs_rty_o;
wire FE_OCPN1822_n_16560;
wire FE_OCPN1823_n_16560;
wire FE_OCPN1824_n_12030;
wire FE_OCPN1825_n_12030;
wire FE_OCPN1827_n_14995;
wire FE_OCPN1831_n_16949;
wire FE_OCPN1832_n_16949;
wire FE_OCPN1833_n_11884;
wire FE_OCPN1834_n_11884;
wire FE_OCPN1835_n_16798;
wire FE_OCPN1836_n_16798;
wire FE_OCPN1837_n_1238;
wire FE_OCPN1838_n_1238;
wire FE_OCPN1839_n_1238;
wire FE_OCPN1840_n_16089;
wire FE_OCPN1841_n_16089;
wire FE_OCPN1842_n_16033;
wire FE_OCPN1843_n_16033;
wire FE_OCPN1844_n_16427;
wire FE_OCPN1845_n_16427;
wire FE_OCPN1846_n_14981;
wire FE_OCPN1847_n_14981;
wire FE_OCPN1848_n_15998;
wire FE_OCPN1849_n_15998;
wire FE_OCPN1850_n_15998;
wire FE_OCPN1851_n_16538;
wire FE_OCPN1852_n_16538;
wire FE_OCPN1853_n_2071;
wire FE_OCPN1854_n_2071;
wire FE_OCPN1855_n_2071;
wire FE_OCPN1856_FE_OFN1774_n_13800;
wire FE_OCPN1860_FE_OFN468_n_15534;
wire FE_OCPN1861_FE_OFN468_n_15534;
wire FE_OCPN1862_FE_OFN474_n_16992;
wire FE_OCPN1863_FE_OFN474_n_16992;
wire FE_OCPN1865_n_12377;
wire FE_OCPN1866_n_12377;
wire FE_OCPN1868_n_16289;
wire FE_OCPN1871_FE_OFN474_n_16992;
wire FE_OCPN1872_FE_OFN474_n_16992;
wire FE_OCPN1873_FE_OFN474_n_16992;
wire FE_OCPN1875_n_14526;
wire FE_OCPN1876_n_13903;
wire FE_OCPN1877_n_13903;
wire FE_OCPN1878_FE_OFN470_n_10588;
wire FE_OCPN1879_FE_OFN470_n_10588;
wire FE_OCPN1880_n_9991;
wire FE_OCPN1881_n_9991;
wire FE_OCPN1882_n_9991;
wire FE_OCPN1883_n_15566;
wire FE_OCPN1884_n_15566;
wire FE_OCPN1885_FE_OFN1508_n_15587;
wire FE_OCPN1886_FE_OFN1508_n_15587;
wire FE_OCPN1887_FE_OFN473_n_16992;
wire FE_OCPN1888_FE_OFN473_n_16992;
wire FE_OCPN1889_n_16553;
wire FE_OCPN1890_n_16553;
wire FE_OCPN1891_FE_OFN1727_n_9975;
wire FE_OCPN1892_FE_OFN1727_n_9975;
wire FE_OCPN1895_FE_OFN1559_n_12042;
wire FE_OCPN1897_n_3231;
wire FE_OCPN1898_n_3231;
wire FE_OCPN1899_n_16810;
wire FE_OCPN1900_n_16810;
wire FE_OCPN1901_n_16810;
wire FE_OCPN1902_FE_OFN1061_n_16720;
wire FE_OCPN1903_FE_OFN1061_n_16720;
wire FE_OCPN1904_n_8927;
wire FE_OCPN1905_n_8927;
wire FE_OCPN1907_n_11767;
wire FE_OCPN1908_n_16497;
wire FE_OCPN1909_n_16497;
wire FE_OCPN1910_FE_OFN1152_n_13249;
wire FE_OCPN1911_FE_OFN1152_n_13249;
wire FE_OCPN1912_FE_OFN1150_n_13249;
wire FE_OCPN1913_FE_OFN1150_n_13249;
wire FE_OCPN1914_FE_OFN1522_n_10892;
wire FE_OCPN1915_FE_OFN1522_n_10892;
wire FE_OCPN2014_n_10195;
wire FE_OCPN2015_n_10195;
wire FE_OCPN2217_n_13997;
wire FE_OCPN2218_n_13997;
wire FE_OCPN2219_n_13997;
wire FE_OCPUNCON1951_FE_OFN697_n_16760;
wire FE_OCPUNCON1952_FE_OFN697_n_16760;
wire FE_OCP_DRV_N1949_n_8660;
wire FE_OCP_DRV_N1950_n_8660;
wire FE_OCP_DRV_N2261_n_8660;
wire FE_OCP_DRV_N2262_n_8660;
wire FE_OCP_RBN1917_wbs_cti_i_1_;
wire FE_OCP_RBN1918_wbs_cti_i_1_;
wire FE_OCP_RBN1921_n_10273;
wire FE_OCP_RBN1922_n_10273;
wire FE_OCP_RBN1923_n_10273;
wire FE_OCP_RBN1924_n_10273;
wire FE_OCP_RBN1925_n_10259;
wire FE_OCP_RBN1926_n_10259;
wire FE_OCP_RBN1927_n_10259;
wire FE_OCP_RBN1928_n_10259;
wire FE_OCP_RBN1929_parchk_pci_trdy_reg_in;
wire FE_OCP_RBN1930_parchk_pci_trdy_reg_in;
wire FE_OCP_RBN1932_FE_OFN1515_n_10538;
wire FE_OCP_RBN1933_FE_OFN1515_n_10538;
wire FE_OCP_RBN1934_FE_OFN1515_n_10538;
wire FE_OCP_RBN1954_FE_RN_462_0;
wire FE_OCP_RBN1955_n_16981;
wire FE_OCP_RBN1956_n_16981;
wire FE_OCP_RBN1961_FE_OFN1591_n_13741;
wire FE_OCP_RBN1962_FE_OFN1591_n_13741;
wire FE_OCP_RBN1963_FE_OFN1591_n_13741;
wire FE_OCP_RBN1964_FE_OFN1591_n_13741;
wire FE_OCP_RBN1965_FE_RN_459_0;
wire FE_OCP_RBN1966_FE_RN_459_0;
wire FE_OCP_RBN1967_FE_RN_459_0;
wire FE_OCP_RBN1968_FE_OFN1532_n_10143;
wire FE_OCP_RBN1969_FE_OFN1532_n_10143;
wire FE_OCP_RBN1970_n_11767;
wire FE_OCP_RBN1971_n_11767;
wire FE_OCP_RBN1972_n_11767;
wire FE_OCP_RBN1973_n_12381;
wire FE_OCP_RBN1974_n_12381;
wire FE_OCP_RBN1975_n_12381;
wire FE_OCP_RBN1976_n_12381;
wire FE_OCP_RBN1977_n_10273;
wire FE_OCP_RBN1978_n_10273;
wire FE_OCP_RBN1979_n_10273;
wire FE_OCP_RBN1980_n_10273;
wire FE_OCP_RBN1981_FE_OFN1591_n_13741;
wire FE_OCP_RBN1983_FE_OFN1591_n_13741;
wire FE_OCP_RBN1984_FE_OFN1591_n_13741;
wire FE_OCP_RBN1985_FE_OFN1591_n_13741;
wire FE_OCP_RBN1994_n_13971;
wire FE_OCP_RBN1995_n_13971;
wire FE_OCP_RBN1996_n_13971;
wire FE_OCP_RBN1997_n_13971;
wire FE_OCP_RBN1998_n_13971;
wire FE_OCP_RBN1999_n_13971;
wire FE_OCP_RBN2000_n_1403;
wire FE_OCP_RBN2003_FE_OFN1026_n_16760;
wire FE_OCP_RBN2004_FE_OFN1026_n_16760;
wire FE_OCP_RBN2005_FE_RN_459_0;
wire FE_OCP_RBN2006_FE_RN_459_0;
wire FE_OCP_RBN2007_n_16698;
wire FE_OCP_RBN2008_n_16698;
wire FE_OCP_RBN2009_n_16698;
wire FE_OCP_RBN2010_n_16698;
wire FE_OCP_RBN2011_n_16698;
wire FE_OCP_RBN2012_n_16698;
wire FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042;
wire FE_OCP_RBN2016_n_16970;
wire FE_OCP_RBN2017_n_16970;
wire FE_OCP_RBN2018_n_16970;
wire FE_OCP_RBN2019_n_16970;
wire FE_OCP_RBN2220_n_15347;
wire FE_OCP_RBN2221_n_15347;
wire FE_OCP_RBN2222_n_15347;
wire FE_OCP_RBN2223_n_15347;
wire FE_OCP_RBN2224_n_16322;
wire FE_OCP_RBN2225_n_16322;
wire FE_OCP_RBN2226_g75174_p;
wire FE_OCP_RBN2227_g75174_p;
wire FE_OCP_RBN2228_n_15969;
wire FE_OCP_RBN2229_n_15969;
wire FE_OCP_RBN2231_FE_RN_390_0;
wire FE_OCP_RBN2232_n_16273;
wire FE_OCP_RBN2233_n_16273;
wire FE_OCP_RBN2237_g74749_p;
wire FE_OCP_RBN2238_g74749_p;
wire FE_OCP_RBN2239_g74749_p;
wire FE_OCP_RBN2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_;
wire FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_;
wire FE_OCP_RBN2270_g75061_p;
wire FE_OCP_RBN2271_g75061_p;
wire FE_OCP_RBN2272_n_10268;
wire FE_OCP_RBN2273_n_10268;
wire FE_OCP_RBN2274_n_10268;
wire FE_OCP_RBN2275_n_10268;
wire FE_OCP_RBN2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_;
wire FE_OCP_RBN2278_n_16974;
wire FE_OCP_RBN2279_n_16974;
wire FE_OCP_RBN2280_g74996_p;
wire FE_OCP_RBN2281_g74996_p;
wire FE_OCP_RBN2282_g74996_p;
wire FE_OCP_RBN2283_g74996_p;
wire FE_OCP_RBN2284_FE_RN_494_0;
wire FE_OCP_RBN2285_FE_RN_494_0;
wire FE_OCP_RBN2286_FE_RN_494_0;
wire FE_OCP_RBN2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_;
wire FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_;
wire FE_OCP_RBN2291_FE_OFN1575_n_12028;
wire FE_OCP_RBN2292_FE_OFN1575_n_12028;
wire FE_OCP_RBN2293_FE_OFN1581_n_12306;
wire FE_OFN1000_n_15978;
wire FE_OFN1001_n_15978;
wire FE_OFN1002_n_2047;
wire FE_OFN1003_n_2047;
wire FE_OFN1004_n_16288;
wire FE_OFN1005_n_16288;
wire FE_OFN1006_n_16288;
wire FE_OFN1007_n_4734;
wire FE_OFN1008_n_4734;
wire FE_OFN1009_n_4734;
wire FE_OFN1010_n_4734;
wire FE_OFN1011_n_4734;
wire FE_OFN1012_n_4734;
wire FE_OFN1013_n_4734;
wire FE_OFN1014_n_2053;
wire FE_OFN1015_n_2053;
wire FE_OFN1016_n_2053;
wire FE_OFN1017_n_2053;
wire FE_OFN1018_n_11877;
wire FE_OFN1019_n_11877;
wire FE_OFN1020_n_11877;
wire FE_OFN1021_n_11877;
wire FE_OFN1022_n_11877;
wire FE_OFN1023_n_11877;
wire FE_OFN1024_n_11877;
wire FE_OFN1025_n_11877;
wire FE_OFN1026_n_16760;
wire FE_OFN1028_n_4732;
wire FE_OFN1029_n_4732;
wire FE_OFN1030_n_4732;
wire FE_OFN1031_n_4732;
wire FE_OFN1032_n_4732;
wire FE_OFN1033_n_4732;
wire FE_OFN1034_n_4732;
wire FE_OFN1035_n_4732;
wire FE_OFN1036_n_4732;
wire FE_OFN1037_n_4732;
wire FE_OFN1038_n_2037;
wire FE_OFN1039_n_2037;
wire FE_OFN1040_n_2037;
wire FE_OFN1041_n_2037;
wire FE_OFN1042_n_2037;
wire FE_OFN1043_n_2037;
wire FE_OFN1044_n_2037;
wire FE_OFN1045_n_16657;
wire FE_OFN1046_n_16657;
wire FE_OFN1047_n_16657;
wire FE_OFN1048_n_16657;
wire FE_OFN1049_n_16657;
wire FE_OFN1050_n_16657;
wire FE_OFN1051_n_16657;
wire FE_OFN1052_n_4727;
wire FE_OFN1053_n_4727;
wire FE_OFN1054_n_4727;
wire FE_OFN1055_n_4727;
wire FE_OFN1056_n_4727;
wire FE_OFN1057_n_4727;
wire FE_OFN1058_n_4727;
wire FE_OFN1059_n_4727;
wire FE_OFN1060_n_16720;
wire FE_OFN1061_n_16720;
wire FE_OFN1062_n_15808;
wire FE_OFN1063_n_15808;
wire FE_OFN1064_n_15808;
wire FE_OFN1065_n_15808;
wire FE_OFN1066_n_15808;
wire FE_OFN1067_n_15729;
wire FE_OFN1068_n_15729;
wire FE_OFN1069_n_15729;
wire FE_OFN1070_n_15729;
wire FE_OFN1071_n_15729;
wire FE_OFN1072_n_4740;
wire FE_OFN1073_n_4740;
wire FE_OFN1074_n_4740;
wire FE_OFN1075_n_4740;
wire FE_OFN1076_n_4740;
wire FE_OFN1077_n_4740;
wire FE_OFN1078_n_4778;
wire FE_OFN1079_n_4778;
wire FE_OFN1080_n_13221;
wire FE_OFN1081_n_13221;
wire FE_OFN1082_n_13221;
wire FE_OFN1083_n_13221;
wire FE_OFN1084_n_13221;
wire FE_OFN1085_n_13221;
wire FE_OFN1086_g64577_p;
wire FE_OFN1087_g64577_p;
wire FE_OFN1088_g64577_p;
wire FE_OFN1089_g64577_p;
wire FE_OFN1090_g64577_p;
wire FE_OFN1091_g64577_p;
wire FE_OFN1092_g64577_p;
wire FE_OFN1093_g64577_p;
wire FE_OFN1094_g64577_p;
wire FE_OFN1095_g64577_p;
wire FE_OFN1096_g64577_p;
wire FE_OFN1097_g64577_p;
wire FE_OFN1098_g64577_p;
wire FE_OFN1099_g64577_p;
wire FE_OFN1100_g64577_p;
wire FE_OFN1101_g64577_p;
wire FE_OFN1102_g64577_p;
wire FE_OFN1103_g64577_p;
wire FE_OFN1104_g64577_p;
wire FE_OFN1105_g64577_p;
wire FE_OFN1106_g64577_p;
wire FE_OFN1107_g64577_p;
wire FE_OFN1108_g64577_p;
wire FE_OFN1109_g64577_p;
wire FE_OFN1110_g64577_p;
wire FE_OFN1111_g64577_p;
wire FE_OFN1112_g64577_p;
wire FE_OFN1113_g64577_p;
wire FE_OFN1114_g64577_p;
wire FE_OFN1115_g64577_p;
wire FE_OFN1116_g64577_p;
wire FE_OFN1117_g64577_p;
wire FE_OFN1118_g64577_p;
wire FE_OFN1119_g64577_p;
wire FE_OFN1120_g64577_p;
wire FE_OFN1121_g64577_p;
wire FE_OFN1122_g64577_p;
wire FE_OFN1123_g64577_p;
wire FE_OFN1124_g64577_p;
wire FE_OFN1125_g64577_p;
wire FE_OFN1126_g64577_p;
wire FE_OFN1127_g64577_p;
wire FE_OFN1128_g64577_p;
wire FE_OFN1129_g64577_p;
wire FE_OFN1130_g64577_p;
wire FE_OFN1131_g64577_p;
wire FE_OFN1132_g64577_p;
wire FE_OFN1133_g64577_p;
wire FE_OFN1134_g64577_p;
wire FE_OFN1135_g64577_p;
wire FE_OFN1136_g64577_p;
wire FE_OFN1137_g64577_p;
wire FE_OFN1138_g64577_p;
wire FE_OFN1139_g64577_p;
wire FE_OFN1140_g64577_p;
wire FE_OFN1141_n_15261;
wire FE_OFN1142_n_15261;
wire FE_OFN1143_n_15261;
wire FE_OFN1144_n_15261;
wire FE_OFN1145_n_15261;
wire FE_OFN1146_n_13249;
wire FE_OFN1147_n_13249;
wire FE_OFN1148_n_13249;
wire FE_OFN1149_n_13249;
wire FE_OFN1150_n_13249;
wire FE_OFN1151_n_13249;
wire FE_OFN1152_n_13249;
wire FE_OFN1153_n_3464;
wire FE_OFN1154_n_3464;
wire FE_OFN1155_n_3464;
wire FE_OFN1156_n_7498;
wire FE_OFN1157_n_15325;
wire FE_OFN1158_n_15325;
wire FE_OFN1159_n_15325;
wire FE_OFN1160_n_5615;
wire FE_OFN1161_n_5615;
wire FE_OFN1162_n_5615;
wire FE_OFN1163_n_5615;
wire FE_OFN1164_n_5615;
wire FE_OFN1165_n_5615;
wire FE_OFN1166_n_5615;
wire FE_OFN1167_n_5592;
wire FE_OFN1168_n_5592;
wire FE_OFN1169_n_5592;
wire FE_OFN1170_n_5592;
wire FE_OFN1171_n_5592;
wire FE_OFN1172_n_5592;
wire FE_OFN1173_n_5592;
wire FE_OFN1174_n_5592;
wire FE_OFN1175_n_3476;
wire FE_OFN1176_n_3476;
wire FE_OFN1177_n_3476;
wire FE_OFN1178_n_3476;
wire FE_OFN1179_n_3476;
wire FE_OFN1180_n_3476;
wire FE_OFN1181_n_3476;
wire FE_OFN1182_n_3476;
wire FE_OFN1183_n_3476;
wire FE_OFN1184_n_3476;
wire FE_OFN1185_n_3476;
wire FE_OFN1186_n_3476;
wire FE_OFN1187_n_5742;
wire FE_OFN1188_n_5742;
wire FE_OFN1189_n_5742;
wire FE_OFN1190_n_6935;
wire FE_OFN1191_n_6935;
wire FE_OFN1192_n_6935;
wire FE_OFN1193_n_6935;
wire FE_OFN1194_n_6935;
wire FE_OFN1195_n_4090;
wire FE_OFN1196_n_4090;
wire FE_OFN1197_n_4090;
wire FE_OFN1198_n_4090;
wire FE_OFN1199_n_4090;
wire FE_OFN1200_n_4090;
wire FE_OFN1201_n_4090;
wire FE_OFN1202_n_4090;
wire FE_OFN1203_n_4090;
wire FE_OFN1204_n_4090;
wire FE_OFN1205_n_6356;
wire FE_OFN1206_n_6356;
wire FE_OFN1207_n_6356;
wire FE_OFN1208_n_6356;
wire FE_OFN1209_n_4151;
wire FE_OFN1210_n_4151;
wire FE_OFN1211_n_4151;
wire FE_OFN1212_n_4151;
wire FE_OFN1213_n_4151;
wire FE_OFN1214_n_4151;
wire FE_OFN1215_n_4151;
wire FE_OFN1216_n_4151;
wire FE_OFN1217_n_6886;
wire FE_OFN1218_n_6886;
wire FE_OFN1219_n_6886;
wire FE_OFN1220_n_6391;
wire FE_OFN1221_n_6391;
wire FE_OFN1222_n_6391;
wire FE_OFN1223_n_6391;
wire FE_OFN1224_n_6391;
wire FE_OFN1225_n_6391;
wire FE_OFN1226_n_6391;
wire FE_OFN1227_n_6391;
wire FE_OFN1228_n_6391;
wire FE_OFN1229_n_6391;
wire FE_OFN1230_n_6391;
wire FE_OFN1231_n_6391;
wire FE_OFN1232_n_6391;
wire FE_OFN1233_n_6391;
wire FE_OFN1234_n_6391;
wire FE_OFN1235_n_6391;
wire FE_OFN1236_n_6391;
wire FE_OFN1237_n_4092;
wire FE_OFN1238_n_4092;
wire FE_OFN1239_n_4092;
wire FE_OFN1240_n_4092;
wire FE_OFN1241_n_4092;
wire FE_OFN1242_n_4092;
wire FE_OFN1243_n_4092;
wire FE_OFN1244_n_4092;
wire FE_OFN1245_n_4093;
wire FE_OFN1246_n_4093;
wire FE_OFN1247_n_4093;
wire FE_OFN1248_n_4093;
wire FE_OFN1249_n_4093;
wire FE_OFN1250_n_4093;
wire FE_OFN1251_n_4143;
wire FE_OFN1252_n_4143;
wire FE_OFN1253_n_4143;
wire FE_OFN1254_n_4143;
wire FE_OFN1255_n_4143;
wire FE_OFN1256_n_4143;
wire FE_OFN1257_n_4143;
wire FE_OFN1258_n_4143;
wire FE_OFN1259_n_4143;
wire FE_OFN1260_n_4143;
wire FE_OFN1261_n_4143;
wire FE_OFN1262_n_4095;
wire FE_OFN1263_n_4095;
wire FE_OFN1264_n_4095;
wire FE_OFN1265_n_4095;
wire FE_OFN1266_n_4095;
wire FE_OFN1267_n_4095;
wire FE_OFN1268_n_4095;
wire FE_OFN1269_n_4095;
wire FE_OFN1270_n_4095;
wire FE_OFN1271_n_4096;
wire FE_OFN1272_n_4096;
wire FE_OFN1273_n_4096;
wire FE_OFN1274_n_4096;
wire FE_OFN1275_n_4096;
wire FE_OFN1276_n_4096;
wire FE_OFN1277_n_4097;
wire FE_OFN1278_n_4097;
wire FE_OFN1279_n_4097;
wire FE_OFN1280_n_4097;
wire FE_OFN1281_n_4097;
wire FE_OFN1282_n_4097;
wire FE_OFN1283_n_4097;
wire FE_OFN1284_n_4097;
wire FE_OFN1285_n_4097;
wire FE_OFN1286_n_4098;
wire FE_OFN1287_n_4098;
wire FE_OFN1288_n_4098;
wire FE_OFN1289_n_4098;
wire FE_OFN1290_n_4098;
wire FE_OFN1291_n_4098;
wire FE_OFN1292_n_4098;
wire FE_OFN1293_n_4098;
wire FE_OFN1294_n_4098;
wire FE_OFN1295_n_4098;
wire FE_OFN1296_n_5763;
wire FE_OFN1297_n_5763;
wire FE_OFN1298_n_5763;
wire FE_OFN1299_n_5763;
wire FE_OFN1300_n_5763;
wire FE_OFN1301_n_5763;
wire FE_OFN1302_n_5763;
wire FE_OFN1303_n_13124;
wire FE_OFN1304_n_13124;
wire FE_OFN1305_n_13124;
wire FE_OFN1306_n_13124;
wire FE_OFN1307_n_6624;
wire FE_OFN1308_n_6624;
wire FE_OFN1309_n_6624;
wire FE_OFN1310_n_6624;
wire FE_OFN1311_n_6624;
wire FE_OFN1312_n_6624;
wire FE_OFN1313_n_6624;
wire FE_OFN1314_n_6624;
wire FE_OFN1315_n_6624;
wire FE_OFN1316_n_6624;
wire FE_OFN1317_n_6624;
wire FE_OFN1318_n_6436;
wire FE_OFN1319_n_6436;
wire FE_OFN1320_n_6436;
wire FE_OFN1321_n_6436;
wire FE_OFN1322_n_6436;
wire FE_OFN1323_n_6436;
wire FE_OFN1324_n_13547;
wire FE_OFN1325_n_13547;
wire FE_OFN1326_n_13547;
wire FE_OFN1327_n_13547;
wire FE_OFN1328_n_13547;
wire FE_OFN1329_n_13547;
wire FE_OFN1330_n_13547;
wire FE_OFN1331_n_13547;
wire FE_OFN1332_n_13547;
wire FE_OFN1333_n_13547;
wire FE_OFN1334_n_13720;
wire FE_OFN1335_n_13720;
wire FE_OFN1336_n_16439;
wire FE_OFN1337_n_16439;
wire FE_OFN1338_n_8567;
wire FE_OFN1339_n_8567;
wire FE_OFN1340_n_8567;
wire FE_OFN1341_n_8567;
wire FE_OFN1342_n_8567;
wire FE_OFN1343_n_8567;
wire FE_OFN1344_n_8567;
wire FE_OFN1345_n_8567;
wire FE_OFN1346_n_8567;
wire FE_OFN1347_n_8567;
wire FE_OFN1348_n_8567;
wire FE_OFN1349_n_8567;
wire FE_OFN1350_n_8567;
wire FE_OFN1351_n_8567;
wire FE_OFN1352_n_8567;
wire FE_OFN1353_n_8567;
wire FE_OFN1354_n_8567;
wire FE_OFN1355_n_8567;
wire FE_OFN1356_n_8567;
wire FE_OFN1357_n_8567;
wire FE_OFN1358_n_8567;
wire FE_OFN1359_n_8567;
wire FE_OFN1360_n_8567;
wire FE_OFN1361_n_8567;
wire FE_OFN1362_n_8567;
wire FE_OFN1363_n_8567;
wire FE_OFN1364_n_8567;
wire FE_OFN1365_n_8567;
wire FE_OFN1366_n_8567;
wire FE_OFN1367_n_8567;
wire FE_OFN1368_n_8567;
wire FE_OFN1369_n_8567;
wire FE_OFN1370_n_8567;
wire FE_OFN1371_n_8567;
wire FE_OFN1372_n_8567;
wire FE_OFN1373_n_8567;
wire FE_OFN1374_n_8567;
wire FE_OFN1376_n_8567;
wire FE_OFN1377_n_8567;
wire FE_OFN1378_n_8567;
wire FE_OFN1379_n_8567;
wire FE_OFN1380_n_8567;
wire FE_OFN1381_n_8567;
wire FE_OFN1382_n_8567;
wire FE_OFN1383_n_8567;
wire FE_OFN1384_n_8567;
wire FE_OFN1385_n_8567;
wire FE_OFN1386_n_8567;
wire FE_OFN1387_n_8567;
wire FE_OFN1388_n_8567;
wire FE_OFN1389_n_8567;
wire FE_OFN1390_n_8567;
wire FE_OFN1391_n_8567;
wire FE_OFN1392_n_8567;
wire FE_OFN1394_n_8567;
wire FE_OFN1396_n_8567;
wire FE_OFN1397_n_8567;
wire FE_OFN1398_n_8567;
wire FE_OFN1399_n_8567;
wire FE_OFN1400_n_8567;
wire FE_OFN1401_n_8567;
wire FE_OFN1402_n_8567;
wire FE_OFN1403_n_8567;
wire FE_OFN1404_n_8567;
wire FE_OFN1405_n_8567;
wire FE_OFN1406_n_8567;
wire FE_OFN1407_n_8567;
wire FE_OFN1408_n_8567;
wire FE_OFN1409_n_8567;
wire FE_OFN1410_n_8567;
wire FE_OFN1411_n_8567;
wire FE_OFN1412_n_8567;
wire FE_OFN1413_n_8567;
wire FE_OFN1414_n_8567;
wire FE_OFN1415_n_8567;
wire FE_OFN1416_n_8567;
wire FE_OFN1417_n_8567;
wire FE_OFN1419_n_8567;
wire FE_OFN1420_n_8567;
wire FE_OFN1421_n_8567;
wire FE_OFN1422_n_8567;
wire FE_OFN1423_n_8567;
wire FE_OFN1424_n_8567;
wire FE_OFN1425_n_8567;
wire FE_OFN1426_n_8567;
wire FE_OFN1427_n_8567;
wire FE_OFN1428_n_8567;
wire FE_OFN1429_n_16779;
wire FE_OFN1430_n_16779;
wire FE_OFN1431_n_16779;
wire FE_OFN1432_n_16779;
wire FE_OFN1433_n_16779;
wire FE_OFN1434_n_9372;
wire FE_OFN1435_n_9372;
wire FE_OFN1436_n_9372;
wire FE_OFN1437_n_9372;
wire FE_OFN1438_n_9372;
wire FE_OFN1439_n_9372;
wire FE_OFN1440_n_9372;
wire FE_OFN1441_n_9372;
wire FE_OFN1442_n_11125;
wire FE_OFN1443_n_11125;
wire FE_OFN1444_n_11125;
wire FE_OFN1445_n_11125;
wire FE_OFN1446_n_11125;
wire FE_OFN1447_n_9163;
wire FE_OFN1448_n_9163;
wire FE_OFN1449_n_9163;
wire FE_OFN1450_n_9163;
wire FE_OFN1451_n_10588;
wire FE_OFN1452_n_10588;
wire FE_OFN1453_n_10588;
wire FE_OFN1454_n_11138;
wire FE_OFN1455_n_11138;
wire FE_OFN1456_n_11138;
wire FE_OFN1457_n_11138;
wire FE_OFN1458_n_11138;
wire FE_OFN1459_n_11795;
wire FE_OFN1460_n_11795;
wire FE_OFN1461_n_11795;
wire FE_OFN1462_n_11795;
wire FE_OFN1463_n_10789;
wire FE_OFN1464_n_10789;
wire FE_OFN1465_n_10789;
wire FE_OFN1466_n_10789;
wire FE_OFN1467_n_10789;
wire FE_OFN1468_n_10789;
wire FE_OFN1469_g52675_p;
wire FE_OFN146_g65530_p;
wire FE_OFN1470_g52675_p;
wire FE_OFN1471_g52675_p;
wire FE_OFN1472_g52675_p;
wire FE_OFN1473_n_16637;
wire FE_OFN1474_n_16637;
wire FE_OFN1475_n_16637;
wire FE_OFN1477_n_16637;
wire FE_OFN1478_n_16637;
wire FE_OFN1479_n_16637;
wire FE_OFN147_g65530_p;
wire FE_OFN1480_n_15534;
wire FE_OFN1481_n_15534;
wire FE_OFN1483_n_15534;
wire FE_OFN1484_n_15534;
wire FE_OFN1485_n_15534;
wire FE_OFN1486_n_16992;
wire FE_OFN1487_n_9320;
wire FE_OFN1488_n_9320;
wire FE_OFN1489_n_9320;
wire FE_OFN1490_n_9320;
wire FE_OFN1491_n_9320;
wire FE_OFN1492_n_9320;
wire FE_OFN1493_n_9320;
wire FE_OFN1495_n_15558;
wire FE_OFN1496_n_15558;
wire FE_OFN1497_n_15558;
wire FE_OFN1498_n_15558;
wire FE_OFN1499_n_15558;
wire FE_OFN1500_n_15558;
wire FE_OFN1501_n_15558;
wire FE_OFN1502_n_15558;
wire FE_OFN1503_n_15768;
wire FE_OFN1505_n_15768;
wire FE_OFN1506_n_15768;
wire FE_OFN1507_n_15587;
wire FE_OFN1508_n_15587;
wire FE_OFN1509_n_15587;
wire FE_OFN1510_n_15587;
wire FE_OFN1511_n_15587;
wire FE_OFN1513_n_14987;
wire FE_OFN1514_n_10538;
wire FE_OFN1519_n_10892;
wire FE_OFN1520_n_10892;
wire FE_OFN1521_n_10892;
wire FE_OFN1522_n_10892;
wire FE_OFN1523_n_10892;
wire FE_OFN1524_n_10853;
wire FE_OFN1525_n_10853;
wire FE_OFN1526_n_10853;
wire FE_OFN1527_n_10853;
wire FE_OFN1528_n_10853;
wire FE_OFN1529_n_10853;
wire FE_OFN1530_n_10853;
wire FE_OFN1531_n_10143;
wire FE_OFN1532_n_10143;
wire FE_OFN1533_n_10143;
wire FE_OFN1535_n_10143;
wire FE_OFN1536_n_10143;
wire FE_OFN1537_n_10595;
wire FE_OFN1538_n_10595;
wire FE_OFN1539_n_10595;
wire FE_OFN1540_n_10595;
wire FE_OFN1541_n_10595;
wire FE_OFN1542_n_10566;
wire FE_OFN1543_n_10566;
wire FE_OFN1544_n_10566;
wire FE_OFN1545_n_10566;
wire FE_OFN1546_n_10566;
wire FE_OFN1547_n_10566;
wire FE_OFN1548_n_10566;
wire FE_OFN1549_n_12104;
wire FE_OFN1550_n_12104;
wire FE_OFN1551_n_12104;
wire FE_OFN1552_n_12104;
wire FE_OFN1553_n_12104;
wire FE_OFN1554_n_12104;
wire FE_OFN1556_n_12042;
wire FE_OFN1558_n_12042;
wire FE_OFN1559_n_12042;
wire FE_OFN1560_n_12502;
wire FE_OFN1561_n_12502;
wire FE_OFN1562_n_12502;
wire FE_OFN1563_n_12502;
wire FE_OFN1564_n_12502;
wire FE_OFN1565_n_12502;
wire FE_OFN1566_n_12502;
wire FE_OFN1568_n_11027;
wire FE_OFN1572_n_11027;
wire FE_OFN1573_n_12028;
wire FE_OFN1574_n_12028;
wire FE_OFN1575_n_12028;
wire FE_OFN1576_n_12028;
wire FE_OFN1577_n_12028;
wire FE_OFN1579_n_12306;
wire FE_OFN1581_n_12306;
wire FE_OFN1583_n_12306;
wire FE_OFN1584_n_12306;
wire FE_OFN1585_n_13736;
wire FE_OFN1586_n_13736;
wire FE_OFN1587_n_13736;
wire FE_OFN1588_n_13736;
wire FE_OFN1589_n_13736;
wire FE_OFN1590_n_13741;
wire FE_OFN1591_n_13741;
wire FE_OFN1592_n_13741;
wire FE_OFN1593_n_13741;
wire FE_OFN1596_n_13741;
wire FE_OFN1598_n_13995;
wire FE_OFN1599_n_13995;
wire FE_OFN1600_n_13995;
wire FE_OFN1601_n_13995;
wire FE_OFN1602_n_13995;
wire FE_OFN1603_n_13997;
wire FE_OFN1604_n_13997;
wire FE_OFN1605_n_13997;
wire FE_OFN1606_n_13997;
wire FE_OFN1607_n_2122;
wire FE_OFN1608_n_2122;
wire FE_OFN1609_n_2122;
wire FE_OFN1610_n_2122;
wire FE_OFN1611_n_2122;
wire FE_OFN1612_n_2122;
wire FE_OFN1613_n_1787;
wire FE_OFN1614_n_1787;
wire FE_OFN1615_n_1787;
wire FE_OFN1616_n_1787;
wire FE_OFN1617_n_1787;
wire FE_OFN1618_n_1787;
wire FE_OFN1619_n_1787;
wire FE_OFN1620_n_1787;
wire FE_OFN1621_n_1787;
wire FE_OFN1622_n_4438;
wire FE_OFN1623_n_4438;
wire FE_OFN1624_n_4438;
wire FE_OFN1625_n_4438;
wire FE_OFN1626_n_4438;
wire FE_OFN1627_n_4438;
wire FE_OFN1628_n_4438;
wire FE_OFN1629_n_9531;
wire FE_OFN1630_n_9531;
wire FE_OFN1631_n_9531;
wire FE_OFN1632_n_9531;
wire FE_OFN1633_n_9531;
wire FE_OFN1634_n_9531;
wire FE_OFN1635_n_9531;
wire FE_OFN1636_n_4460;
wire FE_OFN1637_n_4671;
wire FE_OFN1638_n_4671;
wire FE_OFN1639_n_4671;
wire FE_OFN1640_n_4671;
wire FE_OFN1641_n_4671;
wire FE_OFN1642_n_4671;
wire FE_OFN1643_n_4671;
wire FE_OFN1644_n_4671;
wire FE_OFN1645_n_4671;
wire FE_OFN1646_n_9428;
wire FE_OFN1647_n_9428;
wire FE_OFN1648_n_9428;
wire FE_OFN1649_n_9428;
wire FE_OFN1650_n_9428;
wire FE_OFN1651_n_9428;
wire FE_OFN1652_n_9502;
wire FE_OFN1653_n_9502;
wire FE_OFN1654_n_9502;
wire FE_OFN1655_n_9502;
wire FE_OFN1656_n_9502;
wire FE_OFN1657_n_9502;
wire FE_OFN1658_n_4490;
wire FE_OFN1659_n_4490;
wire FE_OFN1660_n_4490;
wire FE_OFN1661_n_4490;
wire FE_OFN1662_n_4490;
wire FE_OFN1663_n_4490;
wire FE_OFN1664_n_9477;
wire FE_OFN1665_n_9477;
wire FE_OFN1666_n_9477;
wire FE_OFN1667_n_9477;
wire FE_OFN1668_n_9477;
wire FE_OFN1669_n_9477;
wire FE_OFN1670_n_9477;
wire FE_OFN1671_n_9477;
wire FE_OFN1672_n_4655;
wire FE_OFN1673_n_4655;
wire FE_OFN1674_n_4655;
wire FE_OFN1675_n_4655;
wire FE_OFN1676_n_4655;
wire FE_OFN1677_n_4655;
wire FE_OFN1678_n_4655;
wire FE_OFN1679_n_4655;
wire FE_OFN1680_n_4655;
wire FE_OFN1681_n_4669;
wire FE_OFN1682_n_4669;
wire FE_OFN1683_n_9528;
wire FE_OFN1684_n_9528;
wire FE_OFN1685_n_9528;
wire FE_OFN1686_n_9528;
wire FE_OFN1687_n_9528;
wire FE_OFN1688_n_9528;
wire FE_OFN1689_n_9528;
wire FE_OFN1690_n_9528;
wire FE_OFN1691_n_9528;
wire FE_OFN1692_n_9528;
wire FE_OFN1693_n_3368;
wire FE_OFN1694_n_3368;
wire FE_OFN1695_n_3368;
wire FE_OFN1696_n_5751;
wire FE_OFN1697_n_5751;
wire FE_OFN1698_n_5751;
wire FE_OFN1699_n_5751;
wire FE_OFN1700_n_5751;
wire FE_OFN1701_n_4868;
wire FE_OFN1702_n_4868;
wire FE_OFN1703_n_4868;
wire FE_OFN1704_n_4868;
wire FE_OFN1705_n_4868;
wire FE_OFN1706_n_4868;
wire FE_OFN1707_n_4868;
wire FE_OFN1708_n_4868;
wire FE_OFN1709_n_4868;
wire FE_OFN1710_n_4868;
wire FE_OFN1711_n_13563;
wire FE_OFN1712_n_13563;
wire FE_OFN1713_n_13650;
wire FE_OFN1714_n_13650;
wire FE_OFN1716_n_16698;
wire FE_OFN1719_n_16891;
wire FE_OFN1720_n_16891;
wire FE_OFN1721_n_16891;
wire FE_OFN1722_n_16891;
wire FE_OFN1723_n_16891;
wire FE_OFN1724_n_16891;
wire FE_OFN1725_n_16891;
wire FE_OFN1726_n_9975;
wire FE_OFN1727_n_9975;
wire FE_OFN1728_n_9975;
wire FE_OFN1729_n_9975;
wire FE_OFN1730_n_9975;
wire FE_OFN1731_n_9975;
wire FE_OFN1732_n_16317;
wire FE_OFN1733_n_16317;
wire FE_OFN1734_n_16317;
wire FE_OFN1735_n_16317;
wire FE_OFN1736_n_16317;
wire FE_OFN1737_n_11019;
wire FE_OFN1738_n_11019;
wire FE_OFN1739_n_11019;
wire FE_OFN1740_n_11019;
wire FE_OFN1741_n_11019;
wire FE_OFN1742_n_11019;
wire FE_OFN1743_n_12004;
wire FE_OFN1744_n_12004;
wire FE_OFN1745_n_12004;
wire FE_OFN1746_n_12004;
wire FE_OFN1747_n_12004;
wire FE_OFN1748_n_12004;
wire FE_OFN1749_n_12004;
wire FE_OFN1751_n_12086;
wire FE_OFN1752_n_12086;
wire FE_OFN1753_n_12086;
wire FE_OFN1754_n_12681;
wire FE_OFN1755_n_12681;
wire FE_OFN1756_n_12681;
wire FE_OFN1757_n_12681;
wire FE_OFN1758_n_10780;
wire FE_OFN1759_n_10780;
wire FE_OFN1760_n_10780;
wire FE_OFN1761_n_10780;
wire FE_OFN1762_n_10780;
wire FE_OFN1767_n_14054;
wire FE_OFN1768_n_14054;
wire FE_OFN1769_n_14054;
wire FE_OFN1770_n_14054;
wire FE_OFN1771_n_14054;
wire FE_OFN1772_n_13800;
wire FE_OFN1773_n_13800;
wire FE_OFN1774_n_13800;
wire FE_OFN1775_n_13800;
wire FE_OFN1776_parchk_pci_ad_reg_in_1222;
wire FE_OFN1777_parchk_pci_ad_reg_in_1222;
wire FE_OFN1778_parchk_pci_ad_reg_in_1222;
wire FE_OFN1779_parchk_pci_ad_reg_in_1221;
wire FE_OFN1780_parchk_pci_ad_reg_in_1221;
wire FE_OFN1781_parchk_pci_ad_reg_in_1221;
wire FE_OFN1782_n_1699;
wire FE_OFN1783_n_1699;
wire FE_OFN1784_n_1699;
wire FE_OFN1785_n_1699;
wire FE_OFN1786_n_1699;
wire FE_OFN1789_n_9823;
wire FE_OFN1790_n_2687;
wire FE_OFN1791_n_9904;
wire FE_OFN1792_n_9904;
wire FE_OFN1793_n_9904;
wire FE_OFN1794_n_9904;
wire FE_OFN1795_n_9904;
wire FE_OFN1796_n_2299;
wire FE_OFN1797_n_2299;
wire FE_OFN1798_n_9690;
wire FE_OFN1799_n_9690;
wire FE_OFN1800_n_9690;
wire FE_OFN1801_n_9690;
wire FE_OFN1802_n_9690;
wire FE_OFN1803_n_9690;
wire FE_OFN1804_n_4501;
wire FE_OFN1805_n_4501;
wire FE_OFN1806_n_4501;
wire FE_OFN1807_n_4501;
wire FE_OFN1808_n_4454;
wire FE_OFN1809_n_4454;
wire FE_OFN1810_n_4454;
wire FE_OFN1811_n_7845;
wire FE_OFN1812_n_7845;
wire FE_OFN1813_n_2919;
wire FE_OFN1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid;
wire FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid;
wire FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid;
wire FE_OFN1819_n_2919;
wire FE_OFN186_n_15768;
wire FE_OFN190_n_1193;
wire FE_OFN191_n_1193;
wire FE_OFN1935_n_1781;
wire FE_OFN1936_n_1781;
wire FE_OFN1937_g66085_p;
wire FE_OFN1938_g66085_p;
wire FE_OFN1939_g66095_p;
wire FE_OFN1940_g66095_p;
wire FE_OFN1941_n_3241;
wire FE_OFN1942_n_3241;
wire FE_OFN1943_n_15813;
wire FE_OFN1944_n_15813;
wire FE_OFN1945_n_13784;
wire FE_OFN1946_n_13784;
wire FE_OFN196_n_2683;
wire FE_OFN197_n_2683;
wire FE_OFN198_n_3298;
wire FE_OFN199_n_3298;
wire FE_OFN1_n_4778;
wire FE_OFN200_n_9230;
wire FE_OFN201_n_9230;
wire FE_OFN2020_n_4778;
wire FE_OFN2021_n_4778;
wire FE_OFN2022_n_4778;
wire FE_OFN202_n_9228;
wire FE_OFN203_n_9228;
wire FE_OFN204_n_9140;
wire FE_OFN2051_n_6965;
wire FE_OFN2052_n_6965;
wire FE_OFN2053_n_8831;
wire FE_OFN2054_n_8831;
wire FE_OFN2055_n_8831;
wire FE_OFN2056_n_2117;
wire FE_OFN2057_n_2117;
wire FE_OFN2058_n_13447;
wire FE_OFN2059_n_13447;
wire FE_OFN205_n_9140;
wire FE_OFN2060_g66087_p;
wire FE_OFN2061_g66087_p;
wire FE_OFN2062_n_6391;
wire FE_OFN2063_n_6391;
wire FE_OFN2064_n_6391;
wire FE_OFN2069_n_15978;
wire FE_OFN206_n_9865;
wire FE_OFN2070_n_15978;
wire FE_OFN2071_n_15978;
wire FE_OFN2072_n_15978;
wire FE_OFN2073_n_2723;
wire FE_OFN2074_n_2723;
wire FE_OFN2075_FE_OCPUNCON1952_FE_OFN697_n_16760;
wire FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760;
wire FE_OFN2077_n_8069;
wire FE_OFN2079_n_8069;
wire FE_OFN207_n_9865;
wire FE_OFN2080_n_8176;
wire FE_OFN2081_n_8176;
wire FE_OFN2082_n_8407;
wire FE_OFN2083_n_8407;
wire FE_OFN2084_n_8407;
wire FE_OFN2085_n_8448;
wire FE_OFN2086_n_8448;
wire FE_OFN2088_n_13124;
wire FE_OFN208_n_9126;
wire FE_OFN2092_n_2301;
wire FE_OFN2093_n_2301;
wire FE_OFN2094_n_2520;
wire FE_OFN2095_n_2520;
wire FE_OFN2096_n_2520;
wire FE_OFN2099_n_3281;
wire FE_OFN209_n_9126;
wire FE_OFN2100_n_3281;
wire FE_OFN2101_n_2834;
wire FE_OFN2102_n_2834;
wire FE_OFN2103_g64577_p;
wire FE_OFN2104_g64577_p;
wire FE_OFN2105_g64577_p;
wire FE_OFN2106_g64577_p;
wire FE_OFN2107_n_2047;
wire FE_OFN2108_n_2047;
wire FE_OFN2109_n_2047;
wire FE_OFN210_n_9858;
wire FE_OFN2110_n_2248;
wire FE_OFN2111_n_2248;
wire FE_OFN2112_n_2053;
wire FE_OFN2113_n_2053;
wire FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source;
wire FE_OFN211_n_9858;
wire FE_OFN2121_n_2687;
wire FE_OFN2123_n_16497;
wire FE_OFN2124_n_16497;
wire FE_OFN2125_n_16497;
wire FE_OFN2126_n_16497;
wire FE_OFN2127_n_16497;
wire FE_OFN2128_n_16497;
wire FE_OFN2129_n_16720;
wire FE_OFN212_n_9124;
wire FE_OFN2130_n_10588;
wire FE_OFN2131_n_10588;
wire FE_OFN2132_n_13124;
wire FE_OFN2133_n_13124;
wire FE_OFN2134_n_13124;
wire FE_OFN2135_n_13124;
wire FE_OFN2136_n_13124;
wire FE_OFN2137_n_15534;
wire FE_OFN2139_n_16992;
wire FE_OFN213_n_9124;
wire FE_OFN2140_n_16992;
wire FE_OFN2141_n_16992;
wire FE_OFN2142_n_16992;
wire FE_OFN2143_n_16992;
wire FE_OFN2144_n_16992;
wire FE_OFN2145_n_16992;
wire FE_OFN2146_n_9320;
wire FE_OFN2147_n_10595;
wire FE_OFN2148_n_10595;
wire FE_OFN2149_n_10595;
wire FE_OFN214_n_9856;
wire FE_OFN2150_n_10595;
wire FE_OFN2151_n_16439;
wire FE_OFN2152_n_16439;
wire FE_OFN2153_n_16439;
wire FE_OFN2154_n_16439;
wire FE_OFN2155_n_16439;
wire FE_OFN2156_n_16439;
wire FE_OFN2157_n_16439;
wire FE_OFN2158_n_16439;
wire FE_OFN2159_n_16301;
wire FE_OFN215_n_9856;
wire FE_OFN2160_n_16301;
wire FE_OFN2161_n_16301;
wire FE_OFN2162_n_16301;
wire FE_OFN2163_n_16301;
wire FE_OFN2164_n_16301;
wire FE_OFN2165_n_16301;
wire FE_OFN2166_n_8567;
wire FE_OFN2167_n_8567;
wire FE_OFN2168_n_8567;
wire FE_OFN2169_n_8567;
wire FE_OFN216_n_9889;
wire FE_OFN2170_n_8567;
wire FE_OFN2171_n_8567;
wire FE_OFN2172_n_8567;
wire FE_OFN2173_n_8567;
wire FE_OFN2174_n_8567;
wire FE_OFN2175_n_8567;
wire FE_OFN2176_n_8567;
wire FE_OFN2177_n_8567;
wire FE_OFN2178_n_8567;
wire FE_OFN2179_n_8567;
wire FE_OFN217_n_9889;
wire FE_OFN2180_n_8567;
wire FE_OFN2181_n_8567;
wire FE_OFN2182_n_8567;
wire FE_OFN2183_n_8567;
wire FE_OFN2184_n_8567;
wire FE_OFN2185_n_8567;
wire FE_OFN2186_n_8567;
wire FE_OFN2187_n_8567;
wire FE_OFN2188_n_8567;
wire FE_OFN2189_n_8567;
wire FE_OFN218_n_9853;
wire FE_OFN2190_n_8567;
wire FE_OFN2191_n_8567;
wire FE_OFN2192_n_16779;
wire FE_OFN2193_n_9163;
wire FE_OFN2194_n_9163;
wire FE_OFN2195_n_9163;
wire FE_OFN2196_n_9163;
wire FE_OFN2197_n_10256;
wire FE_OFN2198_n_10256;
wire FE_OFN2199_n_10256;
wire FE_OFN219_n_9853;
wire FE_OFN21_n_9372;
wire FE_OFN2200_n_10256;
wire FE_OFN2201_n_12042;
wire FE_OFN2202_n_12042;
wire FE_OFN2203_n_12042;
wire FE_OFN2204_n_12028;
wire FE_OFN2205_n_10538;
wire FE_OFN2206_n_10892;
wire FE_OFN2207_n_10892;
wire FE_OFN2208_n_11795;
wire FE_OFN2209_n_11027;
wire FE_OFN220_n_9846;
wire FE_OFN2210_n_11027;
wire FE_OFN2211_n_8407;
wire FE_OFN2212_n_8407;
wire FE_OFN2213_n_15366;
wire FE_OFN2214_n_15366;
wire FE_OFN2215_n_15366;
wire FE_OFN2216_n_10143;
wire FE_OFN221_n_9846;
wire FE_OFN222_n_9844;
wire FE_OFN223_n_9844;
wire FE_OFN2240_g52675_p;
wire FE_OFN2241_g52675_p;
wire FE_OFN2242_g52675_p;
wire FE_OFN2243_g52675_p;
wire FE_OFN2244_n_4792;
wire FE_OFN2245_n_4792;
wire FE_OFN2246_n_2113;
wire FE_OFN2247_n_2113;
wire FE_OFN2248_n_1790;
wire FE_OFN2249_n_1790;
wire FE_OFN224_n_9122;
wire FE_OFN2250_n_2101;
wire FE_OFN2251_n_2101;
wire FE_OFN2252_n_9687;
wire FE_OFN2253_n_9687;
wire FE_OFN2254_n_9687;
wire FE_OFN2255_n_8060;
wire FE_OFN2256_n_8060;
wire FE_OFN2257_n_8060;
wire FE_OFN2258_n_8060;
wire FE_OFN2259_n_2775;
wire FE_OFN225_n_9122;
wire FE_OFN2260_n_2775;
wire FE_OFN226_n_9841;
wire FE_OFN227_n_9841;
wire FE_OFN228_n_9120;
wire FE_OFN229_n_9120;
wire FE_OFN230_n_9839;
wire FE_OFN231_n_9839;
wire FE_OFN232_n_9876;
wire FE_OFN233_n_9876;
wire FE_OFN234_n_9834;
wire FE_OFN235_n_9834;
wire FE_OFN236_n_9118;
wire FE_OFN237_n_9118;
wire FE_OFN238_n_9832;
wire FE_OFN239_n_9832;
wire FE_OFN240_n_9830;
wire FE_OFN241_n_9830;
wire FE_OFN242_n_9116;
wire FE_OFN243_n_9116;
wire FE_OFN244_n_9114;
wire FE_OFN245_n_9114;
wire FE_OFN246_n_9112;
wire FE_OFN247_n_9112;
wire FE_OFN248_n_9789;
wire FE_OFN250_n_9789;
wire FE_OFN251_n_9868;
wire FE_OFN252_n_9868;
wire FE_OFN253_n_9825;
wire FE_OFN254_n_9825;
wire FE_OFN255_n_8969;
wire FE_OFN256_n_8969;
wire FE_OFN257_n_9862;
wire FE_OFN258_n_9862;
wire FE_OFN259_n_9860;
wire FE_OFN260_n_9860;
wire FE_OFN261_n_9851;
wire FE_OFN262_n_9851;
wire FE_OFN263_n_9849;
wire FE_OFN264_n_9849;
wire FE_OFN265_n_9884;
wire FE_OFN266_n_9884;
wire FE_OFN267_n_9880;
wire FE_OFN268_n_9880;
wire FE_OFN269_n_9836;
wire FE_OFN270_n_9836;
wire FE_OFN271_n_9828;
wire FE_OFN272_n_9828;
wire FE_OFN275_n_9941;
wire FE_OFN276_n_9941;
wire FE_OFN2_n_4778;
wire FE_OFN334_g66081_p;
wire FE_OFN335_g66081_p;
wire FE_OFN336_g66089_p;
wire FE_OFN337_g66089_p;
wire FE_OFN365_n_4093;
wire FE_OFN369_n_4092;
wire FE_OFN3_n_4778;
wire FE_OFN514_n_9697;
wire FE_OFN515_n_9697;
wire FE_OFN516_n_9697;
wire FE_OFN517_n_9697;
wire FE_OFN518_n_9697;
wire FE_OFN519_n_9697;
wire FE_OFN523_n_9428;
wire FE_OFN524_n_9899;
wire FE_OFN525_n_9899;
wire FE_OFN526_n_9899;
wire FE_OFN527_n_9899;
wire FE_OFN528_n_9899;
wire FE_OFN529_n_9899;
wire FE_OFN530_n_9823;
wire FE_OFN531_n_9823;
wire FE_OFN532_n_9823;
wire FE_OFN533_n_9823;
wire FE_OFN534_n_9823;
wire FE_OFN535_n_9823;
wire FE_OFN537_n_9690;
wire FE_OFN539_n_9690;
wire FE_OFN540_n_9690;
wire FE_OFN541_n_9690;
wire FE_OFN542_n_9690;
wire FE_OFN543_n_9690;
wire FE_OFN548_n_9477;
wire FE_OFN549_n_9864;
wire FE_OFN550_n_9864;
wire FE_OFN551_n_9864;
wire FE_OFN552_n_9864;
wire FE_OFN553_n_9864;
wire FE_OFN554_n_9864;
wire FE_OFN555_n_9864;
wire FE_OFN556_n_9864;
wire FE_OFN557_n_9895;
wire FE_OFN558_n_9895;
wire FE_OFN559_n_9895;
wire FE_OFN560_n_9895;
wire FE_OFN561_n_9895;
wire FE_OFN562_n_9895;
wire FE_OFN563_n_9895;
wire FE_OFN564_n_9895;
wire FE_OFN568_n_9528;
wire FE_OFN569_n_9528;
wire FE_OFN572_n_9502;
wire FE_OFN573_n_9902;
wire FE_OFN574_n_9902;
wire FE_OFN575_n_9902;
wire FE_OFN576_n_9902;
wire FE_OFN577_n_9902;
wire FE_OFN579_n_9531;
wire FE_OFN580_n_9531;
wire FE_OFN582_n_9692;
wire FE_OFN583_n_9692;
wire FE_OFN584_n_9692;
wire FE_OFN585_n_9692;
wire FE_OFN587_n_9692;
wire FE_OFN588_n_9692;
wire FE_OFN589_n_9692;
wire FE_OFN590_n_9694;
wire FE_OFN591_n_9694;
wire FE_OFN592_n_9694;
wire FE_OFN593_n_9694;
wire FE_OFN595_n_9694;
wire FE_OFN596_n_9694;
wire FE_OFN597_n_9694;
wire FE_OFN598_n_9687;
wire FE_OFN599_n_9687;
wire FE_OFN600_n_9687;
wire FE_OFN601_n_9687;
wire FE_OFN602_n_9687;
wire FE_OFN603_n_9687;
wire FE_OFN605_n_9904;
wire FE_OFN606_n_9904;
wire FE_OFN607_n_9904;
wire FE_OFN608_n_9904;
wire FE_OFN611_n_4501;
wire FE_OFN612_n_4501;
wire FE_OFN613_n_4501;
wire FE_OFN614_n_4501;
wire FE_OFN615_n_4501;
wire FE_OFN618_n_4490;
wire FE_OFN619_n_4490;
wire FE_OFN620_n_4490;
wire FE_OFN621_n_4409;
wire FE_OFN622_n_4409;
wire FE_OFN623_n_4409;
wire FE_OFN624_n_4409;
wire FE_OFN625_n_4409;
wire FE_OFN627_n_4454;
wire FE_OFN628_n_4454;
wire FE_OFN629_n_4454;
wire FE_OFN630_n_4454;
wire FE_OFN631_n_4454;
wire FE_OFN632_n_4454;
wire FE_OFN633_n_4454;
wire FE_OFN634_n_4454;
wire FE_OFN636_n_4669;
wire FE_OFN638_n_4669;
wire FE_OFN639_n_4669;
wire FE_OFN640_n_4669;
wire FE_OFN641_n_4677;
wire FE_OFN642_n_4677;
wire FE_OFN643_n_4677;
wire FE_OFN644_n_4677;
wire FE_OFN645_n_4497;
wire FE_OFN646_n_4497;
wire FE_OFN647_n_4497;
wire FE_OFN648_n_4497;
wire FE_OFN649_n_4497;
wire FE_OFN650_n_4508;
wire FE_OFN651_n_4508;
wire FE_OFN652_n_4508;
wire FE_OFN653_n_4508;
wire FE_OFN654_n_4508;
wire FE_OFN658_n_4392;
wire FE_OFN659_n_4392;
wire FE_OFN660_n_4392;
wire FE_OFN661_n_4392;
wire FE_OFN662_n_4392;
wire FE_OFN663_n_4495;
wire FE_OFN664_n_4495;
wire FE_OFN665_n_4495;
wire FE_OFN666_n_4495;
wire FE_OFN667_n_4495;
wire FE_OFN668_n_4505;
wire FE_OFN669_n_4505;
wire FE_OFN670_n_4505;
wire FE_OFN671_n_4505;
wire FE_OFN672_n_4505;
wire FE_OFN678_n_4460;
wire FE_OFN679_n_4460;
wire FE_OFN681_n_4460;
wire FE_OFN682_n_4460;
wire FE_OFN683_n_4417;
wire FE_OFN684_n_4417;
wire FE_OFN685_n_4417;
wire FE_OFN686_n_4417;
wire FE_OFN687_n_4417;
wire FE_OFN689_n_4438;
wire FE_OFN697_n_16760;
wire FE_OFN698_n_7845;
wire FE_OFN699_n_7845;
wire FE_OFN700_n_7845;
wire FE_OFN701_n_7845;
wire FE_OFN702_n_7845;
wire FE_OFN703_n_8069;
wire FE_OFN704_n_8069;
wire FE_OFN705_n_8119;
wire FE_OFN706_n_8119;
wire FE_OFN707_n_8119;
wire FE_OFN708_n_8232;
wire FE_OFN709_n_8232;
wire FE_OFN710_n_8232;
wire FE_OFN711_n_8140;
wire FE_OFN712_n_8140;
wire FE_OFN713_n_8140;
wire FE_OFN714_n_8140;
wire FE_OFN715_n_8176;
wire FE_OFN716_n_8176;
wire FE_OFN717_n_8176;
wire FE_OFN718_n_8060;
wire FE_OFN719_n_8060;
wire FE_OFN720_n_8060;
wire FE_OFN732_n_7498;
wire FE_OFN775_n_15366;
wire FE_OFN776_n_15366;
wire FE_OFN777_n_4152;
wire FE_OFN778_n_4152;
wire FE_OFN779_n_2746;
wire FE_OFN780_n_2746;
wire FE_OFN781_n_2746;
wire FE_OFN782_n_2678;
wire FE_OFN783_n_2678;
wire FE_OFN784_n_2678;
wire FE_OFN785_n_2678;
wire FE_OFN786_n_2678;
wire FE_OFN787_n_2678;
wire FE_OFN789_n_2678;
wire FE_OFN792_n_2547;
wire FE_OFN793_n_2547;
wire FE_OFN794_n_2520;
wire FE_OFN795_n_2520;
wire FE_OFN877_g64577_p;
wire FE_OFN881_g64577_p;
wire FE_OFN882_g64577_p;
wire FE_OFN8_n_11877;
wire FE_OFN900_n_4736;
wire FE_OFN901_n_4736;
wire FE_OFN902_n_4736;
wire FE_OFN903_n_4736;
wire FE_OFN904_n_4736;
wire FE_OFN905_n_4736;
wire FE_OFN906_n_4736;
wire FE_OFN908_n_4734;
wire FE_OFN912_n_4727;
wire FE_OFN915_n_4725;
wire FE_OFN916_n_4725;
wire FE_OFN917_n_4725;
wire FE_OFN918_n_4725;
wire FE_OFN923_n_4740;
wire FE_OFN926_n_4730;
wire FE_OFN927_n_4730;
wire FE_OFN928_n_4730;
wire FE_OFN929_n_4730;
wire FE_OFN930_n_4730;
wire FE_OFN934_n_2292;
wire FE_OFN935_n_2292;
wire FE_OFN936_n_2292;
wire FE_OFN937_n_2292;
wire FE_OFN938_n_2292;
wire FE_OFN941_n_2047;
wire FE_OFN944_n_2248;
wire FE_OFN945_n_2248;
wire FE_OFN946_n_2248;
wire FE_OFN947_n_2248;
wire FE_OFN948_n_2248;
wire FE_OFN949_n_2055;
wire FE_OFN950_n_2055;
wire FE_OFN951_n_2055;
wire FE_OFN952_n_2055;
wire FE_OFN953_n_2055;
wire FE_OFN954_n_1699;
wire FE_OFN955_n_1699;
wire FE_OFN956_n_1699;
wire FE_OFN957_n_2299;
wire FE_OFN958_n_2299;
wire FE_OFN959_n_2299;
wire FE_OFN966_n_2233;
wire FE_OFN967_n_2233;
wire FE_OFN968_n_13784;
wire FE_OFN969_n_13784;
wire FE_OFN982_n_2700;
wire FE_OFN983_n_2700;
wire FE_OFN984_n_2697;
wire FE_OFN985_n_2697;
wire FE_OFN986_n_2696;
wire FE_OFN987_n_2696;
wire FE_OFN988_n_574;
wire FE_OFN989_n_574;
wire FE_OFN991_n_2373;
wire FE_OFN992_n_2373;
wire FE_OFN993_n_15366;
wire FE_OFN994_n_15366;
wire FE_OFN995_n_15366;
wire FE_OFN996_n_15366;
wire FE_OFN997_n_15978;
wire FE_OFN999_n_15978;
wire FE_OFN9_n_11877;
wire FE_RN_0_0;
wire FE_RN_100_0;
wire FE_RN_101_0;
wire FE_RN_102_0;
wire FE_RN_103_0;
wire FE_RN_105_0;
wire FE_RN_106_0;
wire FE_RN_107_0;
wire FE_RN_108_0;
wire FE_RN_109_0;
wire FE_RN_110_0;
wire FE_RN_111_0;
wire FE_RN_112_0;
wire FE_RN_113_0;
wire FE_RN_114_0;
wire FE_RN_115_0;
wire FE_RN_116_0;
wire TIMEBOOST_net_184;
wire FE_RN_120_0;
wire FE_RN_121_0;
wire FE_RN_122_0;
wire FE_RN_124_0;
wire TIMEBOOST_net_17013;
wire FE_RN_127_0;
wire TIMEBOOST_net_10415;
wire FE_RN_130_0;
wire TIMEBOOST_net_10414;
wire FE_RN_135_0;
wire FE_RN_136_0;
wire FE_RN_137_0;
wire FE_RN_138_0;
wire FE_RN_139_0;
wire FE_RN_140_0;
wire FE_RN_141_0;
wire FE_RN_142_0;
wire FE_RN_143_0;
wire FE_RN_144_0;
wire FE_RN_145_0;
wire FE_RN_146_0;
wire FE_RN_147_0;
wire FE_RN_148_0;
wire FE_RN_149_0;
wire FE_RN_150_0;
wire FE_RN_151_0;
wire TIMEBOOST_net_340;
wire FE_RN_153_0;
wire FE_RN_154_0;
wire TIMEBOOST_net_17276;
wire FE_RN_156_0;
wire FE_RN_158_0;
wire FE_RN_159_0;
wire FE_RN_15_0;
wire FE_RN_160_0;
wire TIMEBOOST_net_12480;
wire TIMEBOOST_net_23266;
wire FE_RN_176_0;
wire FE_RN_177_0;
wire FE_RN_178_0;
wire FE_RN_179_0;
wire FE_RN_180_0;
wire FE_RN_181_0;
wire FE_RN_182_0;
wire FE_RN_183_0;
wire FE_RN_184_0;
wire FE_RN_185_0;
wire FE_RN_186_0;
wire FE_RN_187_0;
wire FE_RN_188_0;
wire FE_RN_189_0;
wire FE_RN_18_0;
wire FE_RN_190_0;
wire FE_RN_191_0;
wire FE_RN_192_0;
wire FE_RN_193_0;
wire FE_RN_194_0;
wire FE_RN_195_0;
wire FE_RN_196_0;
wire FE_RN_197_0;
wire FE_RN_198_0;
wire FE_RN_199_0;
wire FE_RN_19_0;
wire FE_RN_200_0;
wire FE_RN_201_0;
wire FE_RN_202_0;
wire FE_RN_203_0;
wire FE_RN_207_0;
wire FE_RN_208_0;
wire FE_RN_209_0;
wire FE_RN_20_0;
wire FE_RN_211_0;
wire FE_RN_213_0;
wire FE_RN_214_0;
wire FE_RN_215_0;
wire FE_RN_216_0;
wire FE_RN_217_0;
wire FE_RN_218_0;
wire FE_RN_219_0;
wire FE_RN_220_0;
wire FE_RN_221_0;
wire FE_RN_222_0;
wire FE_RN_223_0;
wire FE_RN_224_0;
wire FE_RN_225_0;
wire FE_RN_226_0;
wire FE_RN_227_0;
wire FE_RN_228_0;
wire FE_RN_229_0;
wire FE_RN_230_0;
wire FE_RN_231_0;
wire FE_RN_232_0;
wire FE_RN_233_0;
wire FE_RN_234_0;
wire FE_RN_235_0;
wire FE_RN_236_0;
wire FE_RN_237_0;
wire FE_RN_238_0;
wire TIMEBOOST_net_12597;
wire FE_RN_23_0;
wire FE_RN_240_0;
wire FE_RN_241_0;
wire FE_RN_243_0;
wire FE_RN_244_0;
wire FE_RN_246_0;
wire FE_RN_247_0;
wire TIMEBOOST_net_13790;
wire FE_RN_249_0;
wire FE_RN_250_0;
wire FE_RN_251_0;
wire FE_RN_259_0;
wire FE_RN_25_0;
wire FE_RN_260_0;
wire FE_RN_261_0;
wire FE_RN_262_0;
wire FE_RN_263_0;
wire FE_RN_264_0;
wire TIMEBOOST_net_10599;
wire TIMEBOOST_net_20745;
wire FE_RN_267_0;
wire FE_RN_268_0;
wire FE_RN_269_0;
wire FE_RN_26_0;
wire FE_RN_270_0;
wire FE_RN_271_0;
wire TIMEBOOST_net_10435;
wire FE_RN_273_0;
wire FE_RN_274_0;
wire FE_RN_275_0;
wire FE_RN_276_0;
wire FE_RN_278_0;
wire FE_RN_279_0;
wire FE_RN_27_0;
wire FE_RN_280_0;
wire FE_RN_281_0;
wire TIMEBOOST_net_16382;
wire FE_RN_284_0;
wire FE_RN_285_0;
wire TIMEBOOST_net_10048;
wire FE_RN_28_0;
wire FE_RN_294_0;
wire FE_RN_295_0;
wire TIMEBOOST_net_6;
wire FE_RN_299_0;
wire FE_RN_29_0;
wire TIMEBOOST_net_16743;
wire FE_RN_303_0;
wire FE_RN_304_0;
wire FE_RN_305_0;
wire FE_RN_307_0;
wire FE_RN_308_0;
wire FE_RN_309_0;
wire FE_RN_30_0;
wire FE_RN_310_0;
wire FE_RN_311_0;
wire FE_RN_312_0;
wire FE_RN_313_0;
wire FE_RN_314_0;
wire FE_RN_315_0;
wire FE_RN_316_0;
wire FE_RN_317_0;
wire FE_RN_318_0;
wire FE_RN_319_0;
wire FE_RN_31_0;
wire FE_RN_320_0;
wire FE_RN_321_0;
wire FE_RN_322_0;
wire FE_RN_323_0;
wire FE_RN_324_0;
wire FE_RN_325_0;
wire FE_RN_326_0;
wire FE_RN_327_0;
wire FE_RN_328_0;
wire FE_RN_329_0;
wire FE_RN_32_0;
wire FE_RN_330_0;
wire FE_RN_331_0;
wire FE_RN_332_0;
wire FE_RN_333_0;
wire FE_RN_334_0;
wire FE_RN_335_0;
wire FE_RN_336_0;
wire FE_RN_337_0;
wire FE_RN_338_0;
wire FE_RN_339_0;
wire FE_RN_33_0;
wire FE_RN_340_0;
wire FE_RN_341_0;
wire FE_RN_342_0;
wire FE_RN_343_0;
wire FE_RN_344_0;
wire FE_RN_345_0;
wire FE_RN_346_0;
wire FE_RN_347_0;
wire FE_RN_348_0;
wire FE_RN_349_0;
wire FE_RN_34_0;
wire FE_RN_350_0;
wire FE_RN_351_0;
wire FE_RN_352_0;
wire FE_RN_353_0;
wire FE_RN_354_0;
wire FE_RN_355_0;
wire FE_RN_356_0;
wire FE_RN_357_0;
wire FE_RN_358_0;
wire FE_RN_359_0;
wire FE_RN_35_0;
wire FE_RN_360_0;
wire FE_RN_361_0;
wire FE_RN_362_0;
wire TIMEBOOST_net_10137;
wire FE_RN_365_0;
wire FE_RN_366_0;
wire FE_RN_368_0;
wire FE_RN_369_0;
wire FE_RN_36_0;
wire FE_RN_370_0;
wire FE_RN_371_0;
wire TIMEBOOST_net_5477;
wire FE_RN_373_0;
wire FE_RN_374_0;
wire TIMEBOOST_net_5478;
wire FE_RN_376_0;
wire FE_RN_377_0;
wire FE_RN_37_0;
wire FE_RN_381_0;
wire FE_RN_382_0;
wire FE_RN_383_0;
wire FE_RN_384_0;
wire FE_RN_385_0;
wire FE_RN_386_0;
wire FE_RN_387_0;
wire FE_RN_388_0;
wire FE_RN_389_0;
wire FE_RN_390_0;
wire FE_RN_392_0;
wire FE_RN_393_0;
wire FE_RN_394_0;
wire FE_RN_395_0;
wire FE_RN_396_0;
wire FE_RN_397_0;
wire FE_RN_398_0;
wire FE_RN_399_0;
wire FE_RN_39_0;
wire FE_RN_400_0;
wire FE_RN_401_0;
wire FE_RN_402_0;
wire FE_RN_403_0;
wire FE_RN_404_0;
wire FE_RN_405_0;
wire FE_RN_406_0;
wire FE_RN_407_0;
wire FE_RN_409_0;
wire FE_RN_40_0;
wire FE_RN_410_0;
wire FE_RN_415_0;
wire FE_RN_416_0;
wire FE_RN_417_0;
wire FE_RN_418_0;
wire FE_RN_419_0;
wire FE_RN_41_0;
wire FE_RN_420_0;
wire FE_RN_421_0;
wire FE_RN_422_0;
wire FE_RN_423_0;
wire TIMEBOOST_net_20381;
wire FE_RN_425_0;
wire FE_RN_426_0;
wire FE_RN_427_0;
wire FE_RN_428_0;
wire FE_RN_429_0;
wire FE_RN_42_0;
wire FE_RN_430_0;
wire FE_RN_431_0;
wire FE_RN_432_0;
wire FE_RN_433_0;
wire FE_RN_434_0;
wire TIMEBOOST_net_16489;
wire FE_RN_437_0;
wire FE_RN_438_0;
wire FE_RN_439_0;
wire FE_RN_43_0;
wire FE_RN_440_0;
wire FE_RN_441_0;
wire FE_RN_442_0;
wire FE_RN_443_0;
wire FE_RN_444_0;
wire FE_RN_445_0;
wire FE_RN_446_0;
wire FE_RN_447_0;
wire FE_RN_448_0;
wire FE_RN_449_0;
wire FE_RN_44_0;
wire FE_RN_450_0;
wire FE_RN_452_0;
wire FE_RN_453_0;
wire FE_RN_454_0;
wire TIMEBOOST_net_13695;
wire FE_RN_456_0;
wire FE_RN_457_0;
wire FE_RN_458_0;
wire FE_RN_459_0;
wire FE_RN_45_0;
wire FE_RN_460_0;
wire FE_RN_462_0;
wire FE_RN_463_0;
wire FE_RN_464_0;
wire FE_RN_465_0;
wire FE_RN_466_0;
wire FE_RN_467_0;
wire FE_RN_468_0;
wire FE_RN_469_0;
wire FE_RN_46_0;
wire FE_RN_470_0;
wire FE_RN_471_0;
wire FE_RN_472_0;
wire FE_RN_473_0;
wire FE_RN_474_0;
wire FE_RN_475_0;
wire FE_RN_476_0;
wire FE_RN_477_0;
wire FE_RN_478_0;
wire FE_RN_479_0;
wire FE_RN_47_0;
wire FE_RN_480_0;
wire FE_RN_481_0;
wire FE_RN_483_0;
wire FE_RN_484_0;
wire FE_RN_489_0;
wire FE_RN_48_0;
wire FE_RN_490_0;
wire FE_RN_491_0;
wire FE_RN_493_0;
wire FE_RN_494_0;
wire TIMEBOOST_net_16810;
wire FE_RN_496_0;
wire TIMEBOOST_net_21462;
wire FE_RN_498_0;
wire FE_RN_49_0;
wire FE_RN_500_0;
wire FE_RN_501_0;
wire FE_RN_502_0;
wire FE_RN_503_0;
wire TIMEBOOST_net_13592;
wire FE_RN_506_0;
wire FE_RN_507_0;
wire FE_RN_508_0;
wire FE_RN_509_0;
wire TIMEBOOST_net_10067;
wire FE_RN_510_0;
wire FE_RN_511_0;
wire FE_RN_512_0;
wire FE_RN_513_0;
wire FE_RN_514_0;
wire FE_RN_515_0;
wire FE_RN_516_0;
wire FE_RN_517_0;
wire FE_RN_518_0;
wire FE_RN_519_0;
wire FE_RN_51_0;
wire FE_RN_520_0;
wire FE_RN_521_0;
wire FE_RN_522_0;
wire FE_RN_523_0;
wire FE_RN_524_0;
wire FE_RN_525_0;
wire FE_RN_526_0;
wire FE_RN_527_0;
wire FE_RN_528_0;
wire FE_RN_529_0;
wire FE_RN_52_0;
wire FE_RN_530_0;
wire FE_RN_531_0;
wire FE_RN_532_0;
wire FE_RN_533_0;
wire TIMEBOOST_net_21753;
wire FE_RN_535_0;
wire TIMEBOOST_net_8791;
wire FE_RN_538_0;
wire FE_RN_539_0;
wire FE_RN_53_0;
wire FE_RN_541_0;
wire FE_RN_542_0;
wire TIMEBOOST_net_5482;
wire FE_RN_544_0;
wire FE_RN_545_0;
wire TIMEBOOST_net_9481;
wire FE_RN_547_0;
wire FE_RN_548_0;
wire FE_RN_549_0;
wire TIMEBOOST_net_7;
wire FE_RN_551_0;
wire FE_RN_552_0;
wire FE_RN_553_0;
wire FE_RN_554_0;
wire FE_RN_555_0;
wire FE_RN_556_0;
wire FE_RN_557_0;
wire FE_RN_558_0;
wire FE_RN_559_0;
wire FE_RN_55_0;
wire FE_RN_560_0;
wire FE_RN_561_0;
wire FE_RN_562_0;
wire TIMEBOOST_net_8823;
wire FE_RN_564_0;
wire FE_RN_565_0;
wire FE_RN_566_0;
wire FE_RN_567_0;
wire FE_RN_569_0;
wire FE_RN_56_0;
wire FE_RN_570_0;
wire FE_RN_571_0;
wire g66401_db;
wire FE_RN_573_0;
wire TIMEBOOST_net_22248;
wire TIMEBOOST_net_16724;
wire FE_RN_577_0;
wire FE_RN_578_0;
wire TIMEBOOST_net_22418;
wire FE_RN_57_0;
wire FE_RN_580_0;
wire FE_RN_581_0;
wire FE_RN_582_0;
wire FE_RN_583_0;
wire FE_RN_584_0;
wire TIMEBOOST_net_16798;
wire TIMEBOOST_net_13752;
wire TIMEBOOST_net_20388;
wire FE_RN_589_0;
wire FE_RN_58_0;
wire FE_RN_590_0;
wire FE_RN_591_0;
wire FE_RN_592_0;
wire FE_RN_593_0;
wire FE_RN_594_0;
wire FE_RN_595_0;
wire FE_RN_596_0;
wire FE_RN_597_0;
wire FE_RN_598_0;
wire TIMEBOOST_net_23018;
wire TIMEBOOST_net_13711;
wire FE_RN_601_0;
wire FE_RN_602_0;
wire FE_RN_603_0;
wire FE_RN_604_0;
wire FE_RN_605_0;
wire FE_RN_606_0;
wire FE_RN_607_0;
wire FE_RN_608_0;
wire FE_RN_609_0;
wire FE_RN_60_0;
wire FE_RN_610_0;
wire FE_RN_611_0;
wire FE_RN_612_0;
wire FE_RN_613_0;
wire FE_RN_614_0;
wire FE_RN_615_0;
wire FE_RN_616_0;
wire FE_RN_617_0;
wire FE_RN_618_0;
wire FE_RN_619_0;
wire FE_RN_61_0;
wire FE_RN_620_0;
wire FE_RN_621_0;
wire FE_RN_622_0;
wire FE_RN_623_0;
wire TIMEBOOST_net_14495;
wire TIMEBOOST_net_14544;
wire FE_RN_626_0;
wire FE_RN_627_0;
wire FE_RN_628_0;
wire TIMEBOOST_net_16169;
wire TIMEBOOST_net_23256;
wire TIMEBOOST_net_13664;
wire FE_RN_631_0;
wire FE_RN_632_0;
wire FE_RN_633_0;
wire TIMEBOOST_net_17452;
wire FE_RN_636_0;
wire FE_RN_637_0;
wire FE_RN_638_0;
wire TIMEBOOST_net_16652;
wire FE_RN_63_0;
wire FE_RN_641_0;
wire FE_RN_642_0;
wire FE_RN_643_0;
wire FE_RN_644_0;
wire FE_RN_645_0;
wire FE_RN_646_0;
wire FE_RN_647_0;
wire FE_RN_648_0;
wire FE_RN_649_0;
wire FE_RN_64_0;
wire FE_RN_650_0;
wire FE_RN_651_0;
wire FE_RN_653_0;
wire FE_RN_654_0;
wire FE_RN_655_0;
wire FE_RN_656_0;
wire FE_RN_657_0;
wire FE_RN_659_0;
wire TIMEBOOST_net_17103;
wire FE_RN_660_0;
wire FE_RN_661_0;
wire FE_RN_662_0;
wire FE_RN_663_0;
wire FE_RN_665_0;
wire FE_RN_666_0;
wire FE_RN_667_0;
wire FE_RN_668_0;
wire FE_RN_669_0;
wire FE_RN_66_0;
wire FE_RN_670_0;
wire FE_RN_672_0;
wire FE_RN_673_0;
wire FE_RN_674_0;
wire FE_RN_675_0;
wire TIMEBOOST_net_32;
wire FE_RN_677_0;
wire FE_RN_678_0;
wire TIMEBOOST_net_14564;
wire FE_RN_67_0;
wire FE_RN_680_0;
wire FE_RN_681_0;
wire FE_RN_682_0;
wire FE_RN_683_0;
wire FE_RN_684_0;
wire FE_RN_685_0;
wire FE_RN_686_0;
wire TIMEBOOST_net_20201;
wire FE_RN_688_0;
wire FE_RN_689_0;
wire FE_RN_691_0;
wire FE_RN_693_0;
wire FE_RN_694_0;
wire FE_RN_695_0;
wire FE_RN_697_0;
wire FE_RN_698_0;
wire FE_RN_699_0;
wire FE_RN_69_0;
wire FE_RN_6_0;
wire FE_RN_700_0;
wire FE_RN_701_0;
wire FE_RN_702_0;
wire FE_RN_703_0;
wire FE_RN_704_0;
wire FE_RN_705_0;
wire TIMEBOOST_net_11501;
wire TIMEBOOST_net_17109;
wire FE_RN_708_0;
wire FE_RN_709_0;
wire FE_RN_70_0;
wire FE_RN_710_0;
wire FE_RN_711_0;
wire TIMEBOOST_net_5476;
wire FE_RN_713_0;
wire FE_RN_714_0;
wire FE_RN_715_0;
wire FE_RN_716_0;
wire FE_RN_717_0;
wire FE_RN_71_0;
wire FE_RN_720_0;
wire FE_RN_722_0;
wire FE_RN_723_0;
wire FE_RN_725_0;
wire FE_RN_726_0;
wire TIMEBOOST_net_22794;
wire FE_RN_728_0;
wire FE_RN_729_0;
wire FE_RN_72_0;
wire TIMEBOOST_net_14323;
wire FE_RN_731_0;
wire FE_RN_732_0;
wire FE_RN_734_0;
wire FE_RN_735_0;
wire FE_RN_737_0;
wire FE_RN_738_0;
wire FE_RN_739_0;
wire FE_RN_73_0;
wire FE_RN_740_0;
wire FE_RN_741_0;
wire FE_RN_743_0;
wire FE_RN_744_0;
wire FE_RN_745_0;
wire FE_RN_746_0;
wire FE_RN_747_0;
wire FE_RN_748_0;
wire FE_RN_749_0;
wire TIMEBOOST_net_22881;
wire FE_RN_750_0;
wire FE_RN_751_0;
wire FE_RN_752_0;
wire FE_RN_753_0;
wire FE_RN_754_0;
wire FE_RN_755_0;
wire FE_RN_756_0;
wire FE_RN_758_0;
wire FE_RN_759_0;
wire FE_RN_764_0;
wire FE_RN_767_0;
wire FE_RN_768_0;
wire FE_RN_769_0;
wire TIMEBOOST_net_16438;
wire FE_RN_772_0;
wire FE_RN_773_0;
wire FE_RN_774_0;
wire FE_RN_775_0;
wire FE_RN_776_0;
wire FE_RN_778_0;
wire FE_RN_779_0;
wire FE_RN_780_0;
wire FE_RN_795_0;
wire FE_RN_796_0;
wire FE_RN_797_0;
wire FE_RN_798_0;
wire FE_RN_7_0;
wire FE_RN_800_0;
wire FE_RN_801_0;
wire FE_RN_802_0;
wire TIMEBOOST_net_10650;
wire TIMEBOOST_net_13713;
wire FE_RN_805_0;
wire FE_RN_806_0;
wire FE_RN_807_0;
wire FE_RN_809_0;
wire FE_RN_810_0;
wire FE_RN_811_0;
wire FE_RN_812_0;
wire FE_RN_814_0;
wire FE_RN_815_0;
wire FE_RN_816_0;
wire FE_RN_817_0;
wire FE_RN_818_0;
wire TIMEBOOST_net_17456;
wire FE_RN_81_0;
wire FE_RN_820_0;
wire FE_RN_821_0;
wire FE_RN_822_0;
wire FE_RN_824_0;
wire TIMEBOOST_net_16866;
wire FE_RN_827_0;
wire FE_RN_828_0;
wire FE_RN_829_0;
wire FE_RN_82_0;
wire TIMEBOOST_net_14657;
wire FE_RN_831_0;
wire FE_RN_832_0;
wire FE_RN_833_0;
wire FE_RN_835_0;
wire FE_RN_836_0;
wire FE_RN_837_0;
wire FE_RN_838_0;
wire FE_RN_839_0;
wire FE_RN_83_0;
wire TIMEBOOST_net_14464;
wire TIMEBOOST_net_16857;
wire FE_RN_843_0;
wire FE_RN_844_0;
wire FE_RN_845_0;
wire TIMEBOOST_net_7255;
wire FE_RN_847_0;
wire FE_RN_862_0;
wire FE_RN_863_0;
wire FE_RN_87_0;
wire FE_RN_880_0;
wire FE_RN_881_0;
wire FE_RN_882_0;
wire TIMEBOOST_net_23550;
wire FE_RN_887_0;
wire FE_RN_888_0;
wire TIMEBOOST_net_13165;
wire FE_RN_88_0;
wire FE_RN_890_0;
wire TIMEBOOST_net_13195;
wire TIMEBOOST_net_23518;
wire FE_RN_893_0;
wire FE_RN_894_0;
wire FE_RN_895_0;
wire FE_RN_896_0;
wire FE_RN_897_0;
wire FE_RN_898_0;
wire FE_RN_899_0;
wire FE_RN_89_0;
wire FE_RN_8_0;
wire FE_RN_900_0;
wire FE_RN_901_0;
wire FE_RN_902_0;
wire FE_RN_904_0;
wire FE_RN_905_0;
wire FE_RN_906_0;
wire FE_RN_907_0;
wire FE_RN_908_0;
wire FE_RN_909_0;
wire FE_RN_90_0;
wire FE_RN_910_0;
wire FE_RN_911_0;
wire FE_RN_912_0;
wire FE_RN_913_0;
wire FE_RN_914_0;
wire FE_RN_915_0;
wire FE_RN_916_0;
wire FE_RN_917_0;
wire FE_RN_91_0;
wire FE_RN_92_0;
wire FE_RN_93_0;
wire FE_RN_94_0;
wire FE_RN_95_0;
wire FE_RN_96_0;
wire FE_RN_97_0;
wire FE_RN_98_0;
wire FE_RN_99_0;
wire FE_RN_9_0;
wire conf_pci_init_complete_out;
wire conf_target_abort_recv_in;
wire conf_w_addr_in;
wire conf_w_addr_in_931;
wire conf_w_addr_in_932;
wire conf_w_addr_in_933;
wire conf_w_addr_in_935;
wire conf_w_addr_in_937;
wire conf_w_addr_in_938;
wire conf_w_addr_in_939;
wire conf_wb_err_addr_in_943;
wire conf_wb_err_addr_in_944;
wire conf_wb_err_addr_in_945;
wire conf_wb_err_addr_in_946;
wire conf_wb_err_addr_in_947;
wire conf_wb_err_addr_in_948;
wire conf_wb_err_addr_in_949;
wire conf_wb_err_addr_in_950;
wire conf_wb_err_addr_in_951;
wire conf_wb_err_addr_in_952;
wire conf_wb_err_addr_in_953;
wire conf_wb_err_addr_in_954;
wire conf_wb_err_addr_in_955;
wire conf_wb_err_addr_in_956;
wire conf_wb_err_addr_in_957;
wire conf_wb_err_addr_in_958;
wire conf_wb_err_addr_in_959;
wire conf_wb_err_addr_in_960;
wire conf_wb_err_addr_in_961;
wire conf_wb_err_addr_in_962;
wire conf_wb_err_addr_in_963;
wire conf_wb_err_addr_in_964;
wire conf_wb_err_addr_in_965;
wire conf_wb_err_addr_in_966;
wire conf_wb_err_addr_in_967;
wire conf_wb_err_addr_in_968;
wire conf_wb_err_addr_in_969;
wire conf_wb_err_addr_in_970;
wire conf_wb_err_addr_in_971;
wire conf_wb_err_bc_in;
wire conf_wb_err_bc_in_846;
wire conf_wb_err_bc_in_847;
wire conf_wb_err_bc_in_848;
wire configuration_cache_line_size_reg;
wire configuration_cache_line_size_reg_2996;
wire configuration_command_bit;
wire configuration_icr_bit2_0;
wire configuration_icr_bit_2961;
wire configuration_icr_bit_2967;
wire configuration_int_meta;
wire configuration_interrupt_line;
wire configuration_interrupt_line_37;
wire configuration_interrupt_line_38;
wire configuration_interrupt_line_39;
wire configuration_interrupt_line_40;
wire configuration_interrupt_line_41;
wire configuration_interrupt_line_42;
wire configuration_interrupt_line_43;
wire configuration_interrupt_out_reg_Q;
wire configuration_isr_bit_1457;
wire configuration_isr_bit_1461;
wire configuration_isr_bit_2975;
wire configuration_isr_bit_618;
wire configuration_isr_bit_631;
wire configuration_meta_cache_lsize_to_wb_bits;
wire configuration_meta_cache_lsize_to_wb_bits_926;
wire configuration_meta_cache_lsize_to_wb_bits_927;
wire configuration_meta_cache_lsize_to_wb_bits_928;
wire configuration_meta_cache_lsize_to_wb_bits_929;
wire configuration_meta_cache_lsize_to_wb_bits_930;
wire configuration_meta_cache_lsize_to_wb_bits_931;
wire configuration_meta_command_bit;
wire configuration_meta_pci_err_cs_bits;
wire configuration_pci_err_addr;
wire configuration_pci_err_addr_471;
wire configuration_pci_err_addr_472;
wire configuration_pci_err_addr_473;
wire configuration_pci_err_addr_474;
wire configuration_pci_err_addr_475;
wire configuration_pci_err_addr_476;
wire configuration_pci_err_addr_477;
wire configuration_pci_err_addr_478;
wire configuration_pci_err_addr_479;
wire configuration_pci_err_addr_480;
wire configuration_pci_err_addr_481;
wire configuration_pci_err_addr_482;
wire configuration_pci_err_addr_483;
wire configuration_pci_err_addr_484;
wire configuration_pci_err_addr_485;
wire configuration_pci_err_addr_486;
wire configuration_pci_err_addr_487;
wire configuration_pci_err_addr_488;
wire configuration_pci_err_addr_489;
wire configuration_pci_err_addr_490;
wire configuration_pci_err_addr_491;
wire configuration_pci_err_addr_492;
wire configuration_pci_err_addr_493;
wire configuration_pci_err_addr_494;
wire configuration_pci_err_addr_495;
wire configuration_pci_err_addr_496;
wire configuration_pci_err_addr_497;
wire configuration_pci_err_addr_498;
wire configuration_pci_err_addr_499;
wire configuration_pci_err_addr_500;
wire configuration_pci_err_addr_501;
wire configuration_pci_err_cs_bit0;
wire configuration_pci_err_cs_bit10;
wire configuration_pci_err_cs_bit31_24;
wire configuration_pci_err_cs_bit8;
wire configuration_pci_err_cs_bit9;
wire configuration_pci_err_cs_bit_464;
wire configuration_pci_err_cs_bit_465;
wire configuration_pci_err_cs_bit_466;
wire configuration_pci_err_cs_bit_467;
wire configuration_pci_err_cs_bit_468;
wire configuration_pci_err_cs_bit_469;
wire configuration_pci_err_cs_bit_470;
wire configuration_pci_err_data;
wire configuration_pci_err_data_502;
wire configuration_pci_err_data_503;
wire configuration_pci_err_data_504;
wire configuration_pci_err_data_505;
wire configuration_pci_err_data_506;
wire configuration_pci_err_data_507;
wire configuration_pci_err_data_508;
wire configuration_pci_err_data_509;
wire configuration_pci_err_data_510;
wire configuration_pci_err_data_511;
wire configuration_pci_err_data_512;
wire configuration_pci_err_data_513;
wire configuration_pci_err_data_514;
wire configuration_pci_err_data_515;
wire configuration_pci_err_data_516;
wire configuration_pci_err_data_517;
wire configuration_pci_err_data_518;
wire configuration_pci_err_data_519;
wire configuration_pci_err_data_520;
wire configuration_pci_err_data_521;
wire configuration_pci_err_data_522;
wire configuration_pci_err_data_523;
wire configuration_pci_err_data_524;
wire configuration_pci_err_data_525;
wire configuration_pci_err_data_526;
wire configuration_pci_err_data_527;
wire configuration_pci_err_data_528;
wire configuration_pci_err_data_529;
wire configuration_pci_err_data_530;
wire configuration_pci_err_data_531;
wire configuration_pci_err_data_532;
wire configuration_rst_inactive;
wire configuration_rst_inactive_sync;
wire configuration_set_isr_bit2;
wire configuration_set_isr_bit2_reg_Q;
wire configuration_set_pci_err_cs_bit8;
wire configuration_set_pci_err_cs_bit8_reg_Q;
wire configuration_status_bit8;
wire configuration_status_bit_322;
wire configuration_status_bit_351;
wire configuration_status_bit_379;
wire configuration_status_bit_407;
wire configuration_status_bit_435;
wire configuration_sync_cache_lsize_to_wb_bits_reg_2__Q;
wire configuration_sync_cache_lsize_to_wb_bits_reg_3__Q;
wire configuration_sync_cache_lsize_to_wb_bits_reg_4__Q;
wire configuration_sync_command_bit0;
wire configuration_sync_command_bit1;
wire configuration_sync_command_bit2;
wire configuration_sync_command_bit6;
wire configuration_sync_command_bit8;
wire configuration_sync_init_complete;
wire configuration_sync_isr_2_del_bit_reg_Q;
wire configuration_sync_isr_2_delayed_bckp_bit;
wire configuration_sync_isr_2_delayed_bckp_bit_reg_Q;
wire configuration_sync_isr_2_delayed_del_bit;
wire configuration_sync_isr_2_delayed_del_bit_reg_Q;
wire configuration_sync_isr_2_meta_bckp_bit;
wire configuration_sync_isr_2_meta_del_bit;
wire configuration_sync_isr_2_sync_bckp_bit;
wire configuration_sync_isr_2_sync_del_bit;
wire configuration_sync_pci_err_cs_8_del_bit_reg_Q;
wire configuration_sync_pci_err_cs_8_delayed_bckp_bit;
wire configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_Q;
wire configuration_sync_pci_err_cs_8_delayed_del_bit;
wire configuration_sync_pci_err_cs_8_delayed_del_bit_reg_Q;
wire configuration_sync_pci_err_cs_8_meta_bckp_bit;
wire configuration_sync_pci_err_cs_8_meta_del_bit;
wire configuration_sync_pci_err_cs_8_sync_bckp_bit;
wire configuration_sync_pci_err_cs_8_sync_del_bit;
wire configuration_wb_err_addr;
wire configuration_wb_err_addr_533;
wire configuration_wb_err_addr_534;
wire configuration_wb_err_addr_535;
wire configuration_wb_err_addr_536;
wire configuration_wb_err_addr_537;
wire configuration_wb_err_addr_538;
wire configuration_wb_err_addr_539;
wire configuration_wb_err_addr_540;
wire configuration_wb_err_addr_541;
wire configuration_wb_err_addr_542;
wire configuration_wb_err_addr_543;
wire configuration_wb_err_addr_544;
wire configuration_wb_err_addr_545;
wire configuration_wb_err_addr_546;
wire configuration_wb_err_addr_547;
wire configuration_wb_err_addr_548;
wire configuration_wb_err_addr_549;
wire configuration_wb_err_addr_550;
wire configuration_wb_err_addr_551;
wire configuration_wb_err_addr_552;
wire configuration_wb_err_addr_553;
wire configuration_wb_err_addr_554;
wire configuration_wb_err_addr_555;
wire configuration_wb_err_addr_556;
wire configuration_wb_err_addr_557;
wire configuration_wb_err_addr_558;
wire configuration_wb_err_addr_559;
wire configuration_wb_err_addr_560;
wire configuration_wb_err_addr_561;
wire configuration_wb_err_addr_562;
wire configuration_wb_err_addr_563;
wire configuration_wb_err_cs_bit0;
wire configuration_wb_err_cs_bit31_24;
wire configuration_wb_err_cs_bit8;
wire configuration_wb_err_cs_bit9;
wire configuration_wb_err_cs_bit_564;
wire configuration_wb_err_cs_bit_565;
wire configuration_wb_err_cs_bit_566;
wire configuration_wb_err_cs_bit_567;
wire configuration_wb_err_cs_bit_568;
wire configuration_wb_err_cs_bit_569;
wire configuration_wb_err_cs_bit_570;
wire configuration_wb_err_data;
wire configuration_wb_err_data_571;
wire configuration_wb_err_data_572;
wire configuration_wb_err_data_573;
wire configuration_wb_err_data_574;
wire configuration_wb_err_data_575;
wire configuration_wb_err_data_576;
wire configuration_wb_err_data_577;
wire configuration_wb_err_data_578;
wire configuration_wb_err_data_579;
wire configuration_wb_err_data_580;
wire configuration_wb_err_data_581;
wire configuration_wb_err_data_582;
wire configuration_wb_err_data_583;
wire configuration_wb_err_data_584;
wire configuration_wb_err_data_585;
wire configuration_wb_err_data_586;
wire configuration_wb_err_data_587;
wire configuration_wb_err_data_588;
wire configuration_wb_err_data_589;
wire configuration_wb_err_data_590;
wire configuration_wb_err_data_591;
wire configuration_wb_err_data_592;
wire configuration_wb_err_data_593;
wire configuration_wb_err_data_594;
wire configuration_wb_err_data_595;
wire configuration_wb_err_data_596;
wire configuration_wb_err_data_597;
wire configuration_wb_err_data_598;
wire configuration_wb_err_data_599;
wire configuration_wb_err_data_600;
wire configuration_wb_err_data_601;
wire g15_p;
wire g17_p;
wire g22_p;
wire g52252_p;
wire g52253_p;
wire g52393_db;
wire g52393_sb;
wire TIMEBOOST_net_23418;
wire g52394_sb;
wire TIMEBOOST_net_10090;
wire TIMEBOOST_net_9704;
wire g52395_sb;
wire TIMEBOOST_net_10091;
wire TIMEBOOST_net_9755;
wire g52396_sb;
wire TIMEBOOST_net_21429;
wire g52397_sb;
wire n_9019;
wire g52398_sb;
wire g52399_db;
wire g52399_sb;
wire TIMEBOOST_net_22378;
wire g52400_sb;
wire g52401_db;
wire g52401_sb;
wire TIMEBOOST_net_21387;
wire g52402_db;
wire g52402_sb;
wire g52403_db;
wire g52403_sb;
wire TIMEBOOST_net_10204;
wire TIMEBOOST_net_20519;
wire g52404_sb;
wire TIMEBOOST_net_23523;
wire g52405_db;
wire g52405_sb;
wire g52439_db;
wire TIMEBOOST_net_10088;
wire TIMEBOOST_net_20458;
wire g52440_sb;
wire TIMEBOOST_net_10089;
wire TIMEBOOST_net_12680;
wire g52441_sb;
wire TIMEBOOST_net_10412;
wire TIMEBOOST_net_12683;
wire g52442_sb;
wire TIMEBOOST_net_21851;
wire g52443_sb;
wire TIMEBOOST_net_10411;
wire TIMEBOOST_net_23463;
wire g52444_sb;
wire TIMEBOOST_net_16522;
wire g52445_db;
wire TIMEBOOST_net_10049;
wire g52446_db;
wire g52446_sb;
wire g52447_db;
wire g52447_sb;
wire TIMEBOOST_net_10904;
wire g52448_sb;
wire TIMEBOOST_net_10079;
wire g52449_sb;
wire TIMEBOOST_net_14387;
wire g52450_sb;
wire TIMEBOOST_net_10098;
wire TIMEBOOST_net_23449;
wire g52451_sb;
wire TIMEBOOST_net_10078;
wire g52452_sb;
wire TIMEBOOST_net_22372;
wire g52454_sb;
wire g52455_da;
wire TIMEBOOST_net_23164;
wire g52455_sb;
wire g52456_da;
wire g52456_sb;
wire TIMEBOOST_net_20769;
wire TIMEBOOST_net_20398;
wire g52457_sb;
wire TIMEBOOST_net_20770;
wire TIMEBOOST_net_16725;
wire g52458_sb;
wire g52459_da;
wire g52459_sb;
wire TIMEBOOST_net_20771;
wire TIMEBOOST_net_20389;
wire g52460_sb;
wire TIMEBOOST_net_20772;
wire g52461_sb;
wire g52462_da;
wire TIMEBOOST_net_16749;
wire g52462_sb;
wire TIMEBOOST_net_20773;
wire TIMEBOOST_net_16518;
wire g52463_sb;
wire g52464_da;
wire TIMEBOOST_net_20377;
wire g52464_sb;
wire TIMEBOOST_net_20774;
wire TIMEBOOST_net_11360;
wire g52466_da;
wire TIMEBOOST_net_16677;
wire g52466_sb;
wire TIMEBOOST_net_20775;
wire g52468_da;
wire TIMEBOOST_net_16674;
wire TIMEBOOST_net_20776;
wire TIMEBOOST_net_20777;
wire g52470_sb;
wire TIMEBOOST_net_20778;
wire g52472_da;
wire TIMEBOOST_net_16517;
wire TIMEBOOST_net_20779;
wire TIMEBOOST_net_12737;
wire TIMEBOOST_net_20780;
wire TIMEBOOST_net_16727;
wire TIMEBOOST_net_20781;
wire TIMEBOOST_net_16054;
wire g52476_da;
wire TIMEBOOST_net_14538;
wire g52476_sb;
wire g52477_da;
wire TIMEBOOST_net_10554;
wire g52477_sb;
wire g52478_da;
wire g64241_db;
wire g52478_sb;
wire g52479_da;
wire TIMEBOOST_net_13718;
wire g52479_sb;
wire TIMEBOOST_net_14454;
wire TIMEBOOST_net_14298;
wire TIMEBOOST_net_14658;
wire g52482_da;
wire g52482_sb;
wire TIMEBOOST_net_20782;
wire TIMEBOOST_net_14266;
wire TIMEBOOST_net_14656;
wire TIMEBOOST_net_20783;
wire TIMEBOOST_net_17362;
wire g52495_p;
wire g52496_p;
wire g52497_p;
wire g52498_p;
wire TIMEBOOST_net_17062;
wire TIMEBOOST_net_16064;
wire g52503_sb;
wire TIMEBOOST_net_12493;
wire TIMEBOOST_net_21185;
wire g52504_sb;
wire TIMEBOOST_net_17063;
wire g52505_sb;
wire TIMEBOOST_net_16594;
wire g52506_sb;
wire TIMEBOOST_net_20344;
wire TIMEBOOST_net_22575;
wire g52507_sb;
wire g52508_sb;
wire TIMEBOOST_net_12494;
wire TIMEBOOST_net_16595;
wire g52509_sb;
wire TIMEBOOST_net_17108;
wire g52510_sb;
wire TIMEBOOST_net_17205;
wire TIMEBOOST_net_14267;
wire g52511_sb;
wire TIMEBOOST_net_14268;
wire g52512_sb;
wire TIMEBOOST_net_6978;
wire TIMEBOOST_net_14269;
wire g52513_sb;
wire TIMEBOOST_net_22588;
wire g52514_sb;
wire TIMEBOOST_net_13722;
wire g52515_sb;
wire TIMEBOOST_net_20271;
wire g52516_sb;
wire TIMEBOOST_net_14602;
wire g52517_sb;
wire TIMEBOOST_net_17375;
wire TIMEBOOST_net_22357;
wire g52518_sb;
wire g52519_sb;
wire TIMEBOOST_net_12590;
wire TIMEBOOST_net_16686;
wire g52520_sb;
wire TIMEBOOST_net_14532;
wire g52521_sb;
wire TIMEBOOST_net_12375;
wire g52522_sb;
wire TIMEBOOST_net_20549;
wire g52523_sb;
wire TIMEBOOST_net_20196;
wire TIMEBOOST_net_13729;
wire g52524_sb;
wire g52525_sb;
wire TIMEBOOST_net_12377;
wire TIMEBOOST_net_16515;
wire g52526_sb;
wire g52527_sb;
wire g52528_sb;
wire TIMEBOOST_net_21949;
wire TIMEBOOST_net_16052;
wire g52529_sb;
wire TIMEBOOST_net_16597;
wire g52530_sb;
wire TIMEBOOST_net_22324;
wire g52531_sb;
wire TIMEBOOST_net_12508;
wire TIMEBOOST_net_20917;
wire g52532_sb;
wire TIMEBOOST_net_22325;
wire g52533_sb;
wire TIMEBOOST_net_23464;
wire g52534_sb;
wire TIMEBOOST_net_13375;
wire TIMEBOOST_net_16922;
wire g52590_sb;
wire TIMEBOOST_net_5465;
wire g52591_sb;
wire TIMEBOOST_net_5466;
wire g52592_sb;
wire TIMEBOOST_net_5467;
wire g52593_sb;
wire TIMEBOOST_net_12411;
wire g52594_sb;
wire TIMEBOOST_net_16440;
wire g52595_sb;
wire g54176_da;
wire g52596_sb;
wire g52597_db;
wire g52597_sb;
wire g52598_sb;
wire TIMEBOOST_net_21435;
wire g52599_sb;
wire TIMEBOOST_net_21903;
wire g52600_db;
wire g52600_sb;
wire TIMEBOOST_net_17001;
wire g52601_sb;
wire TIMEBOOST_net_17002;
wire g52602_sb;
wire TIMEBOOST_net_17246;
wire g52603_sb;
wire TIMEBOOST_net_21747;
wire g52604_sb;
wire TIMEBOOST_net_12251;
wire g52605_sb;
wire g52606_db;
wire g52606_sb;
wire TIMEBOOST_net_9803;
wire g52607_sb;
wire TIMEBOOST_net_22877;
wire TIMEBOOST_net_12790;
wire g52608_sb;
wire TIMEBOOST_net_17407;
wire g52609_sb;
wire g52610_sb;
wire TIMEBOOST_net_13461;
wire TIMEBOOST_net_17415;
wire g52611_sb;
wire TIMEBOOST_net_21585;
wire g52612_sb;
wire TIMEBOOST_net_21529;
wire g52614_sb;
wire TIMEBOOST_net_13850;
wire g52616_sb;
wire TIMEBOOST_net_12405;
wire g52617_sb;
wire g54202_da;
wire TIMEBOOST_net_22745;
wire g52618_sb;
wire g54200_da;
wire g52619_sb;
wire TIMEBOOST_net_12253;
wire TIMEBOOST_net_13849;
wire g52620_sb;
wire TIMEBOOST_net_22746;
wire g52621_sb;
wire TIMEBOOST_net_12254;
wire TIMEBOOST_net_16707;
wire g52622_sb;
wire g52623_p;
wire TIMEBOOST_net_15474;
wire g52624_sb;
wire g52625_sb;
wire TIMEBOOST_net_22494;
wire TIMEBOOST_net_22141;
wire g52626_sb;
wire TIMEBOOST_net_13928;
wire g52627_sb;
wire TIMEBOOST_net_21535;
wire TIMEBOOST_net_17526;
wire g52628_sb;
wire TIMEBOOST_net_21712;
wire g52629_sb;
wire TIMEBOOST_net_13519;
wire TIMEBOOST_net_20450;
wire g52630_sb;
wire TIMEBOOST_net_15986;
wire g60682_da;
wire g52631_sb;
wire TIMEBOOST_net_9504;
wire g52632_sb;
wire TIMEBOOST_net_21558;
wire TIMEBOOST_net_14977;
wire g52633_sb;
wire TIMEBOOST_net_13929;
wire TIMEBOOST_net_14803;
wire g52634_sb;
wire g52635_sb;
wire TIMEBOOST_net_21554;
wire g52636_sb;
wire TIMEBOOST_net_13520;
wire g52637_sb;
wire TIMEBOOST_net_21548;
wire g52638_db;
wire g52638_sb;
wire TIMEBOOST_net_8112;
wire TIMEBOOST_net_17318;
wire g52639_sb;
wire TIMEBOOST_net_20784;
wire TIMEBOOST_net_8111;
wire g52641_sb;
wire TIMEBOOST_net_12569;
wire g52642_sb;
wire TIMEBOOST_net_20256;
wire g64944_db;
wire g52643_sb;
wire TIMEBOOST_net_8118;
wire TIMEBOOST_net_8615;
wire g52644_sb;
wire TIMEBOOST_net_16757;
wire g52645_sb;
wire g52646_sb;
wire TIMEBOOST_net_13245;
wire g52647_sb;
wire TIMEBOOST_net_14978;
wire g52648_sb;
wire TIMEBOOST_net_21997;
wire TIMEBOOST_net_13246;
wire g52650_db;
wire g52650_sb;
wire TIMEBOOST_net_21739;
wire g52651_sb;
wire TIMEBOOST_net_8110;
wire TIMEBOOST_net_12931;
wire g52652_sb;
wire TIMEBOOST_net_21651;
wire TIMEBOOST_net_14979;
wire g52653_sb;
wire g52675_p;
wire g52714_p;
wire g52865_p;
wire TIMEBOOST_net_17509;
wire TIMEBOOST_net_23504;
wire g52876_sb;
wire TIMEBOOST_net_17484;
wire TIMEBOOST_net_14717;
wire g52877_sb;
wire TIMEBOOST_net_14967;
wire TIMEBOOST_net_17448;
wire g52878_sb;
wire g58774_da;
wire TIMEBOOST_net_20181;
wire g52879_sb;
wire g52880_sb;
wire TIMEBOOST_net_10976;
wire g52881_sb;
wire g52_p;
wire g53011_p;
wire g53012_p;
wire g53014_p;
wire g53015_p;
wire g53016_p;
wire g53017_p;
wire g53018_p;
wire g53022_p;
wire g53026_p;
wire g53031_p;
wire g53035_p;
wire g53039_p;
wire g53069_p;
wire g53071_p;
wire g53072_p;
wire g53073_p;
wire g53074_p;
wire g53075_p;
wire g53076_p;
wire g53077_p;
wire g53078_p;
wire g53079_p;
wire g53080_p;
wire g53082_p;
wire g53083_p;
wire g53084_p;
wire g53087_p;
wire g53098_p;
wire TIMEBOOST_net_23115;
wire g53141_p;
wire g53142_p;
wire g53154_p;
wire g53155_p;
wire g53158_p;
wire g53159_p;
wire g53163_p;
wire g53167_p;
wire g53170_p;
wire g53171_p;
wire g53174_p;
wire g53175_p;
wire g53182_p;
wire g53183_p;
wire g53187_p;
wire g53199_p;
wire g53203_p;
wire g53206_p;
wire g53207_p;
wire g53210_p;
wire g53211_p;
wire g53214_p;
wire g53222_p;
wire g53223_p;
wire g53226_p;
wire g53230_p;
wire g53231_p;
wire g53234_p;
wire g53235_p;
wire g53238_p;
wire g53239_p;
wire g53242_p;
wire g53243_p;
wire g53250_p;
wire g53251_p;
wire g53254_p;
wire g53255_p;
wire g53258_p;
wire g53259_p;
wire g53262_p;
wire g53263_p;
wire g53267_p;
wire g53268_p;
wire g53275_p;
wire g53276_p;
wire g53288_p;
wire g53289_p;
wire g53298_p;
wire g53301_p;
wire g53302_p;
wire g53310_p;
wire g53314_p;
wire g53709_p;
wire g53726_p;
wire g53729_p;
wire g53752_p;
wire g53891_da;
wire g53891_db;
wire g53892_sb;
wire g53893_da;
wire g53893_db;
wire TIMEBOOST_net_13515;
wire TIMEBOOST_net_10610;
wire g53897_sb;
wire TIMEBOOST_net_10130;
wire g53898_sb;
wire TIMEBOOST_net_10129;
wire TIMEBOOST_net_20788;
wire g53899_sb;
wire g53900_sb;
wire TIMEBOOST_net_20910;
wire TIMEBOOST_net_16549;
wire g53901_sb;
wire TIMEBOOST_net_22579;
wire TIMEBOOST_net_16550;
wire g53902_sb;
wire TIMEBOOST_net_16942;
wire TIMEBOOST_net_16551;
wire g53903_sb;
wire TIMEBOOST_net_16552;
wire g53904_sb;
wire TIMEBOOST_net_23338;
wire TIMEBOOST_net_16553;
wire g53905_sb;
wire TIMEBOOST_net_16935;
wire TIMEBOOST_net_16554;
wire g53906_sb;
wire TIMEBOOST_net_10120;
wire TIMEBOOST_net_16555;
wire g53907_sb;
wire TIMEBOOST_net_10118;
wire TIMEBOOST_net_16556;
wire g53908_sb;
wire TIMEBOOST_net_10117;
wire TIMEBOOST_net_16557;
wire g53909_sb;
wire TIMEBOOST_net_10116;
wire TIMEBOOST_net_22404;
wire g53910_sb;
wire TIMEBOOST_net_10115;
wire g53911_sb;
wire TIMEBOOST_net_10114;
wire TIMEBOOST_net_22390;
wire g53912_sb;
wire TIMEBOOST_net_10113;
wire TIMEBOOST_net_22391;
wire g53913_sb;
wire TIMEBOOST_net_10112;
wire TIMEBOOST_net_22596;
wire g53914_sb;
wire TIMEBOOST_net_13897;
wire TIMEBOOST_net_16563;
wire g53915_sb;
wire TIMEBOOST_net_10109;
wire g53916_sb;
wire TIMEBOOST_net_10108;
wire TIMEBOOST_net_16565;
wire g53917_sb;
wire TIMEBOOST_net_10107;
wire TIMEBOOST_net_16566;
wire g53918_sb;
wire TIMEBOOST_net_10106;
wire g53919_sb;
wire TIMEBOOST_net_10105;
wire TIMEBOOST_net_10596;
wire g53920_sb;
wire TIMEBOOST_net_10104;
wire g53921_sb;
wire TIMEBOOST_net_10103;
wire g53922_sb;
wire TIMEBOOST_net_10102;
wire TIMEBOOST_net_16880;
wire g53923_sb;
wire TIMEBOOST_net_10100;
wire g53924_sb;
wire TIMEBOOST_net_10099;
wire TIMEBOOST_net_16571;
wire g53925_sb;
wire TIMEBOOST_net_10097;
wire TIMEBOOST_net_16572;
wire g53926_sb;
wire TIMEBOOST_net_10096;
wire TIMEBOOST_net_16573;
wire g53927_sb;
wire TIMEBOOST_net_10095;
wire TIMEBOOST_net_10597;
wire g53928_sb;
wire TIMEBOOST_net_10094;
wire TIMEBOOST_net_14586;
wire g53929_sb;
wire TIMEBOOST_net_10093;
wire TIMEBOOST_net_16574;
wire g53930_sb;
wire TIMEBOOST_net_10092;
wire g53931_sb;
wire TIMEBOOST_net_10381;
wire g53932_sb;
wire g53935_da;
wire g53935_db;
wire TIMEBOOST_net_14105;
wire TIMEBOOST_net_17404;
wire g53937_sb;
wire TIMEBOOST_net_16739;
wire g53939_db;
wire g53939_sb;
wire TIMEBOOST_net_13517;
wire TIMEBOOST_net_10757;
wire g53940_sb;
wire TIMEBOOST_net_13516;
wire TIMEBOOST_net_17471;
wire g53942_db;
wire TIMEBOOST_net_22949;
wire TIMEBOOST_net_22393;
wire TIMEBOOST_net_22950;
wire TIMEBOOST_net_22295;
wire g53945_da;
wire g53946_da;
wire TIMEBOOST_net_5512;
wire g53946_sb;
wire TIMEBOOST_net_22893;
wire TIMEBOOST_net_5513;
wire g53990_p;
wire TIMEBOOST_net_17238;
wire TIMEBOOST_net_13390;
wire g54030_sb;
wire TIMEBOOST_net_34;
wire g54038_db;
wire g54038_sb;
wire TIMEBOOST_net_10413;
wire g54039_sb;
wire TIMEBOOST_net_10409;
wire g54040_sb;
wire g54131_da;
wire TIMEBOOST_net_16499;
wire g54131_sb;
wire TIMEBOOST_net_21415;
wire g54132_sb;
wire g58401_db;
wire g54133_sb;
wire TIMEBOOST_net_9414;
wire TIMEBOOST_net_22182;
wire g54134_sb;
wire TIMEBOOST_net_9415;
wire TIMEBOOST_net_21228;
wire g54135_sb;
wire TIMEBOOST_net_13611;
wire TIMEBOOST_net_14714;
wire g54137_sb;
wire TIMEBOOST_net_9416;
wire TIMEBOOST_net_7999;
wire g54138_sb;
wire g54139_da;
wire TIMEBOOST_net_16782;
wire g54140_sb;
wire TIMEBOOST_net_13532;
wire g54141_sb;
wire TIMEBOOST_net_5438;
wire TIMEBOOST_net_13671;
wire g54143_sb;
wire TIMEBOOST_net_13621;
wire g54144_sb;
wire TIMEBOOST_net_9417;
wire TIMEBOOST_net_14960;
wire g54145_sb;
wire TIMEBOOST_net_15076;
wire g54146_sb;
wire TIMEBOOST_net_23385;
wire g54147_sb;
wire TIMEBOOST_net_12240;
wire g54148_sb;
wire TIMEBOOST_net_9418;
wire TIMEBOOST_net_23415;
wire g54149_sb;
wire TIMEBOOST_net_15951;
wire TIMEBOOST_net_21317;
wire g54150_sb;
wire TIMEBOOST_net_5440;
wire TIMEBOOST_net_13701;
wire g54151_sb;
wire TIMEBOOST_net_5441;
wire TIMEBOOST_net_20895;
wire g54152_sb;
wire TIMEBOOST_net_9419;
wire TIMEBOOST_net_20893;
wire g54153_sb;
wire TIMEBOOST_net_9420;
wire TIMEBOOST_net_7996;
wire g54154_sb;
wire TIMEBOOST_net_9421;
wire g54155_sb;
wire TIMEBOOST_net_9422;
wire TIMEBOOST_net_7995;
wire g54157_sb;
wire TIMEBOOST_net_21261;
wire g54158_sb;
wire TIMEBOOST_net_15352;
wire TIMEBOOST_net_12756;
wire g54160_sb;
wire TIMEBOOST_net_14113;
wire TIMEBOOST_net_14988;
wire g54161_sb;
wire g54163_da;
wire TIMEBOOST_net_22783;
wire TIMEBOOST_net_14987;
wire g54164_sb;
wire TIMEBOOST_net_12783;
wire TIMEBOOST_net_23157;
wire g54167_db;
wire g54167_sb;
wire TIMEBOOST_net_5442;
wire TIMEBOOST_net_20956;
wire g54168_sb;
wire g54169_sb;
wire TIMEBOOST_net_13936;
wire n_1617;
wire g54170_sb;
wire TIMEBOOST_net_13490;
wire TIMEBOOST_net_22788;
wire g54171_sb;
wire g54172_sb;
wire g54173_sb;
wire TIMEBOOST_net_15477;
wire g54174_db;
wire g54174_sb;
wire g54175_da;
wire g54175_sb;
wire TIMEBOOST_net_7530;
wire g54176_sb;
wire TIMEBOOST_net_17302;
wire g54177_sb;
wire g54178_da;
wire TIMEBOOST_net_7529;
wire g54178_sb;
wire g54179_sb;
wire TIMEBOOST_net_17544;
wire g54180_db;
wire g54180_sb;
wire g54181_da;
wire TIMEBOOST_net_7528;
wire g54181_sb;
wire TIMEBOOST_net_14331;
wire g54182_db;
wire g54182_sb;
wire TIMEBOOST_net_13935;
wire TIMEBOOST_net_22263;
wire g54183_sb;
wire TIMEBOOST_net_14625;
wire g54184_db;
wire g54184_sb;
wire TIMEBOOST_net_20241;
wire g54185_db;
wire g54185_sb;
wire TIMEBOOST_net_5449;
wire g66456_da;
wire g54186_sb;
wire TIMEBOOST_net_13938;
wire TIMEBOOST_net_16003;
wire g54187_sb;
wire TIMEBOOST_net_14626;
wire g54188_db;
wire g54188_sb;
wire TIMEBOOST_net_21733;
wire g54189_db;
wire g54189_sb;
wire TIMEBOOST_net_15904;
wire TIMEBOOST_net_13564;
wire g54190_sb;
wire TIMEBOOST_net_21151;
wire TIMEBOOST_net_84;
wire g54191_sb;
wire TIMEBOOST_net_14429;
wire TIMEBOOST_net_13554;
wire g54192_sb;
wire TIMEBOOST_net_7519;
wire g54193_sb;
wire g54194_sb;
wire TIMEBOOST_net_7504;
wire g54195_sb;
wire TIMEBOOST_net_20217;
wire TIMEBOOST_net_23308;
wire g54196_sb;
wire TIMEBOOST_net_21355;
wire g54197_sb;
wire TIMEBOOST_net_17083;
wire TIMEBOOST_net_23307;
wire g54198_sb;
wire g54199_sb;
wire TIMEBOOST_net_21914;
wire TIMEBOOST_net_13551;
wire g54200_sb;
wire TIMEBOOST_net_20920;
wire TIMEBOOST_net_14114;
wire g54201_sb;
wire TIMEBOOST_net_21209;
wire TIMEBOOST_net_13550;
wire g54202_sb;
wire TIMEBOOST_net_21384;
wire g54203_sb;
wire TIMEBOOST_net_27;
wire TIMEBOOST_net_16520;
wire TIMEBOOST_net_51;
wire g54205_sb;
wire TIMEBOOST_net_16718;
wire g54207_sb;
wire TIMEBOOST_net_15975;
wire TIMEBOOST_net_11920;
wire TIMEBOOST_net_20210;
wire g54209_sb;
wire TIMEBOOST_net_10445;
wire TIMEBOOST_net_14667;
wire TIMEBOOST_net_16291;
wire TIMEBOOST_net_16521;
wire TIMEBOOST_net_21172;
wire TIMEBOOST_net_17426;
wire TIMEBOOST_net_28;
wire TIMEBOOST_net_21705;
wire TIMEBOOST_net_12773;
wire g54216_da;
wire g54216_sb;
wire TIMEBOOST_net_21703;
wire TIMEBOOST_net_12820;
wire g54219_sb;
wire TIMEBOOST_net_29;
wire TIMEBOOST_net_20438;
wire TIMEBOOST_net_12507;
wire TIMEBOOST_net_22057;
wire TIMEBOOST_net_22082;
wire TIMEBOOST_net_30;
wire TIMEBOOST_net_14661;
wire TIMEBOOST_net_13746;
wire TIMEBOOST_net_13548;
wire TIMEBOOST_net_22026;
wire TIMEBOOST_net_14530;
wire TIMEBOOST_net_12917;
wire TIMEBOOST_net_13590;
wire TIMEBOOST_net_14986;
wire g54234_sb;
wire TIMEBOOST_net_15066;
wire g54235_sb;
wire TIMEBOOST_net_7684;
wire TIMEBOOST_net_14961;
wire g54236_sb;
wire g54237_sb;
wire TIMEBOOST_net_13605;
wire TIMEBOOST_net_14984;
wire g54238_sb;
wire TIMEBOOST_net_14943;
wire g54239_sb;
wire TIMEBOOST_net_11311;
wire g54244_sb;
wire TIMEBOOST_net_22219;
wire TIMEBOOST_net_15103;
wire g54304_sb;
wire TIMEBOOST_net_14718;
wire g54305_sb;
wire g54306_sb;
wire TIMEBOOST_net_21029;
wire g54309_sb;
wire TIMEBOOST_net_14796;
wire TIMEBOOST_net_22171;
wire g54310_sb;
wire g54311_db;
wire g54311_sb;
wire g54312_sb;
wire TIMEBOOST_net_14942;
wire TIMEBOOST_net_21067;
wire g54314_sb;
wire TIMEBOOST_net_14886;
wire g54315_db;
wire g54315_sb;
wire TIMEBOOST_net_11486;
wire TIMEBOOST_net_20612;
wire g54316_sb;
wire TIMEBOOST_net_14874;
wire g54317_sb;
wire TIMEBOOST_net_20556;
wire TIMEBOOST_net_13526;
wire g54318_sb;
wire TIMEBOOST_net_13689;
wire g65797_db;
wire g54319_sb;
wire g61974_db;
wire TIMEBOOST_net_9507;
wire g54320_sb;
wire TIMEBOOST_net_23461;
wire TIMEBOOST_net_13527;
wire g54321_sb;
wire g61973_db;
wire TIMEBOOST_net_22251;
wire g54322_sb;
wire TIMEBOOST_net_14030;
wire g54323_sb;
wire g61972_db;
wire g54324_sb;
wire TIMEBOOST_net_22170;
wire g54325_sb;
wire g54326_sb;
wire TIMEBOOST_net_21250;
wire TIMEBOOST_net_16500;
wire g54328_sb;
wire g54329_p;
wire TIMEBOOST_net_13581;
wire g54330_sb;
wire g54331_sb;
wire TIMEBOOST_net_20971;
wire TIMEBOOST_net_14912;
wire g54332_sb;
wire TIMEBOOST_net_23391;
wire TIMEBOOST_net_21310;
wire g54333_sb;
wire TIMEBOOST_net_23386;
wire TIMEBOOST_net_21293;
wire g54334_sb;
wire TIMEBOOST_net_21313;
wire g54335_sb;
wire TIMEBOOST_net_22158;
wire g54336_sb;
wire TIMEBOOST_net_12603;
wire TIMEBOOST_net_20331;
wire g54337_sb;
wire TIMEBOOST_net_21339;
wire g54338_sb;
wire TIMEBOOST_net_17395;
wire g54339_sb;
wire g54340_sb;
wire g54341_sb;
wire TIMEBOOST_net_17423;
wire g54342_sb;
wire TIMEBOOST_net_12676;
wire TIMEBOOST_net_15099;
wire g54343_sb;
wire TIMEBOOST_net_13362;
wire g54344_sb;
wire g54345_sb;
wire TIMEBOOST_net_10077;
wire TIMEBOOST_net_16380;
wire g54346_sb;
wire TIMEBOOST_net_10076;
wire g54347_sb;
wire TIMEBOOST_net_10075;
wire TIMEBOOST_net_17296;
wire g54348_sb;
wire TIMEBOOST_net_13518;
wire g52469_da;
wire g54349_sb;
wire TIMEBOOST_net_10074;
wire TIMEBOOST_net_14426;
wire g54350_sb;
wire TIMEBOOST_net_10073;
wire TIMEBOOST_net_10420;
wire g54351_sb;
wire TIMEBOOST_net_10072;
wire g54352_sb;
wire TIMEBOOST_net_13370;
wire g54353_sb;
wire TIMEBOOST_net_10087;
wire g54354_sb;
wire TIMEBOOST_net_10071;
wire g54355_sb;
wire TIMEBOOST_net_10070;
wire g54356_sb;
wire TIMEBOOST_net_10086;
wire g54357_sb;
wire TIMEBOOST_net_10085;
wire TIMEBOOST_net_11317;
wire g54358_sb;
wire TIMEBOOST_net_10084;
wire TIMEBOOST_net_11318;
wire g54359_sb;
wire TIMEBOOST_net_10083;
wire TIMEBOOST_net_15188;
wire g54360_sb;
wire TIMEBOOST_net_10082;
wire g54361_sb;
wire TIMEBOOST_net_10081;
wire TIMEBOOST_net_11321;
wire g54362_sb;
wire TIMEBOOST_net_10080;
wire TIMEBOOST_net_11322;
wire g54363_sb;
wire TIMEBOOST_net_23492;
wire TIMEBOOST_net_17396;
wire g54364_sb;
wire TIMEBOOST_net_21831;
wire g54365_sb;
wire TIMEBOOST_net_21349;
wire g54366_sb;
wire TIMEBOOST_net_15035;
wire g54367_sb;
wire TIMEBOOST_net_10069;
wire TIMEBOOST_net_17459;
wire g54368_sb;
wire TIMEBOOST_net_10068;
wire TIMEBOOST_net_16377;
wire g54369_sb;
wire g54453_p;
wire g54456_p;
wire g54458_p;
wire g54465_p;
wire TIMEBOOST_net_22462;
wire TIMEBOOST_net_21743;
wire g54471_sb;
wire TIMEBOOST_net_12378;
wire g54472_sb;
wire TIMEBOOST_net_9815;
wire g54484_sb;
wire g59231_db;
wire g54485_sb;
wire TIMEBOOST_net_12739;
wire g54486_sb;
wire TIMEBOOST_net_20635;
wire g58800_db;
wire g54487_sb;
wire TIMEBOOST_net_12607;
wire TIMEBOOST_net_22772;
wire g54488_sb;
wire TIMEBOOST_net_13071;
wire g54489_sb;
wire TIMEBOOST_net_12381;
wire g54490_sb;
wire TIMEBOOST_net_17376;
wire g54491_sb;
wire TIMEBOOST_net_13070;
wire g54492_sb;
wire TIMEBOOST_net_17440;
wire g54493_sb;
wire TIMEBOOST_net_12600;
wire TIMEBOOST_net_21794;
wire g54494_sb;
wire g54495_sb;
wire g54568_p;
wire g54569_p;
wire g54572_p;
wire g54573_p;
wire g54574_p;
wire g54579_p;
wire g54580_p;
wire g54581_p;
wire g54586_p;
wire g54587_p;
wire g54591_p;
wire g54593_p;
wire g54594_p;
wire g54595_p;
wire g54596_p;
wire g54597_p;
wire g54601_p;
wire g54603_p;
wire g54606_p;
wire TIMEBOOST_net_20156;
wire g55851_sb;
wire TIMEBOOST_net_20244;
wire TIMEBOOST_net_16180;
wire g55852_sb;
wire g55853_sb;
wire g56933_sb;
wire TIMEBOOST_net_22282;
wire g52475_da;
wire g56934_sb;
wire g57030_p;
wire g57033_p;
wire TIMEBOOST_net_17333;
wire g57034_sb;
wire TIMEBOOST_net_6755;
wire g57035_sb;
wire TIMEBOOST_net_10527;
wire TIMEBOOST_net_16367;
wire g57036_sb;
wire TIMEBOOST_net_17227;
wire g57037_sb;
wire TIMEBOOST_net_10442;
wire g57038_sb;
wire TIMEBOOST_net_6756;
wire TIMEBOOST_net_16152;
wire g57039_sb;
wire TIMEBOOST_net_6757;
wire TIMEBOOST_net_22481;
wire g57040_sb;
wire TIMEBOOST_net_11298;
wire TIMEBOOST_net_20545;
wire g57041_sb;
wire TIMEBOOST_net_20437;
wire g57042_sb;
wire TIMEBOOST_net_10506;
wire g57043_sb;
wire TIMEBOOST_net_21192;
wire TIMEBOOST_net_10066;
wire g57044_sb;
wire TIMEBOOST_net_21143;
wire g57045_sb;
wire TIMEBOOST_net_6758;
wire TIMEBOOST_net_10235;
wire g57046_sb;
wire TIMEBOOST_net_10065;
wire g57047_sb;
wire g57048_sb;
wire TIMEBOOST_net_6759;
wire TIMEBOOST_net_16155;
wire g57049_sb;
wire TIMEBOOST_net_6760;
wire TIMEBOOST_net_16156;
wire g57050_sb;
wire TIMEBOOST_net_17154;
wire TIMEBOOST_net_16371;
wire g57051_sb;
wire TIMEBOOST_net_10531;
wire g57052_sb;
wire TIMEBOOST_net_22740;
wire g57053_sb;
wire TIMEBOOST_net_14104;
wire TIMEBOOST_net_6761;
wire TIMEBOOST_net_15718;
wire g57055_sb;
wire TIMEBOOST_net_17136;
wire TIMEBOOST_net_23420;
wire g57056_sb;
wire TIMEBOOST_net_17153;
wire g57057_sb;
wire TIMEBOOST_net_11894;
wire g57058_sb;
wire TIMEBOOST_net_22457;
wire g57059_sb;
wire TIMEBOOST_net_22456;
wire g57060_sb;
wire TIMEBOOST_net_14397;
wire g57061_sb;
wire TIMEBOOST_net_17150;
wire g57062_sb;
wire TIMEBOOST_net_16183;
wire g57063_sb;
wire TIMEBOOST_net_14213;
wire g57064_sb;
wire TIMEBOOST_net_20535;
wire g57065_sb;
wire TIMEBOOST_net_22959;
wire g57066_sb;
wire TIMEBOOST_net_22360;
wire g57067_sb;
wire g57068_sb;
wire g57069_sb;
wire TIMEBOOST_net_17174;
wire g57070_sb;
wire g57071_sb;
wire g57072_sb;
wire TIMEBOOST_net_10489;
wire g57073_sb;
wire TIMEBOOST_net_11922;
wire TIMEBOOST_net_22671;
wire g57074_sb;
wire TIMEBOOST_net_20539;
wire g57075_sb;
wire TIMEBOOST_net_22334;
wire g57076_sb;
wire TIMEBOOST_net_20318;
wire g57077_sb;
wire TIMEBOOST_net_16729;
wire g57078_sb;
wire TIMEBOOST_net_21193;
wire TIMEBOOST_net_10064;
wire g57079_sb;
wire TIMEBOOST_net_16399;
wire g57080_sb;
wire TIMEBOOST_net_22948;
wire g57081_sb;
wire TIMEBOOST_net_22896;
wire g57082_sb;
wire TIMEBOOST_net_21303;
wire TIMEBOOST_net_21409;
wire g57083_sb;
wire TIMEBOOST_net_23484;
wire TIMEBOOST_net_14413;
wire g57084_sb;
wire TIMEBOOST_net_20659;
wire TIMEBOOST_net_16401;
wire g57085_sb;
wire TIMEBOOST_net_21154;
wire g57086_sb;
wire g57087_sb;
wire TIMEBOOST_net_14471;
wire TIMEBOOST_net_17212;
wire g57088_sb;
wire TIMEBOOST_net_10541;
wire g57089_sb;
wire TIMEBOOST_net_21171;
wire g57090_sb;
wire g57091_sb;
wire TIMEBOOST_net_10517;
wire TIMEBOOST_net_14416;
wire g57092_sb;
wire g57093_sb;
wire TIMEBOOST_net_23313;
wire g57094_sb;
wire TIMEBOOST_net_12747;
wire TIMEBOOST_net_14418;
wire g57095_sb;
wire TIMEBOOST_net_16430;
wire g57096_sb;
wire TIMEBOOST_net_17044;
wire TIMEBOOST_net_14420;
wire g57097_sb;
wire TIMEBOOST_net_22928;
wire TIMEBOOST_net_14421;
wire g57098_sb;
wire g57099_sb;
wire TIMEBOOST_net_16405;
wire g57100_sb;
wire TIMEBOOST_net_10534;
wire TIMEBOOST_net_16406;
wire g57101_sb;
wire TIMEBOOST_net_10535;
wire TIMEBOOST_net_16407;
wire g57102_sb;
wire TIMEBOOST_net_10536;
wire TIMEBOOST_net_16408;
wire g57103_sb;
wire TIMEBOOST_net_23204;
wire TIMEBOOST_net_23270;
wire g57104_sb;
wire TIMEBOOST_net_22737;
wire TIMEBOOST_net_16409;
wire g57105_sb;
wire TIMEBOOST_net_17325;
wire g57106_sb;
wire g57107_sb;
wire TIMEBOOST_net_20555;
wire g57108_sb;
wire TIMEBOOST_net_16137;
wire g57109_sb;
wire TIMEBOOST_net_16411;
wire g57110_sb;
wire TIMEBOOST_net_14218;
wire TIMEBOOST_net_16138;
wire g57111_sb;
wire TIMEBOOST_net_20147;
wire TIMEBOOST_net_14675;
wire g57112_sb;
wire TIMEBOOST_net_23376;
wire TIMEBOOST_net_16412;
wire g57113_sb;
wire TIMEBOOST_net_16394;
wire g57114_sb;
wire TIMEBOOST_net_15349;
wire g57115_sb;
wire TIMEBOOST_net_23254;
wire g57116_sb;
wire TIMEBOOST_net_16730;
wire g57117_sb;
wire TIMEBOOST_net_21840;
wire TIMEBOOST_net_22955;
wire g57118_sb;
wire TIMEBOOST_net_6773;
wire TIMEBOOST_net_22445;
wire g57119_sb;
wire TIMEBOOST_net_21225;
wire TIMEBOOST_net_14407;
wire g57120_sb;
wire TIMEBOOST_net_16404;
wire g57121_sb;
wire TIMEBOOST_net_8776;
wire TIMEBOOST_net_20528;
wire g57122_sb;
wire TIMEBOOST_net_21194;
wire g57123_sb;
wire g57124_sb;
wire g57125_sb;
wire TIMEBOOST_net_21714;
wire g57126_sb;
wire TIMEBOOST_net_20342;
wire TIMEBOOST_net_23155;
wire g57127_sb;
wire TIMEBOOST_net_17127;
wire g57128_sb;
wire TIMEBOOST_net_21070;
wire g57129_sb;
wire TIMEBOOST_net_21227;
wire TIMEBOOST_net_16357;
wire g57130_sb;
wire g57131_sb;
wire g57132_sb;
wire TIMEBOOST_net_9478;
wire g57133_sb;
wire TIMEBOOST_net_13103;
wire TIMEBOOST_net_22854;
wire g57134_sb;
wire TIMEBOOST_net_13104;
wire TIMEBOOST_net_14398;
wire g57135_sb;
wire TIMEBOOST_net_10431;
wire g57136_sb;
wire TIMEBOOST_net_16140;
wire g57137_sb;
wire TIMEBOOST_net_9471;
wire g57138_sb;
wire TIMEBOOST_net_13106;
wire g57139_sb;
wire TIMEBOOST_net_23298;
wire g57140_sb;
wire g57141_sb;
wire TIMEBOOST_net_20529;
wire g57142_sb;
wire TIMEBOOST_net_14500;
wire g57143_sb;
wire TIMEBOOST_net_14596;
wire g57144_sb;
wire TIMEBOOST_net_10572;
wire TIMEBOOST_net_14388;
wire g57145_sb;
wire TIMEBOOST_net_14517;
wire TIMEBOOST_net_14100;
wire g57146_sb;
wire g57147_sb;
wire TIMEBOOST_net_21196;
wire g57148_sb;
wire TIMEBOOST_net_10424;
wire g57149_sb;
wire g57150_sb;
wire TIMEBOOST_net_10581;
wire TIMEBOOST_net_17457;
wire g57151_sb;
wire TIMEBOOST_net_10582;
wire g57152_sb;
wire TIMEBOOST_net_14157;
wire TIMEBOOST_net_16731;
wire g57153_sb;
wire TIMEBOOST_net_22492;
wire g57154_sb;
wire TIMEBOOST_net_10591;
wire g57155_sb;
wire g57156_sb;
wire g57157_sb;
wire g57158_sb;
wire TIMEBOOST_net_23222;
wire g57159_sb;
wire TIMEBOOST_net_15481;
wire g57160_sb;
wire TIMEBOOST_net_10566;
wire g57161_sb;
wire TIMEBOOST_net_10568;
wire TIMEBOOST_net_20607;
wire g57162_sb;
wire TIMEBOOST_net_11884;
wire g57163_sb;
wire TIMEBOOST_net_17292;
wire g57164_sb;
wire TIMEBOOST_net_10571;
wire g57165_sb;
wire g57166_sb;
wire TIMEBOOST_net_10569;
wire g59798_db;
wire g57167_sb;
wire TIMEBOOST_net_10354;
wire g57168_sb;
wire g57169_sb;
wire TIMEBOOST_net_17252;
wire TIMEBOOST_net_14322;
wire g57170_sb;
wire TIMEBOOST_net_21309;
wire TIMEBOOST_net_10353;
wire g57171_sb;
wire TIMEBOOST_net_6780;
wire TIMEBOOST_net_22477;
wire g57172_sb;
wire TIMEBOOST_net_10583;
wire g57173_sb;
wire TIMEBOOST_net_6781;
wire TIMEBOOST_net_20140;
wire g57174_sb;
wire TIMEBOOST_net_15391;
wire TIMEBOOST_net_22627;
wire g57175_sb;
wire TIMEBOOST_net_10567;
wire g57176_sb;
wire TIMEBOOST_net_23246;
wire TIMEBOOST_net_16332;
wire g57177_sb;
wire g57178_sb;
wire TIMEBOOST_net_22760;
wire g57179_sb;
wire TIMEBOOST_net_10577;
wire TIMEBOOST_net_17254;
wire g57180_sb;
wire TIMEBOOST_net_14158;
wire TIMEBOOST_net_10054;
wire g57181_sb;
wire TIMEBOOST_net_10576;
wire g57182_sb;
wire g57183_sb;
wire TIMEBOOST_net_21197;
wire TIMEBOOST_net_10063;
wire g57184_sb;
wire g57185_sb;
wire TIMEBOOST_net_20423;
wire g57186_sb;
wire TIMEBOOST_net_10062;
wire g57187_sb;
wire g57188_sb;
wire TIMEBOOST_net_16203;
wire TIMEBOOST_net_22587;
wire g57189_sb;
wire TIMEBOOST_net_10620;
wire g57190_sb;
wire TIMEBOOST_net_10562;
wire TIMEBOOST_net_17253;
wire g57191_sb;
wire TIMEBOOST_net_23171;
wire TIMEBOOST_net_17255;
wire g57192_sb;
wire TIMEBOOST_net_10615;
wire g57193_sb;
wire TIMEBOOST_net_21635;
wire g57194_sb;
wire TIMEBOOST_net_10179;
wire TIMEBOOST_net_10618;
wire g57195_sb;
wire TIMEBOOST_net_21735;
wire g57196_sb;
wire TIMEBOOST_net_10617;
wire g57197_sb;
wire TIMEBOOST_net_22469;
wire TIMEBOOST_net_15383;
wire g57198_sb;
wire TIMEBOOST_net_6785;
wire TIMEBOOST_net_22509;
wire g57199_sb;
wire g57200_sb;
wire TIMEBOOST_net_20588;
wire TIMEBOOST_net_10613;
wire g57201_sb;
wire g57202_sb;
wire TIMEBOOST_net_14167;
wire TIMEBOOST_net_10502;
wire g57203_sb;
wire TIMEBOOST_net_10520;
wire TIMEBOOST_net_10616;
wire g57204_sb;
wire TIMEBOOST_net_21473;
wire g57205_sb;
wire TIMEBOOST_net_10417;
wire TIMEBOOST_net_17102;
wire g57206_sb;
wire TIMEBOOST_net_6786;
wire g57207_sb;
wire TIMEBOOST_net_10416;
wire TIMEBOOST_net_15498;
wire g57208_sb;
wire TIMEBOOST_net_17521;
wire g57209_sb;
wire TIMEBOOST_net_16208;
wire TIMEBOOST_net_15345;
wire g57210_sb;
wire TIMEBOOST_net_10348;
wire TIMEBOOST_net_10280;
wire g57211_sb;
wire g57212_sb;
wire TIMEBOOST_net_21005;
wire TIMEBOOST_net_23282;
wire g57213_sb;
wire g57214_sb;
wire TIMEBOOST_net_23317;
wire TIMEBOOST_net_14373;
wire g57215_sb;
wire TIMEBOOST_net_8675;
wire g57216_sb;
wire TIMEBOOST_net_12471;
wire TIMEBOOST_net_16270;
wire g57217_sb;
wire TIMEBOOST_net_8677;
wire TIMEBOOST_net_23265;
wire g57218_sb;
wire TIMEBOOST_net_21198;
wire g57219_sb;
wire TIMEBOOST_net_12391;
wire g57220_sb;
wire TIMEBOOST_net_6789;
wire TIMEBOOST_net_22789;
wire g57221_sb;
wire TIMEBOOST_net_14147;
wire TIMEBOOST_net_10061;
wire g57222_sb;
wire TIMEBOOST_net_8741;
wire g57223_sb;
wire TIMEBOOST_net_22638;
wire g57224_sb;
wire TIMEBOOST_net_16934;
wire g57225_sb;
wire g57226_sb;
wire TIMEBOOST_net_17368;
wire g57227_sb;
wire g57228_sb;
wire TIMEBOOST_net_6792;
wire g57229_sb;
wire TIMEBOOST_net_6793;
wire TIMEBOOST_net_16166;
wire g57230_sb;
wire g57231_sb;
wire TIMEBOOST_net_6794;
wire TIMEBOOST_net_22687;
wire g57232_sb;
wire TIMEBOOST_net_16273;
wire g57233_sb;
wire TIMEBOOST_net_16973;
wire g57234_sb;
wire TIMEBOOST_net_16958;
wire TIMEBOOST_net_10281;
wire g57235_sb;
wire TIMEBOOST_net_14553;
wire TIMEBOOST_net_14222;
wire g57236_sb;
wire g52443_da;
wire TIMEBOOST_net_23202;
wire g57237_sb;
wire TIMEBOOST_net_10500;
wire g57238_sb;
wire TIMEBOOST_net_23305;
wire g57239_sb;
wire TIMEBOOST_net_20417;
wire TIMEBOOST_net_14223;
wire g57240_sb;
wire TIMEBOOST_net_13832;
wire TIMEBOOST_net_16274;
wire g57241_sb;
wire g57242_sb;
wire TIMEBOOST_net_22119;
wire TIMEBOOST_net_23237;
wire g57243_sb;
wire TIMEBOOST_net_10254;
wire TIMEBOOST_net_23241;
wire g57244_sb;
wire g57245_sb;
wire g57246_sb;
wire TIMEBOOST_net_23244;
wire g57247_sb;
wire TIMEBOOST_net_10407;
wire TIMEBOOST_net_14224;
wire g57248_sb;
wire TIMEBOOST_net_22476;
wire TIMEBOOST_net_23196;
wire g57249_sb;
wire TIMEBOOST_net_17330;
wire TIMEBOOST_net_20540;
wire g57250_sb;
wire g57251_sb;
wire g57252_sb;
wire g57253_sb;
wire TIMEBOOST_net_14722;
wire g57254_sb;
wire TIMEBOOST_net_20242;
wire g57255_sb;
wire TIMEBOOST_net_17105;
wire g57256_sb;
wire TIMEBOOST_net_23286;
wire g57257_sb;
wire TIMEBOOST_net_6802;
wire g57258_sb;
wire TIMEBOOST_net_6803;
wire g57259_sb;
wire TIMEBOOST_net_22496;
wire TIMEBOOST_net_21693;
wire g57260_sb;
wire TIMEBOOST_net_14233;
wire g57261_sb;
wire g57262_sb;
wire TIMEBOOST_net_14552;
wire g57263_sb;
wire TIMEBOOST_net_16184;
wire g57264_sb;
wire TIMEBOOST_net_17049;
wire TIMEBOOST_net_16185;
wire g57265_sb;
wire TIMEBOOST_net_21556;
wire TIMEBOOST_net_16186;
wire g57266_sb;
wire TIMEBOOST_net_21944;
wire g57267_sb;
wire TIMEBOOST_net_22689;
wire TIMEBOOST_net_14117;
wire g57268_sb;
wire TIMEBOOST_net_9587;
wire g57269_sb;
wire TIMEBOOST_net_10499;
wire g57270_sb;
wire TIMEBOOST_net_6805;
wire g57271_sb;
wire TIMEBOOST_net_6490;
wire TIMEBOOST_net_17106;
wire g57272_sb;
wire TIMEBOOST_net_14159;
wire g57273_sb;
wire TIMEBOOST_net_21658;
wire TIMEBOOST_net_16189;
wire g57274_sb;
wire g57275_sb;
wire n_9006;
wire TIMEBOOST_net_22872;
wire g57276_sb;
wire TIMEBOOST_net_10350;
wire g57277_sb;
wire TIMEBOOST_net_9571;
wire g57278_sb;
wire TIMEBOOST_net_21819;
wire TIMEBOOST_net_23211;
wire g57279_sb;
wire TIMEBOOST_net_12389;
wire g57280_sb;
wire TIMEBOOST_net_17241;
wire g57281_sb;
wire TIMEBOOST_net_12390;
wire TIMEBOOST_net_14057;
wire g57282_sb;
wire TIMEBOOST_net_6807;
wire TIMEBOOST_net_22327;
wire g57283_sb;
wire TIMEBOOST_net_6808;
wire TIMEBOOST_net_23192;
wire g57284_sb;
wire TIMEBOOST_net_23497;
wire g57285_sb;
wire TIMEBOOST_net_13099;
wire TIMEBOOST_net_16193;
wire g57286_sb;
wire TIMEBOOST_net_8728;
wire g57287_sb;
wire TIMEBOOST_net_17258;
wire TIMEBOOST_net_20183;
wire g57288_sb;
wire TIMEBOOST_net_22033;
wire g57289_sb;
wire TIMEBOOST_net_15097;
wire g57290_sb;
wire TIMEBOOST_net_6745;
wire g57291_sb;
wire TIMEBOOST_net_14971;
wire TIMEBOOST_net_22461;
wire g57292_sb;
wire TIMEBOOST_net_9584;
wire TIMEBOOST_net_16196;
wire g57293_sb;
wire TIMEBOOST_net_9585;
wire g57294_sb;
wire TIMEBOOST_net_9586;
wire g57295_sb;
wire TIMEBOOST_net_9582;
wire TIMEBOOST_net_16200;
wire g57296_sb;
wire TIMEBOOST_net_9607;
wire TIMEBOOST_net_16201;
wire g57297_sb;
wire TIMEBOOST_net_9580;
wire g57298_sb;
wire TIMEBOOST_net_9581;
wire TIMEBOOST_net_14162;
wire g57299_sb;
wire TIMEBOOST_net_10432;
wire TIMEBOOST_net_15519;
wire g57300_sb;
wire TIMEBOOST_net_9579;
wire g57301_sb;
wire TIMEBOOST_net_21823;
wire g57302_sb;
wire TIMEBOOST_net_9577;
wire g57303_sb;
wire TIMEBOOST_net_9578;
wire g57304_sb;
wire TIMEBOOST_net_9575;
wire TIMEBOOST_net_17117;
wire g57305_sb;
wire TIMEBOOST_net_21360;
wire g57306_sb;
wire TIMEBOOST_net_21981;
wire TIMEBOOST_net_17107;
wire g57307_sb;
wire TIMEBOOST_net_9564;
wire TIMEBOOST_net_14164;
wire g57308_sb;
wire TIMEBOOST_net_9565;
wire TIMEBOOST_net_17113;
wire g57309_sb;
wire TIMEBOOST_net_9566;
wire TIMEBOOST_net_16205;
wire g57310_sb;
wire TIMEBOOST_net_21988;
wire TIMEBOOST_net_14165;
wire g57311_sb;
wire TIMEBOOST_net_13542;
wire g57312_sb;
wire TIMEBOOST_net_22329;
wire g57313_sb;
wire TIMEBOOST_net_9568;
wire g57314_sb;
wire TIMEBOOST_net_6810;
wire TIMEBOOST_net_23113;
wire g57315_sb;
wire TIMEBOOST_net_6811;
wire TIMEBOOST_net_22388;
wire g57316_sb;
wire TIMEBOOST_net_9569;
wire g57317_sb;
wire TIMEBOOST_net_9570;
wire TIMEBOOST_net_14180;
wire g57318_sb;
wire TIMEBOOST_net_9572;
wire g57319_sb;
wire TIMEBOOST_net_17034;
wire g57320_sb;
wire TIMEBOOST_net_20419;
wire g57321_sb;
wire TIMEBOOST_net_17138;
wire g57322_sb;
wire TIMEBOOST_net_22767;
wire TIMEBOOST_net_6746;
wire g57323_sb;
wire TIMEBOOST_net_14562;
wire TIMEBOOST_net_22709;
wire g57324_sb;
wire TIMEBOOST_net_20158;
wire g57325_sb;
wire TIMEBOOST_net_13589;
wire TIMEBOOST_net_14225;
wire g57326_sb;
wire TIMEBOOST_net_23247;
wire g57327_sb;
wire TIMEBOOST_net_10052;
wire TIMEBOOST_net_20543;
wire g57328_sb;
wire g57329_sb;
wire TIMEBOOST_net_14860;
wire g57330_sb;
wire TIMEBOOST_net_16361;
wire g57331_sb;
wire TIMEBOOST_net_22460;
wire g57332_sb;
wire TIMEBOOST_net_17224;
wire TIMEBOOST_net_23223;
wire g57333_sb;
wire TIMEBOOST_net_13100;
wire TIMEBOOST_net_23224;
wire g57334_sb;
wire g57335_sb;
wire g57336_sb;
wire g57337_sb;
wire TIMEBOOST_net_20480;
wire g57338_sb;
wire TIMEBOOST_net_16290;
wire g57339_sb;
wire TIMEBOOST_net_6812;
wire TIMEBOOST_net_22392;
wire g57340_sb;
wire TIMEBOOST_net_6813;
wire g57341_sb;
wire TIMEBOOST_net_10637;
wire g57342_sb;
wire TIMEBOOST_net_10638;
wire g57343_sb;
wire TIMEBOOST_net_16293;
wire g57344_sb;
wire TIMEBOOST_net_22331;
wire g57345_sb;
wire TIMEBOOST_net_12551;
wire g57346_sb;
wire TIMEBOOST_net_10278;
wire g59230_db;
wire g57347_sb;
wire TIMEBOOST_net_10641;
wire TIMEBOOST_net_23228;
wire g57348_sb;
wire g57349_sb;
wire g57350_sb;
wire TIMEBOOST_net_17408;
wire g57351_sb;
wire TIMEBOOST_net_10645;
wire g57352_sb;
wire TIMEBOOST_net_20436;
wire TIMEBOOST_net_10060;
wire g57353_sb;
wire TIMEBOOST_net_21644;
wire TIMEBOOST_net_14226;
wire g57354_sb;
wire TIMEBOOST_net_10646;
wire TIMEBOOST_net_14227;
wire g57355_sb;
wire TIMEBOOST_net_22382;
wire g57356_sb;
wire TIMEBOOST_net_14228;
wire g57357_sb;
wire TIMEBOOST_net_10648;
wire g57358_sb;
wire TIMEBOOST_net_23421;
wire g57359_sb;
wire TIMEBOOST_net_12434;
wire TIMEBOOST_net_14230;
wire g57360_sb;
wire TIMEBOOST_net_23422;
wire g57361_sb;
wire TIMEBOOST_net_14231;
wire g57362_sb;
wire TIMEBOOST_net_23277;
wire g57363_sb;
wire TIMEBOOST_net_6817;
wire TIMEBOOST_net_22332;
wire g57364_sb;
wire TIMEBOOST_net_14232;
wire g57365_sb;
wire TIMEBOOST_net_9627;
wire TIMEBOOST_net_14381;
wire g57366_sb;
wire TIMEBOOST_net_6818;
wire TIMEBOOST_net_22333;
wire g57367_sb;
wire TIMEBOOST_net_9574;
wire g57368_sb;
wire TIMEBOOST_net_23257;
wire g57369_sb;
wire TIMEBOOST_net_22339;
wire TIMEBOOST_net_6747;
wire g57370_sb;
wire TIMEBOOST_net_22473;
wire TIMEBOOST_net_23424;
wire g57371_sb;
wire TIMEBOOST_net_12318;
wire g57372_sb;
wire g57373_sb;
wire TIMEBOOST_net_20542;
wire g57374_sb;
wire g57375_sb;
wire TIMEBOOST_net_12435;
wire TIMEBOOST_net_23331;
wire g57376_sb;
wire TIMEBOOST_net_6819;
wire TIMEBOOST_net_22395;
wire g57377_sb;
wire TIMEBOOST_net_20618;
wire g57378_sb;
wire TIMEBOOST_net_6820;
wire g57379_sb;
wire TIMEBOOST_net_15165;
wire TIMEBOOST_net_22417;
wire g57380_sb;
wire TIMEBOOST_net_16307;
wire g57381_sb;
wire TIMEBOOST_net_12450;
wire TIMEBOOST_net_16308;
wire g57382_sb;
wire TIMEBOOST_net_20177;
wire TIMEBOOST_net_14136;
wire g57383_sb;
wire TIMEBOOST_net_22658;
wire TIMEBOOST_net_20219;
wire g57384_sb;
wire TIMEBOOST_net_17315;
wire TIMEBOOST_net_20512;
wire g57385_sb;
wire TIMEBOOST_net_22676;
wire g57386_sb;
wire g57387_sb;
wire g57388_sb;
wire TIMEBOOST_net_9588;
wire g57389_sb;
wire TIMEBOOST_net_9649;
wire TIMEBOOST_net_16213;
wire g57390_sb;
wire TIMEBOOST_net_9650;
wire TIMEBOOST_net_23279;
wire g57391_sb;
wire TIMEBOOST_net_9651;
wire TIMEBOOST_net_17193;
wire g57392_sb;
wire TIMEBOOST_net_9652;
wire TIMEBOOST_net_23173;
wire g57393_sb;
wire g57394_sb;
wire g57395_sb;
wire TIMEBOOST_net_17058;
wire g57396_sb;
wire TIMEBOOST_net_9654;
wire TIMEBOOST_net_14170;
wire g57397_sb;
wire TIMEBOOST_net_21220;
wire g57398_sb;
wire TIMEBOOST_net_9656;
wire TIMEBOOST_net_20506;
wire g57399_sb;
wire TIMEBOOST_net_21677;
wire TIMEBOOST_net_14171;
wire g57400_sb;
wire TIMEBOOST_net_12032;
wire g57401_sb;
wire TIMEBOOST_net_6822;
wire g57402_sb;
wire TIMEBOOST_net_21719;
wire g57403_sb;
wire TIMEBOOST_net_10494;
wire g57404_sb;
wire g57405_sb;
wire g57406_sb;
wire TIMEBOOST_net_14172;
wire g57407_sb;
wire TIMEBOOST_net_23293;
wire g57408_sb;
wire TIMEBOOST_net_9662;
wire TIMEBOOST_net_20215;
wire g57409_sb;
wire TIMEBOOST_net_14561;
wire TIMEBOOST_net_20441;
wire g57410_sb;
wire TIMEBOOST_net_9663;
wire TIMEBOOST_net_20185;
wire g57411_sb;
wire TIMEBOOST_net_13627;
wire g57412_sb;
wire TIMEBOOST_net_22550;
wire TIMEBOOST_net_22402;
wire g57413_sb;
wire TIMEBOOST_net_22654;
wire g57414_sb;
wire g57415_sb;
wire TIMEBOOST_net_15818;
wire g57416_sb;
wire TIMEBOOST_net_16175;
wire g57417_sb;
wire TIMEBOOST_net_14177;
wire g57418_sb;
wire TIMEBOOST_net_12239;
wire TIMEBOOST_net_20207;
wire g57419_sb;
wire TIMEBOOST_net_9669;
wire TIMEBOOST_net_20447;
wire g57420_sb;
wire TIMEBOOST_net_20557;
wire TIMEBOOST_net_10059;
wire g57421_sb;
wire TIMEBOOST_net_22222;
wire g57422_sb;
wire TIMEBOOST_net_12275;
wire g57423_sb;
wire TIMEBOOST_net_22706;
wire TIMEBOOST_net_14179;
wire g57424_sb;
wire g57425_sb;
wire g57426_sb;
wire TIMEBOOST_net_15556;
wire g57427_sb;
wire TIMEBOOST_net_9573;
wire TIMEBOOST_net_14135;
wire g57428_sb;
wire TIMEBOOST_net_9473;
wire TIMEBOOST_net_20507;
wire g57429_sb;
wire TIMEBOOST_net_9475;
wire TIMEBOOST_net_23153;
wire g57430_sb;
wire TIMEBOOST_net_22377;
wire TIMEBOOST_net_23524;
wire g57431_sb;
wire TIMEBOOST_net_17316;
wire g57432_sb;
wire TIMEBOOST_net_9590;
wire g57433_sb;
wire TIMEBOOST_net_9591;
wire g57434_sb;
wire TIMEBOOST_net_9592;
wire g57435_sb;
wire TIMEBOOST_net_9593;
wire TIMEBOOST_net_14185;
wire g57436_sb;
wire TIMEBOOST_net_13609;
wire g57437_sb;
wire TIMEBOOST_net_9594;
wire TIMEBOOST_net_20464;
wire g57438_sb;
wire g57439_sb;
wire TIMEBOOST_net_9595;
wire g57440_sb;
wire TIMEBOOST_net_9596;
wire TIMEBOOST_net_23295;
wire g57441_sb;
wire TIMEBOOST_net_22399;
wire g57442_sb;
wire TIMEBOOST_net_9597;
wire TIMEBOOST_net_16232;
wire g57443_sb;
wire TIMEBOOST_net_6748;
wire g57444_sb;
wire TIMEBOOST_net_22341;
wire TIMEBOOST_net_6749;
wire g57445_sb;
wire g57446_sb;
wire TIMEBOOST_net_13610;
wire TIMEBOOST_net_22742;
wire g57447_sb;
wire TIMEBOOST_net_14125;
wire TIMEBOOST_net_17137;
wire g57448_sb;
wire g57449_sb;
wire TIMEBOOST_net_23312;
wire g57450_sb;
wire TIMEBOOST_net_14126;
wire g57451_sb;
wire TIMEBOOST_net_9598;
wire TIMEBOOST_net_20184;
wire g57452_sb;
wire TIMEBOOST_net_9599;
wire TIMEBOOST_net_20424;
wire g57453_sb;
wire TIMEBOOST_net_9600;
wire g57454_sb;
wire TIMEBOOST_net_9601;
wire g57455_sb;
wire TIMEBOOST_net_9603;
wire g57456_sb;
wire TIMEBOOST_net_16362;
wire TIMEBOOST_net_10058;
wire g57457_sb;
wire TIMEBOOST_net_9604;
wire g57458_sb;
wire TIMEBOOST_net_9605;
wire g57459_sb;
wire TIMEBOOST_net_9610;
wire g57460_sb;
wire TIMEBOOST_net_22389;
wire g57461_sb;
wire TIMEBOOST_net_9611;
wire TIMEBOOST_net_16237;
wire g57462_sb;
wire TIMEBOOST_net_9612;
wire TIMEBOOST_net_23259;
wire g57463_sb;
wire TIMEBOOST_net_21622;
wire TIMEBOOST_net_22383;
wire g57464_sb;
wire TIMEBOOST_net_9613;
wire TIMEBOOST_net_16238;
wire g57465_sb;
wire TIMEBOOST_net_9614;
wire TIMEBOOST_net_14191;
wire g57466_sb;
wire TIMEBOOST_net_9615;
wire TIMEBOOST_net_14192;
wire g57467_sb;
wire TIMEBOOST_net_22387;
wire g57468_sb;
wire g57469_sb;
wire g57470_sb;
wire TIMEBOOST_net_22862;
wire g57471_sb;
wire n_3684;
wire g57472_sb;
wire TIMEBOOST_net_14193;
wire g57473_sb;
wire TIMEBOOST_net_15338;
wire g57474_sb;
wire TIMEBOOST_net_22891;
wire g57475_sb;
wire TIMEBOOST_net_9618;
wire g57476_sb;
wire TIMEBOOST_net_9619;
wire TIMEBOOST_net_16240;
wire g57477_sb;
wire TIMEBOOST_net_16141;
wire TIMEBOOST_net_14702;
wire g57478_sb;
wire TIMEBOOST_net_14194;
wire g57479_sb;
wire TIMEBOOST_net_15073;
wire TIMEBOOST_net_16241;
wire g57480_sb;
wire TIMEBOOST_net_15071;
wire TIMEBOOST_net_14195;
wire g57481_sb;
wire TIMEBOOST_net_21446;
wire g57482_sb;
wire TIMEBOOST_net_21416;
wire TIMEBOOST_net_16176;
wire g57483_sb;
wire TIMEBOOST_net_14196;
wire g57484_sb;
wire TIMEBOOST_net_15439;
wire TIMEBOOST_net_10747;
wire g57485_sb;
wire TIMEBOOST_net_21454;
wire g57486_sb;
wire TIMEBOOST_net_11581;
wire TIMEBOOST_net_10748;
wire g57487_sb;
wire TIMEBOOST_net_16243;
wire g57488_sb;
wire TIMEBOOST_net_23079;
wire g57489_sb;
wire TIMEBOOST_net_21456;
wire g57490_sb;
wire TIMEBOOST_net_23294;
wire g57491_sb;
wire TIMEBOOST_net_21599;
wire TIMEBOOST_net_22697;
wire g57492_sb;
wire TIMEBOOST_net_21636;
wire g57493_sb;
wire TIMEBOOST_net_21713;
wire TIMEBOOST_net_16245;
wire g57494_sb;
wire TIMEBOOST_net_21774;
wire g57495_sb;
wire g57496_sb;
wire TIMEBOOST_net_22070;
wire g57497_sb;
wire TIMEBOOST_net_20530;
wire g57498_sb;
wire TIMEBOOST_net_21571;
wire TIMEBOOST_net_20531;
wire g57499_sb;
wire TIMEBOOST_net_21727;
wire TIMEBOOST_net_22930;
wire g57500_sb;
wire TIMEBOOST_net_16954;
wire g57501_sb;
wire TIMEBOOST_net_9644;
wire TIMEBOOST_net_14200;
wire g57502_sb;
wire TIMEBOOST_net_23016;
wire TIMEBOOST_net_23284;
wire g57503_sb;
wire TIMEBOOST_net_22999;
wire TIMEBOOST_net_16249;
wire g57504_sb;
wire TIMEBOOST_net_22967;
wire TIMEBOOST_net_21669;
wire g57505_sb;
wire TIMEBOOST_net_9647;
wire g57506_sb;
wire TIMEBOOST_net_9648;
wire TIMEBOOST_net_22947;
wire g57507_sb;
wire TIMEBOOST_net_23288;
wire g57508_sb;
wire TIMEBOOST_net_9602;
wire TIMEBOOST_net_14202;
wire g57509_sb;
wire TIMEBOOST_net_6750;
wire g57510_sb;
wire g57511_sb;
wire TIMEBOOST_net_20387;
wire TIMEBOOST_net_16251;
wire g57512_sb;
wire TIMEBOOST_net_17304;
wire TIMEBOOST_net_16252;
wire g57513_sb;
wire TIMEBOOST_net_14203;
wire g57514_sb;
wire TIMEBOOST_net_10717;
wire TIMEBOOST_net_23289;
wire g57515_sb;
wire TIMEBOOST_net_10718;
wire TIMEBOOST_net_16732;
wire TIMEBOOST_net_13710;
wire TIMEBOOST_net_16253;
wire g57517_sb;
wire g57518_sb;
wire n_3976;
wire TIMEBOOST_net_14204;
wire g57519_sb;
wire TIMEBOOST_net_10724;
wire g57520_sb;
wire g57521_sb;
wire TIMEBOOST_net_6845;
wire g57522_sb;
wire TIMEBOOST_net_16254;
wire g57523_sb;
wire TIMEBOOST_net_10742;
wire TIMEBOOST_net_20532;
wire g57524_sb;
wire g57525_sb;
wire TIMEBOOST_net_10721;
wire TIMEBOOST_net_20533;
wire g57526_sb;
wire TIMEBOOST_net_10727;
wire TIMEBOOST_net_20473;
wire g57527_sb;
wire TIMEBOOST_net_11886;
wire TIMEBOOST_net_9971;
wire g57528_sb;
wire TIMEBOOST_net_17110;
wire g57529_sb;
wire TIMEBOOST_net_17496;
wire TIMEBOOST_net_16259;
wire g57530_sb;
wire TIMEBOOST_net_17497;
wire g57531_sb;
wire TIMEBOOST_net_10746;
wire g57532_sb;
wire TIMEBOOST_net_17542;
wire TIMEBOOST_net_22436;
wire g57533_sb;
wire TIMEBOOST_net_10735;
wire g57534_sb;
wire TIMEBOOST_net_17498;
wire g57535_sb;
wire TIMEBOOST_net_6848;
wire g57536_sb;
wire TIMEBOOST_net_16143;
wire TIMEBOOST_net_6751;
wire g57537_sb;
wire TIMEBOOST_net_17499;
wire TIMEBOOST_net_16261;
wire g57538_sb;
wire TIMEBOOST_net_17500;
wire TIMEBOOST_net_23213;
wire g57539_sb;
wire TIMEBOOST_net_12648;
wire g57540_sb;
wire g57541_sb;
wire g62450_db;
wire g57542_sb;
wire TIMEBOOST_net_16144;
wire TIMEBOOST_net_16733;
wire g57543_sb;
wire TIMEBOOST_net_15487;
wire g57544_sb;
wire TIMEBOOST_net_23432;
wire TIMEBOOST_net_23209;
wire g57545_sb;
wire TIMEBOOST_net_16468;
wire g57546_sb;
wire TIMEBOOST_net_10464;
wire g57547_sb;
wire g57548_sb;
wire TIMEBOOST_net_10725;
wire TIMEBOOST_net_22468;
wire g57549_sb;
wire TIMEBOOST_net_14703;
wire g57550_sb;
wire TIMEBOOST_net_10726;
wire TIMEBOOST_net_20248;
wire g57551_sb;
wire TIMEBOOST_net_10728;
wire g57552_sb;
wire g57553_sb;
wire TIMEBOOST_net_11294;
wire TIMEBOOST_net_23197;
wire g57554_sb;
wire TIMEBOOST_net_20243;
wire g57555_sb;
wire TIMEBOOST_net_11345;
wire TIMEBOOST_net_22648;
wire g57556_sb;
wire TIMEBOOST_net_15501;
wire TIMEBOOST_net_6765;
wire g57557_sb;
wire g57558_sb;
wire TIMEBOOST_net_10262;
wire g57559_sb;
wire TIMEBOOST_net_23384;
wire TIMEBOOST_net_14214;
wire g57560_sb;
wire TIMEBOOST_net_15527;
wire TIMEBOOST_net_16983;
wire g57561_sb;
wire TIMEBOOST_net_21838;
wire g57562_sb;
wire TIMEBOOST_net_21758;
wire TIMEBOOST_net_22254;
wire g57563_sb;
wire TIMEBOOST_net_21389;
wire TIMEBOOST_net_20293;
wire g57564_sb;
wire TIMEBOOST_net_15693;
wire g57565_sb;
wire TIMEBOOST_net_22774;
wire g60664_db;
wire g57566_sb;
wire TIMEBOOST_net_16145;
wire TIMEBOOST_net_15717;
wire g57567_sb;
wire g65346_da;
wire g57568_sb;
wire g52460_da;
wire TIMEBOOST_net_22471;
wire g57569_sb;
wire TIMEBOOST_net_16265;
wire g57570_sb;
wire TIMEBOOST_net_16363;
wire g57571_sb;
wire TIMEBOOST_net_23505;
wire TIMEBOOST_net_23243;
wire g57572_sb;
wire TIMEBOOST_net_6860;
wire TIMEBOOST_net_23126;
wire g57573_sb;
wire TIMEBOOST_net_11369;
wire TIMEBOOST_net_12545;
wire g57574_sb;
wire TIMEBOOST_net_21393;
wire TIMEBOOST_net_16266;
wire g57575_sb;
wire TIMEBOOST_net_23229;
wire g57576_sb;
wire TIMEBOOST_net_23513;
wire TIMEBOOST_net_23203;
wire g57577_sb;
wire g57578_sb;
wire TIMEBOOST_net_21367;
wire TIMEBOOST_net_16268;
wire g57579_sb;
wire TIMEBOOST_net_22467;
wire g57580_sb;
wire TIMEBOOST_net_9942;
wire g57581_sb;
wire TIMEBOOST_net_22865;
wire TIMEBOOST_net_14217;
wire g57582_sb;
wire TIMEBOOST_net_6772;
wire g57583_sb;
wire g57584_sb;
wire TIMEBOOST_net_16734;
wire g57586_sb;
wire TIMEBOOST_net_11378;
wire g57587_sb;
wire TIMEBOOST_net_22879;
wire TIMEBOOST_net_21853;
wire g57588_sb;
wire TIMEBOOST_net_11379;
wire g57589_sb;
wire TIMEBOOST_net_11468;
wire TIMEBOOST_net_16269;
wire g57590_sb;
wire TIMEBOOST_net_14153;
wire TIMEBOOST_net_16309;
wire g57591_sb;
wire TIMEBOOST_net_11469;
wire g57592_sb;
wire TIMEBOOST_net_11470;
wire TIMEBOOST_net_14236;
wire g57593_sb;
wire TIMEBOOST_net_20631;
wire g57594_sb;
wire TIMEBOOST_net_17235;
wire g57595_sb;
wire TIMEBOOST_net_11472;
wire TIMEBOOST_net_16310;
wire g57596_sb;
wire TIMEBOOST_net_16311;
wire g57597_sb;
wire TIMEBOOST_net_21269;
wire g57598_sb;
wire TIMEBOOST_net_9405;
wire TIMEBOOST_net_16581;
wire TIMEBOOST_net_9499;
wire TIMEBOOST_net_10456;
wire g57780_sb;
wire TIMEBOOST_net_17225;
wire TIMEBOOST_net_17112;
wire TIMEBOOST_net_21351;
wire TIMEBOOST_net_10455;
wire TIMEBOOST_net_21354;
wire TIMEBOOST_net_10266;
wire g57787_da;
wire g57788_da;
wire TIMEBOOST_net_16364;
wire TIMEBOOST_net_16441;
wire TIMEBOOST_net_17194;
wire TIMEBOOST_net_21083;
wire TIMEBOOST_net_16381;
wire g57790_sb;
wire TIMEBOOST_net_16582;
wire TIMEBOOST_net_10627;
wire g57794_db;
wire g57794_sb;
wire TIMEBOOST_net_22291;
wire TIMEBOOST_net_16583;
wire g57795_sb;
wire TIMEBOOST_net_22292;
wire TIMEBOOST_net_21350;
wire TIMEBOOST_net_22288;
wire TIMEBOOST_net_16541;
wire g57797_sb;
wire TIMEBOOST_net_16039;
wire TIMEBOOST_net_20322;
wire TIMEBOOST_net_16040;
wire TIMEBOOST_net_16584;
wire TIMEBOOST_net_13670;
wire TIMEBOOST_net_20323;
wire TIMEBOOST_net_22283;
wire TIMEBOOST_net_10707;
wire TIMEBOOST_net_16029;
wire g57856_p;
wire g57863_p;
wire g57864_p;
wire g57875_sb;
wire g57876_p;
wire g57878_p;
wire TIMEBOOST_net_17043;
wire g57890_sb;
wire g61968_db;
wire g57891_db;
wire g57891_sb;
wire g61962_db;
wire g57892_db;
wire g57892_sb;
wire TIMEBOOST_net_14260;
wire g57893_db;
wire g57893_sb;
wire TIMEBOOST_net_22293;
wire g57894_db;
wire g57894_sb;
wire g61923_db;
wire g57895_db;
wire g57895_sb;
wire TIMEBOOST_net_17139;
wire g57896_sb;
wire TIMEBOOST_net_13578;
wire g57897_db;
wire g57897_sb;
wire g57898_db;
wire g57898_sb;
wire g57899_db;
wire g57899_sb;
wire TIMEBOOST_net_17067;
wire g57900_sb;
wire TIMEBOOST_net_21647;
wire g57901_db;
wire g57901_sb;
wire TIMEBOOST_net_9406;
wire g57902_sb;
wire TIMEBOOST_net_13692;
wire g57903_sb;
wire TIMEBOOST_net_13577;
wire g57904_db;
wire g57904_sb;
wire TIMEBOOST_net_23536;
wire g57905_sb;
wire TIMEBOOST_net_13586;
wire g57906_db;
wire g57906_sb;
wire g57907_db;
wire g57907_sb;
wire g57908_sb;
wire g57909_db;
wire g57909_sb;
wire TIMEBOOST_net_14779;
wire g57910_sb;
wire TIMEBOOST_net_22122;
wire g57911_db;
wire g57911_sb;
wire g57912_db;
wire g57912_sb;
wire TIMEBOOST_net_12690;
wire TIMEBOOST_net_17319;
wire g57913_sb;
wire TIMEBOOST_net_17140;
wire g57914_sb;
wire TIMEBOOST_net_17141;
wire g57915_sb;
wire TIMEBOOST_net_17142;
wire g57916_sb;
wire TIMEBOOST_net_17143;
wire g57917_sb;
wire TIMEBOOST_net_14087;
wire g57918_sb;
wire TIMEBOOST_net_14038;
wire g57919_db;
wire g57919_sb;
wire TIMEBOOST_net_21327;
wire g57920_db;
wire g57920_sb;
wire TIMEBOOST_net_22270;
wire TIMEBOOST_net_17229;
wire g57921_sb;
wire TIMEBOOST_net_22271;
wire g57922_db;
wire g57922_sb;
wire g57923_db;
wire g57923_sb;
wire g57924_db;
wire g57924_sb;
wire TIMEBOOST_net_14849;
wire TIMEBOOST_net_17144;
wire g57925_sb;
wire TIMEBOOST_net_14011;
wire g57926_db;
wire g57926_sb;
wire g57927_db;
wire g57927_sb;
wire TIMEBOOST_net_13964;
wire TIMEBOOST_net_22630;
wire g57928_sb;
wire TIMEBOOST_net_9323;
wire g57929_db;
wire g57929_sb;
wire TIMEBOOST_net_13745;
wire g57930_db;
wire g57930_sb;
wire TIMEBOOST_net_13742;
wire TIMEBOOST_net_17145;
wire g57931_sb;
wire TIMEBOOST_net_14021;
wire TIMEBOOST_net_12263;
wire g57932_sb;
wire TIMEBOOST_net_13851;
wire TIMEBOOST_net_17146;
wire g57933_sb;
wire TIMEBOOST_net_10528;
wire g57934_sb;
wire TIMEBOOST_net_13848;
wire g57935_db;
wire g57935_sb;
wire TIMEBOOST_net_17147;
wire g57936_sb;
wire TIMEBOOST_net_13847;
wire TIMEBOOST_net_21055;
wire g57937_sb;
wire TIMEBOOST_net_13846;
wire g57938_db;
wire g57938_sb;
wire TIMEBOOST_net_17149;
wire g57939_sb;
wire TIMEBOOST_net_13743;
wire g57940_db;
wire g57940_sb;
wire TIMEBOOST_net_21406;
wire g57941_db;
wire g57941_sb;
wire TIMEBOOST_net_13845;
wire TIMEBOOST_net_17151;
wire g57942_sb;
wire TIMEBOOST_net_13843;
wire g57944_db;
wire g57944_sb;
wire TIMEBOOST_net_13792;
wire g57945_db;
wire g57945_sb;
wire TIMEBOOST_net_14205;
wire TIMEBOOST_net_17155;
wire g57946_sb;
wire TIMEBOOST_net_13380;
wire TIMEBOOST_net_15557;
wire g57947_sb;
wire TIMEBOOST_net_14828;
wire g57948_db;
wire g57948_sb;
wire TIMEBOOST_net_13744;
wire TIMEBOOST_net_22128;
wire g57949_sb;
wire n_4307;
wire g57950_db;
wire TIMEBOOST_net_17363;
wire g57951_db;
wire g57951_sb;
wire g57952_db;
wire g57952_sb;
wire TIMEBOOST_net_16329;
wire g57953_db;
wire g57953_sb;
wire TIMEBOOST_net_14261;
wire g57954_db;
wire g57954_sb;
wire TIMEBOOST_net_20735;
wire g57955_db;
wire TIMEBOOST_net_20786;
wire g57956_db;
wire g57956_sb;
wire g65763_da;
wire g57957_db;
wire g57957_sb;
wire g57958_db;
wire g57958_sb;
wire TIMEBOOST_net_14255;
wire g57959_sb;
wire TIMEBOOST_net_13970;
wire g57960_db;
wire g57961_db;
wire g57961_sb;
wire g57962_db;
wire TIMEBOOST_net_14263;
wire TIMEBOOST_net_17158;
wire TIMEBOOST_net_8387;
wire TIMEBOOST_net_17159;
wire g57964_sb;
wire TIMEBOOST_net_13617;
wire g57965_db;
wire g57965_sb;
wire TIMEBOOST_net_14880;
wire TIMEBOOST_net_11386;
wire TIMEBOOST_net_22374;
wire TIMEBOOST_net_22140;
wire TIMEBOOST_net_14264;
wire g57968_db;
wire g57968_sb;
wire g57969_sb;
wire g57970_db;
wire g57970_sb;
wire TIMEBOOST_net_20138;
wire g57971_sb;
wire TIMEBOOST_net_17162;
wire g57972_sb;
wire TIMEBOOST_net_20286;
wire g57973_db;
wire g57973_sb;
wire TIMEBOOST_net_17163;
wire TIMEBOOST_net_17164;
wire g57975_sb;
wire g57976_db;
wire TIMEBOOST_net_13448;
wire TIMEBOOST_net_17119;
wire g57977_sb;
wire TIMEBOOST_net_22597;
wire TIMEBOOST_net_12242;
wire g57978_sb;
wire TIMEBOOST_net_14941;
wire g57979_db;
wire g57979_sb;
wire TIMEBOOST_net_15024;
wire TIMEBOOST_net_17268;
wire g57980_sb;
wire TIMEBOOST_net_13449;
wire g57981_db;
wire g57981_sb;
wire g57982_db;
wire g57982_sb;
wire TIMEBOOST_net_13450;
wire g57983_db;
wire g57983_sb;
wire g57984_db;
wire g57984_sb;
wire TIMEBOOST_net_15657;
wire g57985_db;
wire g57985_sb;
wire TIMEBOOST_net_17120;
wire g57986_sb;
wire TIMEBOOST_net_14891;
wire g57987_db;
wire g57987_sb;
wire g57988_sb;
wire g57989_db;
wire g57989_sb;
wire TIMEBOOST_net_22202;
wire TIMEBOOST_net_17121;
wire g57990_sb;
wire TIMEBOOST_net_20906;
wire g57991_sb;
wire TIMEBOOST_net_21247;
wire g57992_db;
wire g57992_sb;
wire g57993_db;
wire g57993_sb;
wire TIMEBOOST_net_17562;
wire TIMEBOOST_net_17269;
wire g57994_sb;
wire TIMEBOOST_net_17122;
wire g57995_sb;
wire g57996_db;
wire g57996_sb;
wire g57997_db;
wire g57997_sb;
wire TIMEBOOST_net_17563;
wire g57998_db;
wire TIMEBOOST_net_17123;
wire g57999_sb;
wire TIMEBOOST_net_13688;
wire g58000_db;
wire g58000_sb;
wire TIMEBOOST_net_14929;
wire g58001_sb;
wire g58002_sb;
wire TIMEBOOST_net_20365;
wire g58003_db;
wire g58003_sb;
wire TIMEBOOST_net_13707;
wire g58004_sb;
wire TIMEBOOST_net_17293;
wire g58005_sb;
wire TIMEBOOST_net_13706;
wire g58006_db;
wire g58006_sb;
wire TIMEBOOST_net_14434;
wire TIMEBOOST_net_17165;
wire g58008_sb;
wire g58009_db;
wire g58009_sb;
wire TIMEBOOST_net_12276;
wire g58010_db;
wire g58010_sb;
wire TIMEBOOST_net_16587;
wire TIMEBOOST_net_17068;
wire g58011_sb;
wire TIMEBOOST_net_17388;
wire TIMEBOOST_net_21577;
wire g58012_sb;
wire TIMEBOOST_net_23506;
wire g58013_db;
wire g58013_sb;
wire g58014_db;
wire g58014_sb;
wire TIMEBOOST_net_22465;
wire g58015_db;
wire g58015_sb;
wire TIMEBOOST_net_14519;
wire g58016_sb;
wire g58017_sb;
wire g58018_db;
wire g58018_sb;
wire TIMEBOOST_net_21127;
wire g58019_db;
wire g58019_sb;
wire g58020_db;
wire g58020_sb;
wire TIMEBOOST_net_16657;
wire TIMEBOOST_net_17069;
wire g58021_sb;
wire TIMEBOOST_net_13971;
wire TIMEBOOST_net_21580;
wire g58022_sb;
wire g63091_db;
wire g58023_db;
wire g58023_sb;
wire TIMEBOOST_net_17070;
wire g58024_sb;
wire TIMEBOOST_net_8343;
wire g58025_sb;
wire TIMEBOOST_net_21292;
wire TIMEBOOST_net_21694;
wire g58026_sb;
wire g58027_db;
wire g58027_sb;
wire g58028_db;
wire g58028_sb;
wire TIMEBOOST_net_14547;
wire TIMEBOOST_net_22867;
wire g58029_sb;
wire g58030_sb;
wire TIMEBOOST_net_17071;
wire g58031_sb;
wire TIMEBOOST_net_21040;
wire g58032_db;
wire g58032_sb;
wire g63089_db;
wire g58033_db;
wire g58033_sb;
wire TIMEBOOST_net_17370;
wire g58034_db;
wire g58034_sb;
wire TIMEBOOST_net_17072;
wire g58035_sb;
wire TIMEBOOST_net_20249;
wire TIMEBOOST_net_17073;
wire g58036_sb;
wire TIMEBOOST_net_12682;
wire g58037_db;
wire g58037_sb;
wire g58038_db;
wire TIMEBOOST_net_13952;
wire g58039_db;
wire g58039_sb;
wire TIMEBOOST_net_21200;
wire g58040_db;
wire g58040_sb;
wire g58041_db;
wire g58041_sb;
wire TIMEBOOST_net_187;
wire TIMEBOOST_net_23163;
wire g58042_sb;
wire TIMEBOOST_net_8336;
wire g58043_db;
wire g58043_sb;
wire TIMEBOOST_net_21291;
wire g58044_db;
wire g58044_sb;
wire TIMEBOOST_net_8334;
wire g58045_db;
wire g58045_sb;
wire TIMEBOOST_net_23423;
wire g58046_db;
wire g58046_sb;
wire TIMEBOOST_net_21177;
wire g58047_sb;
wire g58048_db;
wire g58048_sb;
wire TIMEBOOST_net_20742;
wire g58049_db;
wire g58049_sb;
wire TIMEBOOST_net_21290;
wire g58050_db;
wire g58050_sb;
wire g63056_db;
wire g58051_db;
wire g58051_sb;
wire g58052_sb;
wire TIMEBOOST_net_21934;
wire g58053_sb;
wire TIMEBOOST_net_180;
wire g58054_db;
wire TIMEBOOST_net_8332;
wire TIMEBOOST_net_21935;
wire g58055_sb;
wire TIMEBOOST_net_21267;
wire g58056_db;
wire g58056_sb;
wire TIMEBOOST_net_8331;
wire g58057_db;
wire g58057_sb;
wire g58058_db;
wire g58058_sb;
wire TIMEBOOST_net_12488;
wire g58059_sb;
wire TIMEBOOST_net_21559;
wire g58060_sb;
wire TIMEBOOST_net_15582;
wire g58061_db;
wire g58062_db;
wire g58062_sb;
wire g63052_db;
wire g58063_db;
wire g58063_sb;
wire g58064_db;
wire TIMEBOOST_net_22763;
wire TIMEBOOST_net_12681;
wire g58066_db;
wire g58066_sb;
wire g58067_db;
wire TIMEBOOST_net_14826;
wire g58068_sb;
wire g58069_sb;
wire TIMEBOOST_net_20885;
wire g58070_sb;
wire TIMEBOOST_net_21817;
wire g58071_db;
wire g58071_sb;
wire TIMEBOOST_net_14292;
wire TIMEBOOST_net_20599;
wire g58072_sb;
wire TIMEBOOST_net_8325;
wire TIMEBOOST_net_16605;
wire g58073_sb;
wire TIMEBOOST_net_8324;
wire g58074_db;
wire g58074_sb;
wire g58075_sb;
wire g58076_db;
wire g58076_sb;
wire TIMEBOOST_net_22190;
wire g58077_db;
wire g58077_sb;
wire g58078_db;
wire g58078_sb;
wire TIMEBOOST_net_17047;
wire g58079_sb;
wire TIMEBOOST_net_8322;
wire g58080_db;
wire g58080_sb;
wire g58081_db;
wire g58081_sb;
wire TIMEBOOST_net_13800;
wire g58082_db;
wire g58082_sb;
wire g58083_db;
wire g58083_sb;
wire g63013_db;
wire g58084_db;
wire g58084_sb;
wire g58085_db;
wire g58086_sb;
wire g58087_db;
wire g58087_sb;
wire g58088_db;
wire g58088_sb;
wire g58089_db;
wire g58089_sb;
wire g58090_db;
wire g58090_sb;
wire TIMEBOOST_net_13386;
wire TIMEBOOST_net_21718;
wire g58091_sb;
wire TIMEBOOST_net_12679;
wire g58092_db;
wire g58092_sb;
wire g58093_sb;
wire TIMEBOOST_net_14293;
wire g58094_db;
wire g58094_sb;
wire g62852_db;
wire g58095_db;
wire g58095_sb;
wire TIMEBOOST_net_23544;
wire TIMEBOOST_net_17048;
wire g58096_sb;
wire TIMEBOOST_net_14571;
wire g58097_db;
wire g58097_sb;
wire g58098_db;
wire TIMEBOOST_net_8316;
wire g58099_db;
wire g58099_sb;
wire TIMEBOOST_net_21448;
wire TIMEBOOST_net_14151;
wire g58100_sb;
wire TIMEBOOST_net_22052;
wire TIMEBOOST_net_17074;
wire g58101_sb;
wire g62843_db;
wire g58102_db;
wire g58102_sb;
wire TIMEBOOST_net_14435;
wire g58103_sb;
wire TIMEBOOST_net_14436;
wire TIMEBOOST_net_6961;
wire g58104_sb;
wire TIMEBOOST_net_8109;
wire g58105_db;
wire g58105_sb;
wire TIMEBOOST_net_21626;
wire TIMEBOOST_net_22590;
wire g58106_sb;
wire g58107_db;
wire g58107_sb;
wire TIMEBOOST_net_22080;
wire TIMEBOOST_net_22540;
wire g58108_sb;
wire g62833_db;
wire TIMEBOOST_net_17004;
wire TIMEBOOST_net_22045;
wire g58110_sb;
wire TIMEBOOST_net_22020;
wire g58111_db;
wire g58111_sb;
wire TIMEBOOST_net_21707;
wire g58112_db;
wire g58112_sb;
wire g62811_db;
wire g58113_db;
wire g58113_sb;
wire g58114_sb;
wire g58115_sb;
wire g58116_db;
wire g58116_sb;
wire TIMEBOOST_net_14822;
wire g58117_sb;
wire TIMEBOOST_net_21673;
wire g58118_sb;
wire g62803_db;
wire g58119_sb;
wire TIMEBOOST_net_13797;
wire TIMEBOOST_net_17133;
wire g58120_sb;
wire TIMEBOOST_net_12257;
wire g58121_db;
wire g58122_db;
wire TIMEBOOST_net_182;
wire TIMEBOOST_net_10425;
wire g58123_sb;
wire TIMEBOOST_net_306;
wire g58124_sb;
wire TIMEBOOST_net_21536;
wire g58125_sb;
wire TIMEBOOST_net_12256;
wire g58126_db;
wire g58126_sb;
wire g58127_sb;
wire g58128_db;
wire g58128_sb;
wire TIMEBOOST_net_17005;
wire g58129_sb;
wire TIMEBOOST_net_17393;
wire g58130_db;
wire g58130_sb;
wire TIMEBOOST_net_20724;
wire TIMEBOOST_net_22541;
wire n_9735;
wire g58132_db;
wire g58132_sb;
wire TIMEBOOST_net_14296;
wire g58133_db;
wire g58133_sb;
wire TIMEBOOST_net_23404;
wire TIMEBOOST_net_178;
wire TIMEBOOST_net_183;
wire TIMEBOOST_net_8311;
wire TIMEBOOST_net_22183;
wire g58136_sb;
wire TIMEBOOST_net_17392;
wire g58137_db;
wire g58138_db;
wire g58138_sb;
wire TIMEBOOST_net_14842;
wire g58139_db;
wire g58139_sb;
wire TIMEBOOST_net_15554;
wire g58140_db;
wire g58140_sb;
wire g58141_db;
wire g58141_sb;
wire g58142_db;
wire g58142_sb;
wire g58143_db;
wire g58143_sb;
wire TIMEBOOST_net_12650;
wire g58144_db;
wire g58144_sb;
wire TIMEBOOST_net_16588;
wire g58145_db;
wire g58145_sb;
wire TIMEBOOST_net_16589;
wire g58146_db;
wire g58146_sb;
wire TIMEBOOST_net_14856;
wire g58147_db;
wire g58147_sb;
wire TIMEBOOST_net_14952;
wire g58148_db;
wire g58148_sb;
wire TIMEBOOST_net_12255;
wire g58149_db;
wire g58149_sb;
wire g58150_sb;
wire TIMEBOOST_net_14690;
wire g58151_db;
wire TIMEBOOST_net_13801;
wire TIMEBOOST_net_21604;
wire g58152_sb;
wire TIMEBOOST_net_21270;
wire g58153_db;
wire g58153_sb;
wire TIMEBOOST_net_16590;
wire g58154_db;
wire g58154_sb;
wire g58155_db;
wire TIMEBOOST_net_23430;
wire TIMEBOOST_net_17075;
wire g58156_sb;
wire TIMEBOOST_net_13953;
wire TIMEBOOST_net_17076;
wire TIMEBOOST_net_14947;
wire g58158_db;
wire g58158_sb;
wire TIMEBOOST_net_13226;
wire g58159_db;
wire g58159_sb;
wire g58160_db;
wire g58160_sb;
wire g58161_sb;
wire TIMEBOOST_net_12641;
wire g58162_db;
wire g58162_sb;
wire TIMEBOOST_net_22695;
wire g58163_sb;
wire TIMEBOOST_net_16667;
wire TIMEBOOST_net_17077;
wire g58164_sb;
wire TIMEBOOST_net_16670;
wire g58165_db;
wire g58165_sb;
wire g58166_db;
wire TIMEBOOST_net_17078;
wire g58167_sb;
wire g58168_db;
wire TIMEBOOST_net_10516;
wire g58169_sb;
wire TIMEBOOST_net_14726;
wire g58170_db;
wire g58170_sb;
wire g58171_db;
wire g58171_sb;
wire g58172_sb;
wire TIMEBOOST_net_23541;
wire g58173_db;
wire g58173_sb;
wire g58382_da;
wire g58174_db;
wire g58174_sb;
wire g58175_db;
wire g58175_sb;
wire g58176_db;
wire g58176_sb;
wire TIMEBOOST_net_20880;
wire g58177_db;
wire g58177_sb;
wire FE_RN_579_0;
wire g58178_sb;
wire TIMEBOOST_net_23545;
wire g58179_db;
wire g58179_sb;
wire TIMEBOOST_net_20362;
wire g58180_sb;
wire TIMEBOOST_net_21849;
wire g58181_sb;
wire TIMEBOOST_net_15558;
wire g58182_sb;
wire TIMEBOOST_net_14438;
wire g58183_db;
wire g58183_sb;
wire TIMEBOOST_net_20288;
wire g58184_sb;
wire g64319_db;
wire TIMEBOOST_net_15401;
wire g58185_sb;
wire TIMEBOOST_net_17387;
wire g58186_sb;
wire TIMEBOOST_net_15692;
wire g58187_db;
wire g58187_sb;
wire TIMEBOOST_net_13090;
wire g58188_sb;
wire TIMEBOOST_net_17171;
wire g58189_sb;
wire TIMEBOOST_net_12634;
wire g58190_db;
wire g58190_sb;
wire TIMEBOOST_net_20363;
wire g58191_db;
wire g58191_sb;
wire g58192_sb;
wire g58193_db;
wire g58193_sb;
wire TIMEBOOST_net_17172;
wire g58194_sb;
wire TIMEBOOST_net_14441;
wire TIMEBOOST_net_17173;
wire g58195_sb;
wire TIMEBOOST_net_20608;
wire g58196_sb;
wire TIMEBOOST_net_15882;
wire g58197_db;
wire g58197_sb;
wire g58198_db;
wire g58198_sb;
wire g58199_db;
wire g58199_sb;
wire g58200_db;
wire g58200_sb;
wire g61958_db;
wire g58201_db;
wire g58201_sb;
wire g58202_db;
wire g58202_sb;
wire TIMEBOOST_net_12625;
wire g58203_db;
wire g58203_sb;
wire TIMEBOOST_net_12624;
wire g58204_db;
wire g58204_sb;
wire TIMEBOOST_net_16719;
wire g58205_sb;
wire TIMEBOOST_net_21011;
wire TIMEBOOST_net_14576;
wire g58206_sb;
wire g58207_db;
wire g58207_sb;
wire TIMEBOOST_net_14775;
wire g58208_db;
wire g58208_sb;
wire g58209_db;
wire g58209_sb;
wire TIMEBOOST_net_21994;
wire g58210_db;
wire g58210_sb;
wire TIMEBOOST_net_22336;
wire g58211_sb;
wire TIMEBOOST_net_23329;
wire g58212_sb;
wire TIMEBOOST_net_14593;
wire g58213_db;
wire g58213_sb;
wire g58214_db;
wire g58214_sb;
wire TIMEBOOST_net_12622;
wire g58215_sb;
wire TIMEBOOST_net_21000;
wire TIMEBOOST_net_22807;
wire g58216_sb;
wire TIMEBOOST_net_14946;
wire g58217_db;
wire g58217_sb;
wire TIMEBOOST_net_12620;
wire TIMEBOOST_net_15387;
wire g58218_sb;
wire g58219_db;
wire g58219_sb;
wire TIMEBOOST_net_17079;
wire g58220_sb;
wire TIMEBOOST_net_17381;
wire g58221_sb;
wire g58222_db;
wire g58222_sb;
wire g58223_db;
wire g58223_sb;
wire TIMEBOOST_net_20537;
wire g58224_db;
wire g58224_sb;
wire TIMEBOOST_net_17380;
wire g58225_db;
wire g58225_sb;
wire TIMEBOOST_net_20525;
wire TIMEBOOST_net_17080;
wire g58227_db;
wire g58227_sb;
wire TIMEBOOST_net_8289;
wire g58228_db;
wire g58228_sb;
wire g58229_db;
wire g58229_sb;
wire TIMEBOOST_net_14442;
wire TIMEBOOST_net_17176;
wire g58230_sb;
wire TIMEBOOST_net_8108;
wire TIMEBOOST_net_12933;
wire g58231_sb;
wire TIMEBOOST_net_8288;
wire TIMEBOOST_net_22243;
wire g58232_sb;
wire g58233_db;
wire g58233_sb;
wire TIMEBOOST_net_22030;
wire g58234_db;
wire g58234_sb;
wire TIMEBOOST_net_8107;
wire TIMEBOOST_net_21697;
wire g58235_sb;
wire TIMEBOOST_net_14443;
wire TIMEBOOST_net_22240;
wire g58236_sb;
wire g58237_sb;
wire TIMEBOOST_net_14837;
wire g58238_sb;
wire g58239_sb;
wire TIMEBOOST_net_13539;
wire TIMEBOOST_net_16972;
wire g58240_sb;
wire TIMEBOOST_net_21952;
wire g58241_db;
wire TIMEBOOST_net_8105;
wire TIMEBOOST_net_21169;
wire g58242_sb;
wire TIMEBOOST_net_13789;
wire g58243_db;
wire g58243_sb;
wire TIMEBOOST_net_9324;
wire g58244_sb;
wire TIMEBOOST_net_22047;
wire g58245_db;
wire TIMEBOOST_net_16463;
wire TIMEBOOST_net_22237;
wire TIMEBOOST_net_21458;
wire TIMEBOOST_net_12618;
wire g58248_db;
wire TIMEBOOST_net_13607;
wire g58249_db;
wire TIMEBOOST_net_14594;
wire g58251_db;
wire g58251_sb;
wire TIMEBOOST_net_21253;
wire g58252_sb;
wire TIMEBOOST_net_13545;
wire TIMEBOOST_net_10380;
wire TIMEBOOST_net_8104;
wire g58254_sb;
wire g58255_db;
wire g58255_sb;
wire TIMEBOOST_net_22014;
wire TIMEBOOST_net_22238;
wire g58256_sb;
wire TIMEBOOST_net_20280;
wire TIMEBOOST_net_22257;
wire g58257_sb;
wire TIMEBOOST_net_8103;
wire g58258_db;
wire g58258_sb;
wire TIMEBOOST_net_8272;
wire TIMEBOOST_net_13537;
wire g58260_db;
wire g58260_sb;
wire TIMEBOOST_net_9480;
wire TIMEBOOST_net_10131;
wire g58261_sb;
wire TIMEBOOST_net_22581;
wire TIMEBOOST_net_15488;
wire g58262_sb;
wire TIMEBOOST_net_15807;
wire g58263_sb;
wire TIMEBOOST_net_13803;
wire TIMEBOOST_net_17248;
wire g58264_sb;
wire TIMEBOOST_net_12619;
wire TIMEBOOST_net_20642;
wire g58265_sb;
wire TIMEBOOST_net_12817;
wire g58266_sb;
wire TIMEBOOST_net_17249;
wire g58267_sb;
wire TIMEBOOST_net_13585;
wire g58268_db;
wire g58268_sb;
wire TIMEBOOST_net_13576;
wire g58269_db;
wire g58269_sb;
wire TIMEBOOST_net_15667;
wire g58270_sb;
wire TIMEBOOST_net_20443;
wire TIMEBOOST_net_15342;
wire g58271_sb;
wire TIMEBOOST_net_21275;
wire TIMEBOOST_net_7726;
wire g58272_sb;
wire TIMEBOOST_net_14763;
wire TIMEBOOST_net_13538;
wire g58273_sb;
wire TIMEBOOST_net_22037;
wire g58274_sb;
wire g58275_sb;
wire TIMEBOOST_net_16513;
wire g58276_db;
wire g58276_sb;
wire TIMEBOOST_net_13835;
wire g58277_db;
wire g58277_sb;
wire TIMEBOOST_net_13844;
wire g58278_db;
wire g58278_sb;
wire TIMEBOOST_net_13842;
wire TIMEBOOST_net_17441;
wire g58279_sb;
wire n_13175;
wire TIMEBOOST_net_21841;
wire g58280_sb;
wire g58281_sb;
wire TIMEBOOST_net_14861;
wire g58282_sb;
wire TIMEBOOST_net_13841;
wire g58283_db;
wire g58283_sb;
wire TIMEBOOST_net_13840;
wire TIMEBOOST_net_16663;
wire g58284_sb;
wire TIMEBOOST_net_17586;
wire TIMEBOOST_net_21730;
wire g58285_sb;
wire TIMEBOOST_net_14685;
wire g58286_sb;
wire TIMEBOOST_net_13839;
wire g58287_db;
wire g58287_sb;
wire TIMEBOOST_net_13838;
wire TIMEBOOST_net_22058;
wire g58288_sb;
wire TIMEBOOST_net_13837;
wire g58289_sb;
wire TIMEBOOST_net_13836;
wire g58290_db;
wire g58290_sb;
wire TIMEBOOST_net_22106;
wire g58291_sb;
wire TIMEBOOST_net_14380;
wire g58292_db;
wire g58292_sb;
wire TIMEBOOST_net_17520;
wire g58293_sb;
wire TIMEBOOST_net_22159;
wire g58294_sb;
wire TIMEBOOST_net_15473;
wire g58295_db;
wire g58295_sb;
wire TIMEBOOST_net_13460;
wire g58296_sb;
wire g58297_sb;
wire g58298_sb;
wire TIMEBOOST_net_13881;
wire g58299_sb;
wire TIMEBOOST_net_13028;
wire TIMEBOOST_net_20144;
wire g58300_sb;
wire TIMEBOOST_net_12695;
wire TIMEBOOST_net_22054;
wire g58301_sb;
wire TIMEBOOST_net_23465;
wire g58302_sb;
wire TIMEBOOST_net_15865;
wire g58303_sb;
wire TIMEBOOST_net_17443;
wire g58304_sb;
wire TIMEBOOST_net_12771;
wire g58305_sb;
wire g58306_db;
wire g58306_sb;
wire TIMEBOOST_net_13862;
wire g58307_sb;
wire TIMEBOOST_net_17383;
wire g58308_sb;
wire g58309_da;
wire g58309_sb;
wire TIMEBOOST_net_13863;
wire TIMEBOOST_net_21938;
wire g58310_sb;
wire TIMEBOOST_net_23519;
wire TIMEBOOST_net_12770;
wire g58311_sb;
wire TIMEBOOST_net_12621;
wire g58312_db;
wire g58312_sb;
wire TIMEBOOST_net_13856;
wire g58313_db;
wire g58313_sb;
wire TIMEBOOST_net_13867;
wire g58314_db;
wire g58314_sb;
wire TIMEBOOST_net_17384;
wire TIMEBOOST_net_13606;
wire g58315_sb;
wire TIMEBOOST_net_12623;
wire TIMEBOOST_net_7714;
wire g58316_sb;
wire TIMEBOOST_net_17385;
wire g52463_da;
wire g58317_sb;
wire g58318_db;
wire g58318_sb;
wire g65888_db;
wire g58319_db;
wire g58319_sb;
wire g58320_db;
wire g58320_sb;
wire TIMEBOOST_net_13613;
wire g58321_sb;
wire TIMEBOOST_net_13993;
wire TIMEBOOST_net_14862;
wire g58322_sb;
wire TIMEBOOST_net_8223;
wire TIMEBOOST_net_21930;
wire g58323_sb;
wire TIMEBOOST_net_12626;
wire TIMEBOOST_net_12769;
wire g58324_sb;
wire TIMEBOOST_net_12627;
wire TIMEBOOST_net_15866;
wire g58325_sb;
wire g58326_da;
wire TIMEBOOST_net_13612;
wire g58326_sb;
wire TIMEBOOST_net_12628;
wire g58327_sb;
wire TIMEBOOST_net_21168;
wire g58328_sb;
wire TIMEBOOST_net_17386;
wire g58329_db;
wire g58329_sb;
wire TIMEBOOST_net_16464;
wire g58330_db;
wire g58330_sb;
wire TIMEBOOST_net_22502;
wire g58331_db;
wire g58331_sb;
wire TIMEBOOST_net_22500;
wire TIMEBOOST_net_17250;
wire g58332_sb;
wire g58333_da;
wire g58333_sb;
wire TIMEBOOST_net_12631;
wire TIMEBOOST_net_13618;
wire g58334_sb;
wire TIMEBOOST_net_22532;
wire g58335_db;
wire g58335_sb;
wire g58336_db;
wire g58336_sb;
wire TIMEBOOST_net_13956;
wire TIMEBOOST_net_15867;
wire g58337_sb;
wire TIMEBOOST_net_21544;
wire TIMEBOOST_net_17251;
wire g58338_sb;
wire TIMEBOOST_net_13972;
wire g58339_db;
wire g58339_sb;
wire TIMEBOOST_net_13948;
wire g58340_db;
wire g58340_sb;
wire TIMEBOOST_net_14229;
wire TIMEBOOST_net_23429;
wire g58341_sb;
wire g58342_sb;
wire TIMEBOOST_net_13614;
wire g58343_sb;
wire TIMEBOOST_net_23125;
wire TIMEBOOST_net_20789;
wire g58344_sb;
wire TIMEBOOST_net_12767;
wire g58345_sb;
wire g58346_db;
wire g58346_sb;
wire g58347_sb;
wire g58348_db;
wire g58348_sb;
wire TIMEBOOST_net_14670;
wire g58349_db;
wire g58349_sb;
wire TIMEBOOST_net_12760;
wire g58350_sb;
wire TIMEBOOST_net_9325;
wire TIMEBOOST_net_21787;
wire g58351_sb;
wire TIMEBOOST_net_12766;
wire g58352_sb;
wire TIMEBOOST_net_13559;
wire TIMEBOOST_net_17445;
wire g58353_sb;
wire g58354_db;
wire g58354_sb;
wire TIMEBOOST_net_14768;
wire TIMEBOOST_net_21356;
wire g58355_sb;
wire TIMEBOOST_net_13686;
wire g58356_db;
wire g58356_sb;
wire TIMEBOOST_net_20747;
wire g58357_sb;
wire TIMEBOOST_net_8262;
wire g58358_sb;
wire n_3506;
wire TIMEBOOST_net_21775;
wire g58359_sb;
wire TIMEBOOST_net_14761;
wire g58360_sb;
wire TIMEBOOST_net_12617;
wire g58361_sb;
wire TIMEBOOST_net_20664;
wire TIMEBOOST_net_17447;
wire g58362_sb;
wire TIMEBOOST_net_21623;
wire g58363_sb;
wire TIMEBOOST_net_12228;
wire g58364_sb;
wire g58365_sb;
wire TIMEBOOST_net_13635;
wire g58366_sb;
wire g58367_da;
wire g58368_sb;
wire TIMEBOOST_net_13462;
wire g58369_db;
wire g58369_sb;
wire TIMEBOOST_net_21616;
wire g58370_db;
wire g58370_sb;
wire TIMEBOOST_net_16434;
wire g58371_db;
wire g58371_sb;
wire TIMEBOOST_net_16435;
wire g58372_sb;
wire TIMEBOOST_net_22932;
wire TIMEBOOST_net_23472;
wire g58373_sb;
wire TIMEBOOST_net_16429;
wire g58374_db;
wire g58374_sb;
wire TIMEBOOST_net_21512;
wire g58375_db;
wire g58375_sb;
wire TIMEBOOST_net_7706;
wire g58376_sb;
wire g58377_sb;
wire TIMEBOOST_net_13947;
wire g58378_sb;
wire TIMEBOOST_net_15162;
wire TIMEBOOST_net_22160;
wire g58379_sb;
wire g58380_db;
wire g58380_sb;
wire TIMEBOOST_net_15114;
wire TIMEBOOST_net_20933;
wire g58381_sb;
wire TIMEBOOST_net_13946;
wire g58382_sb;
wire TIMEBOOST_net_16659;
wire g58383_sb;
wire TIMEBOOST_net_17389;
wire TIMEBOOST_net_22300;
wire g58384_sb;
wire TIMEBOOST_net_12639;
wire TIMEBOOST_net_10587;
wire g58385_sb;
wire TIMEBOOST_net_22589;
wire g58386_sb;
wire TIMEBOOST_net_21539;
wire g58387_db;
wire g58387_sb;
wire TIMEBOOST_net_21159;
wire g58388_db;
wire g58388_sb;
wire TIMEBOOST_net_13949;
wire g58389_db;
wire g58389_sb;
wire TIMEBOOST_net_21839;
wire g58390_sb;
wire TIMEBOOST_net_22698;
wire g58391_db;
wire g58391_sb;
wire TIMEBOOST_net_13950;
wire TIMEBOOST_net_21918;
wire g58392_sb;
wire TIMEBOOST_net_20361;
wire TIMEBOOST_net_21594;
wire g58393_sb;
wire TIMEBOOST_net_15184;
wire g58394_db;
wire g58394_sb;
wire g58395_db;
wire g58395_sb;
wire TIMEBOOST_net_13984;
wire TIMEBOOST_net_21916;
wire g58396_sb;
wire g58397_db;
wire g58397_sb;
wire TIMEBOOST_net_13930;
wire TIMEBOOST_net_21925;
wire g58398_sb;
wire TIMEBOOST_net_13227;
wire g58399_db;
wire g58399_sb;
wire g58400_db;
wire g58400_sb;
wire TIMEBOOST_net_14558;
wire g58401_sb;
wire TIMEBOOST_net_13877;
wire g58402_sb;
wire TIMEBOOST_net_13568;
wire g58403_sb;
wire TIMEBOOST_net_13961;
wire g58404_db;
wire g58404_sb;
wire g58405_db;
wire g58405_sb;
wire TIMEBOOST_net_23482;
wire TIMEBOOST_net_21581;
wire g58406_sb;
wire TIMEBOOST_net_15179;
wire g58407_db;
wire g58407_sb;
wire TIMEBOOST_net_14813;
wire TIMEBOOST_net_12386;
wire g58408_sb;
wire TIMEBOOST_net_12647;
wire TIMEBOOST_net_12385;
wire g58409_sb;
wire TIMEBOOST_net_13575;
wire g58410_db;
wire g58410_sb;
wire TIMEBOOST_net_13584;
wire g58411_db;
wire g58411_sb;
wire TIMEBOOST_net_13712;
wire g58412_db;
wire g58412_sb;
wire TIMEBOOST_net_13588;
wire g58413_db;
wire g58413_sb;
wire TIMEBOOST_net_16451;
wire TIMEBOOST_net_22262;
wire g58414_sb;
wire g58415_db;
wire g58415_sb;
wire TIMEBOOST_net_13709;
wire g58416_db;
wire g58416_sb;
wire TIMEBOOST_net_13374;
wire g58417_sb;
wire TIMEBOOST_net_8835;
wire g58418_sb;
wire g65375_db;
wire g58419_sb;
wire TIMEBOOST_net_21920;
wire TIMEBOOST_net_7700;
wire g58420_sb;
wire g58421_da;
wire TIMEBOOST_net_14536;
wire g58421_sb;
wire TIMEBOOST_net_14248;
wire TIMEBOOST_net_12616;
wire g58422_sb;
wire TIMEBOOST_net_17390;
wire g58423_db;
wire g58423_sb;
wire TIMEBOOST_net_8309;
wire TIMEBOOST_net_12615;
wire g58424_sb;
wire TIMEBOOST_net_8837;
wire g58425_db;
wire g58425_sb;
wire TIMEBOOST_net_17391;
wire g58426_sb;
wire TIMEBOOST_net_12927;
wire TIMEBOOST_net_13634;
wire g58427_sb;
wire g58428_db;
wire g58428_sb;
wire TIMEBOOST_net_8840;
wire TIMEBOOST_net_21915;
wire g58429_sb;
wire TIMEBOOST_net_13885;
wire g58430_db;
wire g58430_sb;
wire TIMEBOOST_net_21907;
wire g58431_sb;
wire g58432_sb;
wire g58433_sb;
wire g58434_da;
wire TIMEBOOST_net_7697;
wire g58434_sb;
wire g58435_sb;
wire g58436_sb;
wire TIMEBOOST_net_8250;
wire g58437_sb;
wire g58438_db;
wire g58438_sb;
wire TIMEBOOST_net_21266;
wire g58439_db;
wire g58439_sb;
wire TIMEBOOST_net_13870;
wire g58440_sb;
wire TIMEBOOST_net_13633;
wire g58441_sb;
wire TIMEBOOST_net_21600;
wire TIMEBOOST_net_23389;
wire g58442_sb;
wire TIMEBOOST_net_20402;
wire g58443_sb;
wire TIMEBOOST_net_13487;
wire TIMEBOOST_net_17273;
wire g58444_sb;
wire g58445_sb;
wire TIMEBOOST_net_7424;
wire g58446_db;
wire g58446_sb;
wire g58447_db;
wire g58447_sb;
wire TIMEBOOST_net_22554;
wire g58448_db;
wire g58448_sb;
wire TIMEBOOST_net_22663;
wire g58449_sb;
wire g58450_sb;
wire g58451_sb;
wire TIMEBOOST_net_14901;
wire g58452_db;
wire g58452_sb;
wire TIMEBOOST_net_23360;
wire TIMEBOOST_net_21957;
wire g58453_sb;
wire g58454_sb;
wire TIMEBOOST_net_17217;
wire TIMEBOOST_net_20227;
wire g58455_sb;
wire TIMEBOOST_net_22664;
wire g58456_sb;
wire TIMEBOOST_net_22595;
wire n_16565;
wire g58457_sb;
wire TIMEBOOST_net_10343;
wire TIMEBOOST_net_10708;
wire g58458_sb;
wire FE_RN_302_0;
wire g58459_sb;
wire TIMEBOOST_net_21465;
wire g58460_sb;
wire TIMEBOOST_net_17064;
wire TIMEBOOST_net_10703;
wire g58461_sb;
wire TIMEBOOST_net_14121;
wire TIMEBOOST_net_20790;
wire g58462_sb;
wire TIMEBOOST_net_10405;
wire g58463_sb;
wire g58464_sb;
wire TIMEBOOST_net_14682;
wire g58465_sb;
wire g58466_sb;
wire TIMEBOOST_net_10339;
wire g58467_sb;
wire TIMEBOOST_net_20186;
wire g58468_sb;
wire TIMEBOOST_net_17100;
wire g58469_sb;
wire TIMEBOOST_net_10338;
wire TIMEBOOST_net_10702;
wire g58470_sb;
wire TIMEBOOST_net_20195;
wire g58471_sb;
wire g58472_sb;
wire TIMEBOOST_net_10337;
wire TIMEBOOST_net_17468;
wire g58473_sb;
wire TIMEBOOST_net_10336;
wire g58474_sb;
wire TIMEBOOST_net_10335;
wire g58475_sb;
wire TIMEBOOST_net_20367;
wire g58476_sb;
wire TIMEBOOST_net_10333;
wire g58477_sb;
wire TIMEBOOST_net_14290;
wire TIMEBOOST_net_10684;
wire g58478_sb;
wire TIMEBOOST_net_17099;
wire TIMEBOOST_net_15049;
wire g58479_sb;
wire TIMEBOOST_net_10401;
wire g58480_sb;
wire TIMEBOOST_net_10332;
wire g58481_sb;
wire TIMEBOOST_net_15046;
wire g58482_sb;
wire TIMEBOOST_net_17098;
wire TIMEBOOST_net_17466;
wire g58483_sb;
wire TIMEBOOST_net_17467;
wire g58484_sb;
wire TIMEBOOST_net_10398;
wire TIMEBOOST_net_12440;
wire g58485_sb;
wire TIMEBOOST_net_10397;
wire g58486_sb;
wire TIMEBOOST_net_13543;
wire g58487_sb;
wire TIMEBOOST_net_17394;
wire TIMEBOOST_net_13628;
wire g58488_sb;
wire TIMEBOOST_net_17101;
wire TIMEBOOST_net_10712;
wire g58489_sb;
wire g58490_p;
wire g58569_p;
wire TIMEBOOST_net_11473;
wire TIMEBOOST_net_16312;
wire g58574_sb;
wire TIMEBOOST_net_11474;
wire TIMEBOOST_net_17199;
wire g58576_sb;
wire g58582_p;
wire TIMEBOOST_net_16147;
wire TIMEBOOST_net_16735;
wire g58586_sb;
wire g58587_sb;
wire TIMEBOOST_net_12445;
wire g58588_sb;
wire TIMEBOOST_net_11475;
wire TIMEBOOST_net_16255;
wire g58589_sb;
wire TIMEBOOST_net_11476;
wire g58590_sb;
wire TIMEBOOST_net_23240;
wire g58591_sb;
wire TIMEBOOST_net_16736;
wire g58592_sb;
wire TIMEBOOST_net_15183;
wire g58593_sb;
wire TIMEBOOST_net_16737;
wire g58594_sb;
wire TIMEBOOST_net_15341;
wire TIMEBOOST_net_17403;
wire g58595_sb;
wire TIMEBOOST_net_15446;
wire TIMEBOOST_net_23411;
wire g58596_sb;
wire g58597_sb;
wire TIMEBOOST_net_22130;
wire g58598_sb;
wire g58599_p;
wire TIMEBOOST_net_16542;
wire g58600_sb;
wire TIMEBOOST_net_16543;
wire g58601_sb;
wire TIMEBOOST_net_21223;
wire TIMEBOOST_net_21662;
wire g58605_sb;
wire TIMEBOOST_net_22373;
wire g58606_sb;
wire TIMEBOOST_net_16150;
wire TIMEBOOST_net_16738;
wire g58607_sb;
wire TIMEBOOST_net_16313;
wire g58608_sb;
wire TIMEBOOST_net_12360;
wire TIMEBOOST_net_9860;
wire g58609_sb;
wire g58610_sb;
wire TIMEBOOST_net_20182;
wire g58611_sb;
wire TIMEBOOST_net_16314;
wire g58616_sb;
wire g58617_sb;
wire TIMEBOOST_net_16316;
wire g58618_sb;
wire TIMEBOOST_net_6735;
wire TIMEBOOST_net_16317;
wire g58619_sb;
wire TIMEBOOST_net_6736;
wire g58620_sb;
wire g58621_sb;
wire TIMEBOOST_net_11301;
wire g58622_sb;
wire TIMEBOOST_net_11302;
wire g58630_sb;
wire g58631_sb;
wire TIMEBOOST_net_23160;
wire g58632_sb;
wire g58633_sb;
wire TIMEBOOST_net_23538;
wire g58634_sb;
wire g58635_sb;
wire TIMEBOOST_net_16985;
wire g58636_sb;
wire TIMEBOOST_net_16544;
wire g58640_sb;
wire TIMEBOOST_net_16545;
wire TIMEBOOST_net_15471;
wire g58652_sb;
wire TIMEBOOST_net_16546;
wire TIMEBOOST_net_6908;
wire g58653_sb;
wire TIMEBOOST_net_16547;
wire g58654_sb;
wire g58655_sb;
wire g58656_p;
wire g58692_p;
wire g58695_p;
wire g58742_p;
wire g58744_p;
wire g58759_p;
wire g58760_p;
wire g58761_p;
wire g58763_p;
wire g58764_p;
wire TIMEBOOST_net_21628;
wire TIMEBOOST_net_21645;
wire g58767_sb;
wire TIMEBOOST_net_21464;
wire g58768_sb;
wire g58769_sb;
wire g58770_sb;
wire g58771_sb;
wire TIMEBOOST_net_13668;
wire g58772_sb;
wire TIMEBOOST_net_16653;
wire TIMEBOOST_net_13557;
wire g58773_sb;
wire TIMEBOOST_net_14542;
wire g58774_sb;
wire TIMEBOOST_net_22414;
wire g58775_sb;
wire TIMEBOOST_net_9326;
wire TIMEBOOST_net_17458;
wire g58776_sb;
wire TIMEBOOST_net_9354;
wire TIMEBOOST_net_114;
wire g58777_sb;
wire TIMEBOOST_net_9355;
wire TIMEBOOST_net_14144;
wire g58778_sb;
wire TIMEBOOST_net_20514;
wire g58779_sb;
wire TIMEBOOST_net_21;
wire TIMEBOOST_net_20623;
wire TIMEBOOST_net_9356;
wire TIMEBOOST_net_116;
wire g58782_sb;
wire TIMEBOOST_net_22;
wire g58783_sb;
wire TIMEBOOST_net_23;
wire TIMEBOOST_net_71;
wire g58785_sb;
wire g58786_sb;
wire TIMEBOOST_net_22161;
wire TIMEBOOST_net_117;
wire g58787_sb;
wire TIMEBOOST_net_22110;
wire g58788_sb;
wire TIMEBOOST_net_9793;
wire TIMEBOOST_net_22343;
wire g58789_sb;
wire TIMEBOOST_net_13552;
wire g58790_sb;
wire TIMEBOOST_net_13553;
wire g58791_sb;
wire TIMEBOOST_net_9357;
wire TIMEBOOST_net_118;
wire g58792_sb;
wire TIMEBOOST_net_37;
wire TIMEBOOST_net_13122;
wire g58793_sb;
wire TIMEBOOST_net_13368;
wire g58794_sb;
wire TIMEBOOST_net_16043;
wire g58795_sb;
wire TIMEBOOST_net_15539;
wire TIMEBOOST_net_17451;
wire TIMEBOOST_net_22287;
wire g58797_sb;
wire TIMEBOOST_net_16041;
wire g58798_db;
wire g58798_sb;
wire TIMEBOOST_net_23558;
wire TIMEBOOST_net_5468;
wire g58799_sb;
wire TIMEBOOST_net_5469;
wire g58800_sb;
wire TIMEBOOST_net_6914;
wire TIMEBOOST_net_22142;
wire g58801_sb;
wire TIMEBOOST_net_6915;
wire g58802_sb;
wire TIMEBOOST_net_17050;
wire TIMEBOOST_net_13719;
wire g58803_sb;
wire g58804_sb;
wire TIMEBOOST_net_21688;
wire TIMEBOOST_net_13720;
wire g58805_sb;
wire TIMEBOOST_net_10603;
wire g58806_sb;
wire TIMEBOOST_net_16708;
wire g58807_sb;
wire TIMEBOOST_net_16447;
wire TIMEBOOST_net_21369;
wire g58808_sb;
wire TIMEBOOST_net_21671;
wire g58809_sb;
wire g58810_sb;
wire TIMEBOOST_net_16982;
wire TIMEBOOST_net_17327;
wire g58811_sb;
wire g58812_sb;
wire TIMEBOOST_net_16471;
wire g58813_sb;
wire TIMEBOOST_net_12550;
wire g58814_sb;
wire TIMEBOOST_net_21768;
wire g58815_sb;
wire g58816_sb;
wire TIMEBOOST_net_20538;
wire TIMEBOOST_net_14449;
wire g58817_sb;
wire g58818_sb;
wire g58819_sb;
wire g58820_sb;
wire g58821_sb;
wire TIMEBOOST_net_23194;
wire TIMEBOOST_net_16714;
wire g58822_sb;
wire TIMEBOOST_net_21711;
wire TIMEBOOST_net_14674;
wire g58823_sb;
wire TIMEBOOST_net_16715;
wire g58824_sb;
wire TIMEBOOST_net_12542;
wire TIMEBOOST_net_16709;
wire g58825_sb;
wire TIMEBOOST_net_16710;
wire g58826_sb;
wire TIMEBOOST_net_21833;
wire g58827_sb;
wire TIMEBOOST_net_16716;
wire g58828_sb;
wire TIMEBOOST_net_21315;
wire TIMEBOOST_net_16711;
wire g58829_sb;
wire TIMEBOOST_net_16712;
wire g58830_sb;
wire TIMEBOOST_net_14672;
wire g58831_sb;
wire TIMEBOOST_net_16056;
wire g58832_sb;
wire g58833_sb;
wire g58834_sb;
wire g58835_sb;
wire TIMEBOOST_net_12504;
wire TIMEBOOST_net_16057;
wire g58836_sb;
wire TIMEBOOST_net_17097;
wire TIMEBOOST_net_17469;
wire g58837_sb;
wire TIMEBOOST_net_22634;
wire TIMEBOOST_net_10696;
wire g58838_sb;
wire TIMEBOOST_net_17096;
wire g58839_sb;
wire TIMEBOOST_net_17095;
wire g58840_sb;
wire TIMEBOOST_net_10393;
wire g58841_sb;
wire TIMEBOOST_net_16548;
wire TIMEBOOST_net_20204;
wire g58842_sb;
wire TIMEBOOST_net_17023;
wire g58843_sb;
wire TIMEBOOST_net_9329;
wire g59082_sb;
wire g59086_p;
wire TIMEBOOST_net_21519;
wire g59089_sb;
wire TIMEBOOST_net_10870;
wire g59090_sb;
wire TIMEBOOST_net_17006;
wire TIMEBOOST_net_13521;
wire g59092_sb;
wire TIMEBOOST_net_16697;
wire TIMEBOOST_net_21480;
wire g59093_sb;
wire g59095_p;
wire TIMEBOOST_net_9476;
wire TIMEBOOST_net_10111;
wire g59096_sb;
wire g61987_db;
wire TIMEBOOST_net_16694;
wire g59097_sb;
wire TIMEBOOST_net_10180;
wire g59098_sb;
wire TIMEBOOST_net_13899;
wire TIMEBOOST_net_10873;
wire g59109_sb;
wire TIMEBOOST_net_10177;
wire TIMEBOOST_net_10874;
wire g59110_sb;
wire TIMEBOOST_net_10875;
wire g59111_sb;
wire TIMEBOOST_net_10174;
wire TIMEBOOST_net_10876;
wire g59112_sb;
wire TIMEBOOST_net_10173;
wire g59113_sb;
wire TIMEBOOST_net_16984;
wire TIMEBOOST_net_10171;
wire TIMEBOOST_net_14963;
wire TIMEBOOST_net_10168;
wire TIMEBOOST_net_21437;
wire TIMEBOOST_net_10166;
wire g59118_sb;
wire TIMEBOOST_net_10163;
wire TIMEBOOST_net_10882;
wire TIMEBOOST_net_16327;
wire TIMEBOOST_net_14924;
wire TIMEBOOST_net_21656;
wire g59121_sb;
wire TIMEBOOST_net_11524;
wire g59122_sb;
wire TIMEBOOST_net_17524;
wire TIMEBOOST_net_5475;
wire g59123_sb;
wire g59124_p;
wire g59125_p;
wire TIMEBOOST_net_16752;
wire g59126_db;
wire g59126_sb;
wire g59127_p;
wire g59128_p;
wire g59196_p;
wire g59198_p;
wire g59199_p;
wire g59201_p;
wire g59206_p;
wire g59226_da;
wire g59226_sb;
wire g59227_p;
wire g59228_p;
wire g59229_p;
wire TIMEBOOST_net_22308;
wire TIMEBOOST_net_21474;
wire g59230_sb;
wire TIMEBOOST_net_5470;
wire g59231_sb;
wire g59232_BP;
wire g59232_p;
wire TIMEBOOST_net_21287;
wire TIMEBOOST_net_13968;
wire g59234_sb;
wire g59239_sb;
wire g59240_sb;
wire g59296_p;
wire g59300_p;
wire g59331_p;
wire g59344_p;
wire g59345_p;
wire g59346_p;
wire g59347_p;
wire TIMEBOOST_net_10461;
wire g59350_sb;
wire g59364_p;
wire g59367_p;
wire TIMEBOOST_net_778;
wire g59368_sb;
wire TIMEBOOST_net_12764;
wire TIMEBOOST_net_779;
wire g59369_sb;
wire TIMEBOOST_net_21222;
wire g59370_sb;
wire TIMEBOOST_net_13620;
wire g59371_sb;
wire TIMEBOOST_net_21542;
wire g59372_sb;
wire TIMEBOOST_net_13623;
wire g59373_sb;
wire g59374_p;
wire g59377_p;
wire TIMEBOOST_net_7423;
wire g59378_sb;
wire TIMEBOOST_net_13622;
wire g59379_sb;
wire TIMEBOOST_net_13680;
wire TIMEBOOST_net_10709;
wire g59380_sb;
wire TIMEBOOST_net_13679;
wire g59381_sb;
wire TIMEBOOST_net_21301;
wire TIMEBOOST_net_10053;
wire g59382_sb;
wire TIMEBOOST_net_20729;
wire TIMEBOOST_net_21803;
wire g59383_sb;
wire TIMEBOOST_net_21672;
wire g59384_sb;
wire g59385_p;
wire g59386_p;
wire TIMEBOOST_net_13682;
wire TIMEBOOST_net_10267;
wire g59387_sb;
wire g59388_p;
wire g59389_p;
wire g59622_p;
wire g59623_p;
wire g59627_p;
wire g59659_p;
wire g59665_p;
wire g59666_p;
wire g59670_p;
wire g59674_p;
wire g59721_p;
wire g59761_p;
wire TIMEBOOST_net_20257;
wire g59763_sb;
wire TIMEBOOST_net_9358;
wire TIMEBOOST_net_20579;
wire TIMEBOOST_net_16745;
wire g59783_p;
wire g59785_p;
wire g59790_p;
wire g59791_p;
wire g59793_p;
wire g59794_p;
wire g59795_p;
wire TIMEBOOST_net_16693;
wire g59796_db;
wire g59796_sb;
wire TIMEBOOST_net_13378;
wire TIMEBOOST_net_21517;
wire g59797_sb;
wire TIMEBOOST_net_9477;
wire TIMEBOOST_net_10101;
wire g59798_sb;
wire TIMEBOOST_net_9404;
wire TIMEBOOST_net_13547;
wire g59799_sb;
wire g59800_db;
wire g59800_sb;
wire TIMEBOOST_net_15312;
wire g59801_sb;
wire g59802_p;
wire g59803_p;
wire TIMEBOOST_net_11410;
wire g61985_db;
wire g59804_sb;
wire TIMEBOOST_net_16623;
wire g59805_sb;
wire TIMEBOOST_net_13690;
wire g59806_sb;
wire TIMEBOOST_net_21344;
wire g61981_db;
wire g59807_sb;
wire g61980_db;
wire g59808_sb;
wire TIMEBOOST_net_13579;
wire g59809_sb;
wire g60298_p;
wire g60304_p;
wire g60307_p;
wire g60310_p;
wire g60319_p;
wire g60321_p;
wire g60330_p;
wire g60339_p;
wire g60345_p;
wire TIMEBOOST_net_331;
wire g60407_sb;
wire TIMEBOOST_net_14744;
wire TIMEBOOST_net_9322;
wire TIMEBOOST_net_14513;
wire TIMEBOOST_net_22489;
wire g60409_sb;
wire g60414_p;
wire g60415_p;
wire g60557_p;
wire g60591_p;
wire g60603_da;
wire g60603_sb;
wire TIMEBOOST_net_10905;
wire TIMEBOOST_net_9479;
wire g60604_sb;
wire TIMEBOOST_net_5550;
wire TIMEBOOST_net_11420;
wire g60605_sb;
wire TIMEBOOST_net_10705;
wire TIMEBOOST_net_21346;
wire g60606_sb;
wire TIMEBOOST_net_23532;
wire g60607_sb;
wire g60608_sb;
wire TIMEBOOST_net_11389;
wire g60609_sb;
wire TIMEBOOST_net_16953;
wire TIMEBOOST_net_23390;
wire g60610_sb;
wire g58406_db;
wire g60611_sb;
wire TIMEBOOST_net_11175;
wire TIMEBOOST_net_11392;
wire g60612_sb;
wire g60613_sb;
wire TIMEBOOST_net_21254;
wire g60614_sb;
wire TIMEBOOST_net_10906;
wire TIMEBOOST_net_21294;
wire g60615_sb;
wire TIMEBOOST_net_5560;
wire g60616_sb;
wire TIMEBOOST_net_21381;
wire g60617_sb;
wire TIMEBOOST_net_11353;
wire TIMEBOOST_net_21394;
wire g60618_sb;
wire TIMEBOOST_net_11352;
wire g60619_sb;
wire TIMEBOOST_net_23511;
wire TIMEBOOST_net_11399;
wire g60620_sb;
wire TIMEBOOST_net_23525;
wire TIMEBOOST_net_11400;
wire g60621_sb;
wire TIMEBOOST_net_21390;
wire g60622_sb;
wire TIMEBOOST_net_21357;
wire g60623_sb;
wire TIMEBOOST_net_23517;
wire g60624_sb;
wire TIMEBOOST_net_15367;
wire TIMEBOOST_net_23455;
wire g60625_sb;
wire g60626_sb;
wire TIMEBOOST_net_11340;
wire TIMEBOOST_net_21396;
wire g60627_sb;
wire g60628_sb;
wire TIMEBOOST_net_15370;
wire g60629_sb;
wire TIMEBOOST_net_5572;
wire TIMEBOOST_net_21471;
wire g60630_sb;
wire TIMEBOOST_net_11637;
wire g60631_sb;
wire TIMEBOOST_net_21573;
wire TIMEBOOST_net_11362;
wire g60632_sb;
wire TIMEBOOST_net_21361;
wire g60633_sb;
wire n_3623;
wire g60634_sb;
wire TIMEBOOST_net_11526;
wire TIMEBOOST_net_23542;
wire g60635_sb;
wire TIMEBOOST_net_10907;
wire g60636_sb;
wire TIMEBOOST_net_21398;
wire g60637_sb;
wire TIMEBOOST_net_12970;
wire TIMEBOOST_net_15069;
wire g60638_sb;
wire g60639_sb;
wire TIMEBOOST_net_11444;
wire TIMEBOOST_net_16780;
wire g60640_sb;
wire TIMEBOOST_net_23515;
wire TIMEBOOST_net_21380;
wire g60641_sb;
wire TIMEBOOST_net_11443;
wire TIMEBOOST_net_21372;
wire g60642_sb;
wire TIMEBOOST_net_17052;
wire g60643_sb;
wire TIMEBOOST_net_11577;
wire TIMEBOOST_net_11201;
wire g60644_sb;
wire g75178_da;
wire g60645_sb;
wire TIMEBOOST_net_12630;
wire TIMEBOOST_net_15056;
wire g60646_sb;
wire g59382_db;
wire TIMEBOOST_net_16777;
wire g60647_sb;
wire TIMEBOOST_net_16776;
wire g60648_sb;
wire TIMEBOOST_net_21689;
wire g60649_sb;
wire g60650_sb;
wire TIMEBOOST_net_10908;
wire g60651_sb;
wire TIMEBOOST_net_23549;
wire g60652_sb;
wire TIMEBOOST_net_21240;
wire g60653_sb;
wire TIMEBOOST_net_5592;
wire g60654_sb;
wire g60655_sb;
wire TIMEBOOST_net_21242;
wire g60656_sb;
wire TIMEBOOST_net_5595;
wire TIMEBOOST_net_21243;
wire g60657_sb;
wire g60658_sb;
wire TIMEBOOST_net_11467;
wire TIMEBOOST_net_15057;
wire g60659_sb;
wire TIMEBOOST_net_21300;
wire TIMEBOOST_net_15058;
wire g60660_sb;
wire TIMEBOOST_net_15059;
wire g60661_sb;
wire TIMEBOOST_net_11482;
wire TIMEBOOST_net_15060;
wire g60662_sb;
wire TIMEBOOST_net_21489;
wire TIMEBOOST_net_15061;
wire g60663_sb;
wire TIMEBOOST_net_10909;
wire g60664_sb;
wire TIMEBOOST_net_11623;
wire g60665_sb;
wire TIMEBOOST_net_21545;
wire TIMEBOOST_net_11339;
wire g60666_sb;
wire TIMEBOOST_net_21174;
wire g60667_sb;
wire TIMEBOOST_net_23400;
wire TIMEBOOST_net_15980;
wire g60668_sb;
wire g60669_sb;
wire TIMEBOOST_net_10910;
wire TIMEBOOST_net_9472;
wire g60670_sb;
wire g60671_sb;
wire TIMEBOOST_net_11525;
wire g60672_sb;
wire TIMEBOOST_net_10911;
wire g60673_sb;
wire g60674_sb;
wire TIMEBOOST_net_20723;
wire g60675_sb;
wire g60676_sb;
wire TIMEBOOST_net_16647;
wire TIMEBOOST_net_15314;
wire g60677_sb;
wire TIMEBOOST_net_13973;
wire g60678_sb;
wire TIMEBOOST_net_22728;
wire TIMEBOOST_net_5472;
wire g60679_sb;
wire TIMEBOOST_net_12961;
wire g60681_db;
wire g60681_sb;
wire TIMEBOOST_net_10185;
wire g60682_sb;
wire g60686_sb;
wire TIMEBOOST_net_22507;
wire TIMEBOOST_net_22024;
wire g60687_sb;
wire TIMEBOOST_net_152;
wire TIMEBOOST_net_16174;
wire g60688_sb;
wire TIMEBOOST_net_20260;
wire g60689_sb;
wire TIMEBOOST_net_23201;
wire g60690_sb;
wire TIMEBOOST_net_16997;
wire g60691_sb;
wire TIMEBOOST_net_15531;
wire g60692_sb;
wire g60693_p;
wire g60694_p;
wire g60695_p;
wire g60696_p;
wire TIMEBOOST_net_91;
wire TIMEBOOST_net_21621;
wire g61569_p;
wire g61570_p;
wire g61572_p;
wire g61575_p;
wire g61581_p;
wire g61582_p;
wire g61597_p;
wire g61606_p;
wire g61617_p;
wire TIMEBOOST_net_15220;
wire TIMEBOOST_net_9500;
wire g61618_p;
wire g61622_p;
wire g61636_p;
wire g61637_p;
wire g61654_p;
wire g61676_sb;
wire g61689_p;
wire g61693_p;
wire TIMEBOOST_net_14983;
wire g61697_sb;
wire TIMEBOOST_net_23493;
wire g61698_db;
wire g61698_sb;
wire TIMEBOOST_net_22732;
wire TIMEBOOST_net_585;
wire g61699_sb;
wire TIMEBOOST_net_15065;
wire TIMEBOOST_net_343;
wire g61700_sb;
wire TIMEBOOST_net_21501;
wire g61701_sb;
wire TIMEBOOST_net_23332;
wire g61702_db;
wire g61702_sb;
wire TIMEBOOST_net_269;
wire g61703_db;
wire g61703_sb;
wire TIMEBOOST_net_15067;
wire g61704_sb;
wire TIMEBOOST_net_9366;
wire g61705_db;
wire g61705_sb;
wire TIMEBOOST_net_15064;
wire TIMEBOOST_net_345;
wire g61706_sb;
wire TIMEBOOST_net_21195;
wire TIMEBOOST_net_9346;
wire g61707_sb;
wire TIMEBOOST_net_271;
wire g61708_db;
wire g61708_sb;
wire g65784_db;
wire g61709_db;
wire g61709_sb;
wire TIMEBOOST_net_273;
wire g61710_db;
wire g61710_sb;
wire TIMEBOOST_net_22753;
wire g61711_sb;
wire g61712_sb;
wire TIMEBOOST_net_9367;
wire g61713_db;
wire g61714_sb;
wire TIMEBOOST_net_10634;
wire g61715_db;
wire g61715_sb;
wire TIMEBOOST_net_13379;
wire TIMEBOOST_net_587;
wire g61716_sb;
wire TIMEBOOST_net_275;
wire g61717_db;
wire g61717_sb;
wire TIMEBOOST_net_22351;
wire g61718_sb;
wire TIMEBOOST_net_15047;
wire g61719_sb;
wire TIMEBOOST_net_15048;
wire TIMEBOOST_net_350;
wire g61720_sb;
wire TIMEBOOST_net_13439;
wire g61721_sb;
wire g61722_sb;
wire TIMEBOOST_net_14680;
wire g61723_sb;
wire TIMEBOOST_net_21161;
wire g61724_sb;
wire TIMEBOOST_net_109;
wire g61725_sb;
wire TIMEBOOST_net_276;
wire g61726_db;
wire g61726_sb;
wire TIMEBOOST_net_21176;
wire g61727_sb;
wire TIMEBOOST_net_16769;
wire TIMEBOOST_net_13510;
wire g61728_sb;
wire TIMEBOOST_net_15013;
wire g61729_sb;
wire TIMEBOOST_net_20264;
wire g61730_sb;
wire TIMEBOOST_net_21179;
wire TIMEBOOST_net_13509;
wire g61731_sb;
wire TIMEBOOST_net_319;
wire g61732_db;
wire g61732_sb;
wire TIMEBOOST_net_20444;
wire g61733_sb;
wire TIMEBOOST_net_321;
wire g61734_db;
wire g61734_sb;
wire TIMEBOOST_net_322;
wire g61735_db;
wire g61735_sb;
wire TIMEBOOST_net_12387;
wire g61736_db;
wire g61736_sb;
wire TIMEBOOST_net_7630;
wire TIMEBOOST_net_13915;
wire g61737_sb;
wire TIMEBOOST_net_14840;
wire TIMEBOOST_net_9347;
wire g61738_sb;
wire TIMEBOOST_net_21165;
wire TIMEBOOST_net_13508;
wire g61739_sb;
wire g61740_db;
wire g61740_sb;
wire TIMEBOOST_net_326;
wire g61741_db;
wire g61741_sb;
wire TIMEBOOST_net_327;
wire g61742_db;
wire g61742_sb;
wire TIMEBOOST_net_328;
wire g61743_db;
wire g61743_sb;
wire TIMEBOOST_net_14469;
wire g61744_sb;
wire TIMEBOOST_net_360;
wire g61745_sb;
wire TIMEBOOST_net_14908;
wire g61746_db;
wire g61746_sb;
wire TIMEBOOST_net_14903;
wire g61747_sb;
wire TIMEBOOST_net_329;
wire g61748_db;
wire g61748_sb;
wire TIMEBOOST_net_17059;
wire g61749_db;
wire g61749_sb;
wire TIMEBOOST_net_20524;
wire TIMEBOOST_net_362;
wire g61750_sb;
wire TIMEBOOST_net_14940;
wire TIMEBOOST_net_363;
wire g61751_sb;
wire TIMEBOOST_net_9348;
wire g61752_sb;
wire TIMEBOOST_net_14935;
wire TIMEBOOST_net_9259;
wire g61753_sb;
wire TIMEBOOST_net_21273;
wire TIMEBOOST_net_365;
wire g61754_sb;
wire TIMEBOOST_net_14913;
wire n_8746;
wire g61755_sb;
wire TIMEBOOST_net_23226;
wire TIMEBOOST_net_14079;
wire g61756_sb;
wire g61757_sb;
wire TIMEBOOST_net_14931;
wire TIMEBOOST_net_15726;
wire g61758_sb;
wire TIMEBOOST_net_21042;
wire TIMEBOOST_net_369;
wire g61759_sb;
wire TIMEBOOST_net_21182;
wire TIMEBOOST_net_370;
wire g61760_sb;
wire TIMEBOOST_net_21942;
wire g61761_sb;
wire TIMEBOOST_net_16490;
wire TIMEBOOST_net_16654;
wire g61762_sb;
wire TIMEBOOST_net_16354;
wire g61763_sb;
wire TIMEBOOST_net_330;
wire g61764_db;
wire g61764_sb;
wire g61765_db;
wire g61765_sb;
wire TIMEBOOST_net_15028;
wire TIMEBOOST_net_20871;
wire g61766_sb;
wire g61767_db;
wire g61767_sb;
wire TIMEBOOST_net_9349;
wire g61768_sb;
wire TIMEBOOST_net_5434;
wire g61769_sb;
wire TIMEBOOST_net_21234;
wire TIMEBOOST_net_12677;
wire g61770_sb;
wire TIMEBOOST_net_15189;
wire g61771_db;
wire g61771_sb;
wire TIMEBOOST_net_14653;
wire g61772_db;
wire g61772_sb;
wire TIMEBOOST_net_14613;
wire g61773_sb;
wire TIMEBOOST_net_376;
wire g61774_sb;
wire g61775_db;
wire g61775_sb;
wire TIMEBOOST_net_23327;
wire g61776_db;
wire TIMEBOOST_net_15192;
wire g61777_db;
wire g61777_sb;
wire TIMEBOOST_net_593;
wire g61778_sb;
wire g61779_db;
wire g61779_sb;
wire g61780_sb;
wire g61781_sb;
wire TIMEBOOST_net_20472;
wire TIMEBOOST_net_594;
wire g61782_sb;
wire g61783_db;
wire g61783_sb;
wire TIMEBOOST_net_21153;
wire TIMEBOOST_net_378;
wire g61784_sb;
wire TIMEBOOST_net_379;
wire g61785_sb;
wire TIMEBOOST_net_15014;
wire TIMEBOOST_net_380;
wire g61786_sb;
wire TIMEBOOST_net_21160;
wire g61787_sb;
wire TIMEBOOST_net_382;
wire g61788_sb;
wire TIMEBOOST_net_383;
wire g61789_sb;
wire g61790_sb;
wire TIMEBOOST_net_21219;
wire TIMEBOOST_net_21148;
wire g61791_sb;
wire TIMEBOOST_net_386;
wire g61792_sb;
wire TIMEBOOST_net_387;
wire g61793_sb;
wire TIMEBOOST_net_21010;
wire TIMEBOOST_net_388;
wire g61794_sb;
wire TIMEBOOST_net_21217;
wire TIMEBOOST_net_13674;
wire g61795_sb;
wire TIMEBOOST_net_501;
wire g61796_db;
wire g61796_sb;
wire g61797_db;
wire g61797_sb;
wire g61798_db;
wire g61798_sb;
wire TIMEBOOST_net_13675;
wire g61799_sb;
wire TIMEBOOST_net_21183;
wire TIMEBOOST_net_12277;
wire g61800_sb;
wire TIMEBOOST_net_9501;
wire g61801_db;
wire g61801_sb;
wire TIMEBOOST_net_14936;
wire TIMEBOOST_net_13287;
wire g61802_sb;
wire TIMEBOOST_net_14883;
wire TIMEBOOST_net_392;
wire g61803_sb;
wire TIMEBOOST_net_13206;
wire g61804_db;
wire g61804_sb;
wire TIMEBOOST_net_14955;
wire TIMEBOOST_net_393;
wire g61805_sb;
wire TIMEBOOST_net_13598;
wire g61806_sb;
wire TIMEBOOST_net_575;
wire TIMEBOOST_net_9350;
wire g61807_sb;
wire TIMEBOOST_net_315;
wire g61808_db;
wire g61808_sb;
wire TIMEBOOST_net_22095;
wire g61809_sb;
wire TIMEBOOST_net_576;
wire g61810_db;
wire g61810_sb;
wire TIMEBOOST_net_17490;
wire g61811_sb;
wire TIMEBOOST_net_316;
wire g61812_db;
wire g61812_sb;
wire TIMEBOOST_net_21248;
wire TIMEBOOST_net_16959;
wire g61813_sb;
wire TIMEBOOST_net_397;
wire g61814_sb;
wire g65709_db;
wire TIMEBOOST_net_9781;
wire g61815_sb;
wire TIMEBOOST_net_530;
wire g61816_db;
wire g61816_sb;
wire g61817_sb;
wire TIMEBOOST_net_577;
wire g61818_sb;
wire TIMEBOOST_net_21666;
wire g61819_sb;
wire TIMEBOOST_net_317;
wire g61820_db;
wire g61820_sb;
wire TIMEBOOST_net_15037;
wire TIMEBOOST_net_399;
wire g61821_sb;
wire g61822_sb;
wire TIMEBOOST_net_21166;
wire TIMEBOOST_net_400;
wire g61823_sb;
wire TIMEBOOST_net_14854;
wire TIMEBOOST_net_23425;
wire g61824_sb;
wire TIMEBOOST_net_20471;
wire TIMEBOOST_net_597;
wire g61825_sb;
wire TIMEBOOST_net_13135;
wire g61826_sb;
wire TIMEBOOST_net_20994;
wire g61827_sb;
wire TIMEBOOST_net_107;
wire g61828_sb;
wire TIMEBOOST_net_20620;
wire TIMEBOOST_net_21634;
wire g61829_sb;
wire TIMEBOOST_net_403;
wire g61830_sb;
wire TIMEBOOST_net_11497;
wire g54194_db;
wire g61832_p;
wire g61833_p;
wire g61834_p;
wire g61835_sb;
wire TIMEBOOST_net_608;
wire g61836_sb;
wire TIMEBOOST_net_609;
wire g61837_db;
wire g61837_sb;
wire g61838_p;
wire g61839_p;
wire TIMEBOOST_net_769;
wire TIMEBOOST_net_14973;
wire g61840_sb;
wire TIMEBOOST_net_9193;
wire g61841_sb;
wire TIMEBOOST_net_13787;
wire g61842_sb;
wire TIMEBOOST_net_13684;
wire g61843_sb;
wire g61846_p;
wire g61850_p;
wire g61851_p;
wire TIMEBOOST_net_13754;
wire g61855_db;
wire g61855_sb;
wire TIMEBOOST_net_13751;
wire TIMEBOOST_net_13755;
wire g61856_sb;
wire g61857_p;
wire TIMEBOOST_net_536;
wire g61858_db;
wire g61858_sb;
wire n_4374;
wire g61859_db;
wire g61859_sb;
wire TIMEBOOST_net_16351;
wire g61860_sb;
wire TIMEBOOST_net_23410;
wire TIMEBOOST_net_404;
wire g61861_sb;
wire TIMEBOOST_net_405;
wire g61862_sb;
wire TIMEBOOST_net_538;
wire g61863_db;
wire g61863_sb;
wire TIMEBOOST_net_539;
wire g61864_db;
wire g61864_sb;
wire TIMEBOOST_net_9351;
wire g61865_sb;
wire TIMEBOOST_net_7548;
wire g61866_db;
wire g61866_sb;
wire TIMEBOOST_net_23334;
wire g61867_sb;
wire TIMEBOOST_net_20787;
wire TIMEBOOST_net_407;
wire g61868_sb;
wire TIMEBOOST_net_21653;
wire TIMEBOOST_net_408;
wire g61869_sb;
wire TIMEBOOST_net_13445;
wire g61870_db;
wire g61870_sb;
wire g61871_sb;
wire TIMEBOOST_net_14857;
wire TIMEBOOST_net_20926;
wire g61872_sb;
wire TIMEBOOST_net_22470;
wire g61873_sb;
wire TIMEBOOST_net_12466;
wire g61874_sb;
wire TIMEBOOST_net_412;
wire g61875_sb;
wire TIMEBOOST_net_16528;
wire g61876_sb;
wire TIMEBOOST_net_9352;
wire g61877_sb;
wire TIMEBOOST_net_736;
wire g61878_sb;
wire g61879_db;
wire g61879_sb;
wire TIMEBOOST_net_21848;
wire TIMEBOOST_net_9794;
wire g61880_sb;
wire TIMEBOOST_net_7611;
wire TIMEBOOST_net_414;
wire g61881_sb;
wire TIMEBOOST_net_20744;
wire TIMEBOOST_net_415;
wire g61882_sb;
wire TIMEBOOST_net_416;
wire g61883_sb;
wire TIMEBOOST_net_16010;
wire g61884_sb;
wire TIMEBOOST_net_14958;
wire TIMEBOOST_net_13580;
wire g61885_sb;
wire TIMEBOOST_net_10379;
wire g61886_sb;
wire TIMEBOOST_net_649;
wire g61887_db;
wire g61887_sb;
wire TIMEBOOST_net_418;
wire g61888_sb;
wire TIMEBOOST_net_650;
wire g61889_db;
wire g61889_sb;
wire TIMEBOOST_net_14870;
wire g61890_sb;
wire g61891_db;
wire g61891_sb;
wire TIMEBOOST_net_13604;
wire TIMEBOOST_net_420;
wire g61892_sb;
wire TIMEBOOST_net_9353;
wire g61893_sb;
wire TIMEBOOST_net_21971;
wire g61894_db;
wire g61894_sb;
wire TIMEBOOST_net_21972;
wire g61895_db;
wire g61895_sb;
wire TIMEBOOST_net_655;
wire g61896_db;
wire TIMEBOOST_net_664;
wire g61897_db;
wire g61897_sb;
wire TIMEBOOST_net_23218;
wire g61898_db;
wire TIMEBOOST_net_657;
wire g61899_db;
wire g61899_sb;
wire TIMEBOOST_net_13603;
wire TIMEBOOST_net_421;
wire g61900_sb;
wire TIMEBOOST_net_658;
wire TIMEBOOST_net_16439;
wire g61901_sb;
wire g61902_sb;
wire TIMEBOOST_net_9309;
wire g61903_sb;
wire TIMEBOOST_net_660;
wire g61904_db;
wire g61904_sb;
wire TIMEBOOST_net_422;
wire g61905_sb;
wire TIMEBOOST_net_17019;
wire TIMEBOOST_net_22250;
wire g61906_sb;
wire g61907_sb;
wire TIMEBOOST_net_176;
wire TIMEBOOST_net_5471;
wire g61908_sb;
wire TIMEBOOST_net_9310;
wire g61909_sb;
wire TIMEBOOST_net_17020;
wire TIMEBOOST_net_17012;
wire g61910_sb;
wire TIMEBOOST_net_13602;
wire g61911_sb;
wire TIMEBOOST_net_170;
wire g61912_sb;
wire g61913_sb;
wire TIMEBOOST_net_13600;
wire TIMEBOOST_net_10057;
wire g61914_sb;
wire TIMEBOOST_net_430;
wire g61915_sb;
wire TIMEBOOST_net_13596;
wire TIMEBOOST_net_431;
wire g61916_sb;
wire TIMEBOOST_net_12991;
wire g61917_sb;
wire TIMEBOOST_net_21180;
wire g61918_db;
wire g61918_sb;
wire g64912_db;
wire g61919_sb;
wire TIMEBOOST_net_22916;
wire g61920_db;
wire TIMEBOOST_net_14389;
wire g61921_sb;
wire TIMEBOOST_net_13447;
wire g61922_db;
wire TIMEBOOST_net_11498;
wire g61923_sb;
wire g61924_db;
wire g61924_sb;
wire g61925_db;
wire g61925_sb;
wire TIMEBOOST_net_21331;
wire g61926_sb;
wire TIMEBOOST_net_531;
wire TIMEBOOST_net_13884;
wire g61927_sb;
wire TIMEBOOST_net_22514;
wire g61928_db;
wire TIMEBOOST_net_13632;
wire g61929_sb;
wire TIMEBOOST_net_16004;
wire g61930_sb;
wire TIMEBOOST_net_284;
wire g61931_db;
wire g61931_sb;
wire TIMEBOOST_net_11599;
wire g61932_db;
wire g61932_sb;
wire TIMEBOOST_net_286;
wire g61933_db;
wire g61933_sb;
wire TIMEBOOST_net_287;
wire g61934_db;
wire g61934_sb;
wire TIMEBOOST_net_23436;
wire g61935_db;
wire g61936_sb;
wire TIMEBOOST_net_435;
wire g61937_sb;
wire TIMEBOOST_net_9706;
wire g61938_db;
wire TIMEBOOST_net_17278;
wire g61939_sb;
wire TIMEBOOST_net_14472;
wire g61940_sb;
wire TIMEBOOST_net_15419;
wire g61941_sb;
wire TIMEBOOST_net_21295;
wire TIMEBOOST_net_14007;
wire g61942_sb;
wire g61943_sb;
wire TIMEBOOST_net_21233;
wire TIMEBOOST_net_10110;
wire g61944_sb;
wire TIMEBOOST_net_23447;
wire TIMEBOOST_net_22526;
wire g61945_sb;
wire TIMEBOOST_net_13708;
wire TIMEBOOST_net_438;
wire g61946_sb;
wire TIMEBOOST_net_15659;
wire TIMEBOOST_net_21164;
wire g61947_sb;
wire TIMEBOOST_net_7113;
wire TIMEBOOST_net_16427;
wire g61948_sb;
wire TIMEBOOST_net_22498;
wire TIMEBOOST_net_12963;
wire g61949_sb;
wire TIMEBOOST_net_23487;
wire TIMEBOOST_net_14006;
wire g61950_sb;
wire g61951_sb;
wire TIMEBOOST_net_17317;
wire TIMEBOOST_net_17470;
wire g61952_sb;
wire TIMEBOOST_net_12259;
wire g61953_db;
wire TIMEBOOST_net_8004;
wire TIMEBOOST_net_16767;
wire g61954_sb;
wire TIMEBOOST_net_16861;
wire TIMEBOOST_net_14797;
wire g61955_sb;
wire TIMEBOOST_net_21167;
wire g61956_db;
wire g61956_sb;
wire g61957_sb;
wire TIMEBOOST_net_20798;
wire g61958_sb;
wire g61959_db;
wire g61959_sb;
wire TIMEBOOST_net_21786;
wire TIMEBOOST_net_13582;
wire g61961_sb;
wire TIMEBOOST_net_20218;
wire g61962_sb;
wire TIMEBOOST_net_12984;
wire g61963_sb;
wire g61964_db;
wire TIMEBOOST_net_22191;
wire g61965_db;
wire g61965_sb;
wire TIMEBOOST_net_20253;
wire TIMEBOOST_net_13678;
wire TIMEBOOST_net_20254;
wire TIMEBOOST_net_13677;
wire TIMEBOOST_net_10832;
wire TIMEBOOST_net_21928;
wire g61969_db;
wire TIMEBOOST_net_17425;
wire TIMEBOOST_net_11480;
wire TIMEBOOST_net_21710;
wire g54489_da;
wire TIMEBOOST_net_13714;
wire TIMEBOOST_net_14570;
wire TIMEBOOST_net_16792;
wire TIMEBOOST_net_12736;
wire TIMEBOOST_net_745;
wire n_4383;
wire TIMEBOOST_net_16793;
wire TIMEBOOST_net_13703;
wire TIMEBOOST_net_16789;
wire TIMEBOOST_net_12546;
wire TIMEBOOST_net_21374;
wire TIMEBOOST_net_17369;
wire TIMEBOOST_net_16794;
wire TIMEBOOST_net_16795;
wire TIMEBOOST_net_17364;
wire TIMEBOOST_net_16796;
wire TIMEBOOST_net_13574;
wire TIMEBOOST_net_11477;
wire TIMEBOOST_net_20431;
wire TIMEBOOST_net_20255;
wire TIMEBOOST_net_13583;
wire TIMEBOOST_net_11478;
wire TIMEBOOST_net_20460;
wire TIMEBOOST_net_748;
wire TIMEBOOST_net_13619;
wire TIMEBOOST_net_11479;
wire TIMEBOOST_net_14324;
wire g61990_db;
wire g61990_sb;
wire TIMEBOOST_net_7619;
wire g61991_sb;
wire TIMEBOOST_net_21531;
wire g61992_db;
wire g61992_sb;
wire g61993_sb;
wire TIMEBOOST_net_14473;
wire g61994_sb;
wire TIMEBOOST_net_21155;
wire TIMEBOOST_net_17583;
wire g61995_sb;
wire TIMEBOOST_net_22017;
wire g61996_db;
wire TIMEBOOST_net_23267;
wire g61997_db;
wire g61997_sb;
wire TIMEBOOST_net_14736;
wire g61998_sb;
wire TIMEBOOST_net_14325;
wire g61999_db;
wire g61999_sb;
wire TIMEBOOST_net_532;
wire g62000_db;
wire g62000_sb;
wire TIMEBOOST_net_14794;
wire g62001_sb;
wire g62002_sb;
wire g62003_db;
wire g62003_sb;
wire TIMEBOOST_net_22545;
wire g62004_db;
wire g62005_sb;
wire TIMEBOOST_net_21943;
wire TIMEBOOST_net_448;
wire g62006_sb;
wire TIMEBOOST_net_23471;
wire g62007_db;
wire g62007_sb;
wire g62008_db;
wire TIMEBOOST_net_20896;
wire TIMEBOOST_net_449;
wire g62009_sb;
wire g62010_sb;
wire TIMEBOOST_net_21022;
wire TIMEBOOST_net_451;
wire g62011_sb;
wire TIMEBOOST_net_13555;
wire g62012_db;
wire g62012_sb;
wire TIMEBOOST_net_452;
wire g62013_sb;
wire TIMEBOOST_net_582;
wire g62014_sb;
wire TIMEBOOST_net_21769;
wire TIMEBOOST_net_453;
wire g62015_sb;
wire TIMEBOOST_net_14841;
wire TIMEBOOST_net_454;
wire g62016_sb;
wire TIMEBOOST_net_7618;
wire TIMEBOOST_net_603;
wire g62017_sb;
wire TIMEBOOST_net_534;
wire TIMEBOOST_net_14954;
wire g62018_sb;
wire TIMEBOOST_net_7617;
wire TIMEBOOST_net_14371;
wire g62019_sb;
wire TIMEBOOST_net_22523;
wire g62020_sb;
wire TIMEBOOST_net_16797;
wire TIMEBOOST_net_12574;
wire TIMEBOOST_net_455;
wire g62022_sb;
wire TIMEBOOST_net_7616;
wire g62023_sb;
wire g62024_sb;
wire TIMEBOOST_net_21002;
wire g62025_sb;
wire TIMEBOOST_net_7615;
wire g62026_sb;
wire g62027_sb;
wire TIMEBOOST_net_12370;
wire g62028_sb;
wire TIMEBOOST_net_14892;
wire TIMEBOOST_net_22441;
wire g62029_sb;
wire g62030_da;
wire g62030_db;
wire g62030_sb;
wire TIMEBOOST_net_15460;
wire g62031_sb;
wire TIMEBOOST_net_5516;
wire g52470_da;
wire g62032_sb;
wire TIMEBOOST_net_20245;
wire TIMEBOOST_net_8278;
wire g62033_sb;
wire g52457_da;
wire g62034_sb;
wire TIMEBOOST_net_10282;
wire g62035_sb;
wire TIMEBOOST_net_23543;
wire g62036_sb;
wire g62037_sb;
wire TIMEBOOST_net_11461;
wire g62038_sb;
wire TIMEBOOST_net_10268;
wire TIMEBOOST_net_11462;
wire g62039_sb;
wire n_9099;
wire g62040_sb;
wire g62041_sb;
wire TIMEBOOST_net_23398;
wire TIMEBOOST_net_15798;
wire g62042_sb;
wire TIMEBOOST_net_8785;
wire g62043_sb;
wire g62044_sb;
wire TIMEBOOST_net_16529;
wire g62045_sb;
wire TIMEBOOST_net_5529;
wire g62046_sb;
wire g62047_sb;
wire TIMEBOOST_net_14609;
wire TIMEBOOST_net_11430;
wire g62048_sb;
wire TIMEBOOST_net_16600;
wire TIMEBOOST_net_21395;
wire g62049_sb;
wire TIMEBOOST_net_5533;
wire g62050_sb;
wire TIMEBOOST_net_15078;
wire g62051_sb;
wire TIMEBOOST_net_15079;
wire g62052_sb;
wire g62053_sb;
wire TIMEBOOST_net_15194;
wire TIMEBOOST_net_15081;
wire g62054_sb;
wire TIMEBOOST_net_15082;
wire g62055_sb;
wire TIMEBOOST_net_21221;
wire g62056_sb;
wire TIMEBOOST_net_9521;
wire TIMEBOOST_net_20785;
wire g62057_sb;
wire g65781_da;
wire g61976_db;
wire g62058_sb;
wire TIMEBOOST_net_16007;
wire TIMEBOOST_net_15085;
wire g62059_sb;
wire TIMEBOOST_net_5542;
wire TIMEBOOST_net_15086;
wire g62060_sb;
wire TIMEBOOST_net_15087;
wire g62061_sb;
wire TIMEBOOST_net_9700;
wire TIMEBOOST_net_21311;
wire g62062_sb;
wire TIMEBOOST_net_9589;
wire g62063_sb;
wire TIMEBOOST_net_21281;
wire g62064_sb;
wire TIMEBOOST_net_22748;
wire TIMEBOOST_net_21299;
wire g62065_sb;
wire TIMEBOOST_net_21770;
wire TIMEBOOST_net_461;
wire g62066_sb;
wire TIMEBOOST_net_13625;
wire TIMEBOOST_net_9503;
wire g62067_sb;
wire TIMEBOOST_net_22894;
wire g62068_db;
wire g62068_sb;
wire TIMEBOOST_net_21661;
wire TIMEBOOST_net_21259;
wire g62069_sb;
wire TIMEBOOST_net_22079;
wire TIMEBOOST_net_463;
wire g62070_sb;
wire TIMEBOOST_net_21610;
wire TIMEBOOST_net_16787;
wire g62071_sb;
wire TIMEBOOST_net_546;
wire TIMEBOOST_net_16512;
wire g62072_sb;
wire TIMEBOOST_net_20760;
wire TIMEBOOST_net_665;
wire g62073_sb;
wire TIMEBOOST_net_23272;
wire TIMEBOOST_net_666;
wire g62074_sb;
wire TIMEBOOST_net_21136;
wire g62075_sb;
wire TIMEBOOST_net_140;
wire TIMEBOOST_net_668;
wire g62076_sb;
wire TIMEBOOST_net_547;
wire TIMEBOOST_net_14299;
wire g62077_sb;
wire TIMEBOOST_net_14310;
wire g62078_sb;
wire TIMEBOOST_net_13784;
wire g62079_sb;
wire TIMEBOOST_net_21419;
wire TIMEBOOST_net_670;
wire g62080_sb;
wire TIMEBOOST_net_21729;
wire TIMEBOOST_net_14486;
wire g62081_sb;
wire TIMEBOOST_net_22957;
wire TIMEBOOST_net_16173;
wire g62082_sb;
wire g62083_sb;
wire TIMEBOOST_net_674;
wire g62084_sb;
wire TIMEBOOST_net_16995;
wire g62085_sb;
wire TIMEBOOST_net_16994;
wire TIMEBOOST_net_7094;
wire g62086_sb;
wire g62087_sb;
wire TIMEBOOST_net_22901;
wire g62088_sb;
wire TIMEBOOST_net_23193;
wire TIMEBOOST_net_22612;
wire g62089_sb;
wire TIMEBOOST_net_22501;
wire TIMEBOOST_net_14309;
wire g62090_sb;
wire TIMEBOOST_net_7587;
wire g62091_sb;
wire TIMEBOOST_net_681;
wire g62092_sb;
wire g62093_sb;
wire TIMEBOOST_net_15414;
wire g62094_sb;
wire TIMEBOOST_net_551;
wire TIMEBOOST_net_16420;
wire g62095_sb;
wire n_2389;
wire g62096_sb;
wire TIMEBOOST_net_7584;
wire TIMEBOOST_net_683;
wire g62097_sb;
wire TIMEBOOST_net_20466;
wire TIMEBOOST_net_684;
wire g62098_sb;
wire TIMEBOOST_net_14140;
wire TIMEBOOST_net_685;
wire g62099_sb;
wire TIMEBOOST_net_14139;
wire g62100_sb;
wire TIMEBOOST_net_20934;
wire TIMEBOOST_net_22843;
wire g62101_sb;
wire TIMEBOOST_net_20137;
wire TIMEBOOST_net_5515;
wire g62102_sb;
wire TIMEBOOST_net_14160;
wire TIMEBOOST_net_688;
wire g62103_sb;
wire TIMEBOOST_net_13873;
wire TIMEBOOST_net_689;
wire g62104_sb;
wire TIMEBOOST_net_23498;
wire g62105_sb;
wire TIMEBOOST_net_553;
wire g62106_db;
wire g62106_sb;
wire TIMEBOOST_net_691;
wire g62107_sb;
wire TIMEBOOST_net_692;
wire g62108_sb;
wire TIMEBOOST_net_119;
wire TIMEBOOST_net_693;
wire g62109_sb;
wire TIMEBOOST_net_21736;
wire TIMEBOOST_net_694;
wire g62110_sb;
wire TIMEBOOST_net_22319;
wire g62111_db;
wire g62111_sb;
wire TIMEBOOST_net_543;
wire TIMEBOOST_net_695;
wire g62112_sb;
wire TIMEBOOST_net_21533;
wire TIMEBOOST_net_696;
wire g62113_sb;
wire TIMEBOOST_net_555;
wire g62114_db;
wire g62114_sb;
wire TIMEBOOST_net_697;
wire g62115_sb;
wire TIMEBOOST_net_16478;
wire TIMEBOOST_net_23521;
wire g62116_sb;
wire g64963_db;
wire TIMEBOOST_net_698;
wire g62117_sb;
wire TIMEBOOST_net_699;
wire g62118_sb;
wire TIMEBOOST_net_557;
wire g62119_db;
wire g62119_sb;
wire TIMEBOOST_net_700;
wire g62120_sb;
wire TIMEBOOST_net_21615;
wire TIMEBOOST_net_701;
wire g62121_sb;
wire TIMEBOOST_net_21691;
wire TIMEBOOST_net_702;
wire g62122_sb;
wire TIMEBOOST_net_12027;
wire TIMEBOOST_net_703;
wire g62123_sb;
wire TIMEBOOST_net_558;
wire g62124_sb;
wire TIMEBOOST_net_704;
wire g62125_sb;
wire TIMEBOOST_net_705;
wire g62126_sb;
wire TIMEBOOST_net_706;
wire g62127_sb;
wire TIMEBOOST_net_707;
wire g62128_sb;
wire g57798_da;
wire TIMEBOOST_net_708;
wire g62129_sb;
wire TIMEBOOST_net_709;
wire g62130_sb;
wire TIMEBOOST_net_23033;
wire TIMEBOOST_net_710;
wire g62131_sb;
wire TIMEBOOST_net_23469;
wire g62132_sb;
wire TIMEBOOST_net_13954;
wire TIMEBOOST_net_17478;
wire g62133_sb;
wire TIMEBOOST_net_14005;
wire g62134_db;
wire g62134_sb;
wire TIMEBOOST_net_13834;
wire TIMEBOOST_net_711;
wire g62135_sb;
wire TIMEBOOST_net_712;
wire g62136_sb;
wire TIMEBOOST_net_23268;
wire TIMEBOOST_net_713;
wire g62137_sb;
wire TIMEBOOST_net_16907;
wire g62138_sb;
wire g62139_sb;
wire TIMEBOOST_net_22577;
wire g62140_sb;
wire g62141_sb;
wire g62219_p;
wire g62220_p;
wire g62221_p;
wire g62223_p;
wire g62254_p;
wire g62264_p;
wire g62285_p;
wire g62312_p;
wire g62318_p;
wire g62319_p;
wire TIMEBOOST_net_10912;
wire g62326_db;
wire g62326_sb;
wire TIMEBOOST_net_16865;
wire TIMEBOOST_net_11211;
wire g62333_sb;
wire TIMEBOOST_net_16863;
wire g62334_sb;
wire TIMEBOOST_net_16862;
wire g62335_sb;
wire TIMEBOOST_net_11863;
wire TIMEBOOST_net_13235;
wire g62336_sb;
wire TIMEBOOST_net_10047;
wire TIMEBOOST_net_11133;
wire g62337_sb;
wire TIMEBOOST_net_10046;
wire TIMEBOOST_net_15227;
wire g62338_sb;
wire TIMEBOOST_net_10045;
wire g62339_sb;
wire g62340_sb;
wire TIMEBOOST_net_17184;
wire g62341_sb;
wire g62342_sb;
wire TIMEBOOST_net_15708;
wire TIMEBOOST_net_23557;
wire g62343_sb;
wire TIMEBOOST_net_10884;
wire g62344_sb;
wire TIMEBOOST_net_16698;
wire g62345_sb;
wire g62346_sb;
wire g62347_sb;
wire g62348_sb;
wire TIMEBOOST_net_23433;
wire g62349_sb;
wire TIMEBOOST_net_21751;
wire g62350_sb;
wire TIMEBOOST_net_10391;
wire TIMEBOOST_net_16699;
wire g62351_sb;
wire TIMEBOOST_net_23310;
wire g62352_sb;
wire TIMEBOOST_net_13624;
wire n_12116;
wire g62353_sb;
wire TIMEBOOST_net_21427;
wire g62354_sb;
wire TIMEBOOST_net_21574;
wire g62355_sb;
wire TIMEBOOST_net_7532;
wire g62356_sb;
wire TIMEBOOST_net_13556;
wire g62357_sb;
wire g62358_sb;
wire TIMEBOOST_net_7508;
wire TIMEBOOST_net_11178;
wire g62359_sb;
wire TIMEBOOST_net_13566;
wire TIMEBOOST_net_16762;
wire g62360_sb;
wire TIMEBOOST_net_22261;
wire g62361_sb;
wire TIMEBOOST_net_17291;
wire TIMEBOOST_net_10133;
wire g62362_sb;
wire TIMEBOOST_net_21740;
wire g62363_sb;
wire TIMEBOOST_net_13599;
wire TIMEBOOST_net_11195;
wire g62364_sb;
wire g62365_sb;
wire g62366_db;
wire g62366_sb;
wire TIMEBOOST_net_21592;
wire TIMEBOOST_net_21202;
wire g62367_sb;
wire g62368_sb;
wire TIMEBOOST_net_11196;
wire g62369_sb;
wire TIMEBOOST_net_22317;
wire TIMEBOOST_net_17516;
wire g62370_sb;
wire TIMEBOOST_net_20844;
wire TIMEBOOST_net_11197;
wire g62371_sb;
wire g64866_db;
wire TIMEBOOST_net_11198;
wire g62372_sb;
wire TIMEBOOST_net_22904;
wire TIMEBOOST_net_23426;
wire g62373_sb;
wire TIMEBOOST_net_12039;
wire g62374_sb;
wire TIMEBOOST_net_5638;
wire g62375_sb;
wire TIMEBOOST_net_14003;
wire g62376_sb;
wire TIMEBOOST_net_14919;
wire TIMEBOOST_net_21147;
wire g62377_sb;
wire TIMEBOOST_net_17517;
wire g62378_sb;
wire TIMEBOOST_net_21278;
wire g62379_sb;
wire TIMEBOOST_net_14751;
wire g62380_sb;
wire TIMEBOOST_net_15063;
wire TIMEBOOST_net_17419;
wire g62381_sb;
wire TIMEBOOST_net_15431;
wire TIMEBOOST_net_14972;
wire g62382_sb;
wire TIMEBOOST_net_5642;
wire TIMEBOOST_net_17573;
wire g62383_sb;
wire TIMEBOOST_net_5643;
wire TIMEBOOST_net_17574;
wire g62384_sb;
wire TIMEBOOST_net_5644;
wire TIMEBOOST_net_17575;
wire g62385_sb;
wire TIMEBOOST_net_14710;
wire TIMEBOOST_net_17576;
wire g62386_sb;
wire TIMEBOOST_net_13188;
wire TIMEBOOST_net_10902;
wire g62387_sb;
wire TIMEBOOST_net_22922;
wire g62388_sb;
wire TIMEBOOST_net_10892;
wire g62389_sb;
wire g62390_sb;
wire TIMEBOOST_net_17486;
wire g62391_sb;
wire TIMEBOOST_net_12537;
wire g62392_sb;
wire TIMEBOOST_net_14175;
wire TIMEBOOST_net_17028;
wire g62393_sb;
wire TIMEBOOST_net_21407;
wire g62394_sb;
wire TIMEBOOST_net_16705;
wire g62395_sb;
wire TIMEBOOST_net_10026;
wire g62396_sb;
wire g62397_sb;
wire g62398_sb;
wire TIMEBOOST_net_14207;
wire TIMEBOOST_net_23440;
wire g62399_sb;
wire TIMEBOOST_net_21178;
wire g62400_sb;
wire TIMEBOOST_net_16703;
wire g62401_sb;
wire TIMEBOOST_net_10019;
wire TIMEBOOST_net_11171;
wire g62402_sb;
wire TIMEBOOST_net_10018;
wire g62403_sb;
wire TIMEBOOST_net_21272;
wire g62404_sb;
wire TIMEBOOST_net_17406;
wire g62405_sb;
wire TIMEBOOST_net_10801;
wire g62406_sb;
wire TIMEBOOST_net_10327;
wire TIMEBOOST_net_16704;
wire g62407_sb;
wire TIMEBOOST_net_17027;
wire TIMEBOOST_net_16706;
wire g62408_sb;
wire TIMEBOOST_net_21821;
wire TIMEBOOST_net_11102;
wire g62409_sb;
wire g62410_sb;
wire TIMEBOOST_net_12678;
wire g62411_sb;
wire TIMEBOOST_net_14215;
wire g62412_sb;
wire g52467_da;
wire g62413_sb;
wire TIMEBOOST_net_23402;
wire g62414_sb;
wire TIMEBOOST_net_8271;
wire g62415_sb;
wire TIMEBOOST_net_10325;
wire TIMEBOOST_net_16701;
wire g62416_sb;
wire TIMEBOOST_net_5664;
wire g62417_sb;
wire g62418_sb;
wire TIMEBOOST_net_5666;
wire g62419_sb;
wire TIMEBOOST_net_5667;
wire g62420_sb;
wire TIMEBOOST_net_10013;
wire g62421_sb;
wire TIMEBOOST_net_5668;
wire g62422_sb;
wire TIMEBOOST_net_21218;
wire TIMEBOOST_net_5500;
wire g62423_sb;
wire TIMEBOOST_net_23362;
wire TIMEBOOST_net_21834;
wire g62424_sb;
wire TIMEBOOST_net_10324;
wire TIMEBOOST_net_16702;
wire g62425_sb;
wire g62426_sb;
wire TIMEBOOST_net_10323;
wire TIMEBOOST_net_16700;
wire g62427_sb;
wire TIMEBOOST_net_10918;
wire TIMEBOOST_net_13615;
wire g62428_sb;
wire g62429_sb;
wire g62430_sb;
wire TIMEBOOST_net_14689;
wire g62431_sb;
wire TIMEBOOST_net_10009;
wire g62432_sb;
wire TIMEBOOST_net_10390;
wire TIMEBOOST_net_16696;
wire g62433_sb;
wire TIMEBOOST_net_17358;
wire g62434_sb;
wire TIMEBOOST_net_20511;
wire g62435_sb;
wire TIMEBOOST_net_8784;
wire g62436_sb;
wire TIMEBOOST_net_8783;
wire g62437_sb;
wire g62438_sb;
wire TIMEBOOST_net_17082;
wire TIMEBOOST_net_23095;
wire g62439_sb;
wire TIMEBOOST_net_9327;
wire g62440_sb;
wire TIMEBOOST_net_17357;
wire g62441_sb;
wire g62442_sb;
wire TIMEBOOST_net_12993;
wire TIMEBOOST_net_16998;
wire g62443_sb;
wire TIMEBOOST_net_10389;
wire TIMEBOOST_net_14648;
wire g62444_sb;
wire TIMEBOOST_net_13373;
wire g62445_sb;
wire g62446_sb;
wire TIMEBOOST_net_21619;
wire g62447_sb;
wire g62448_sb;
wire TIMEBOOST_net_15167;
wire g62449_sb;
wire g54239_db;
wire g52483_da;
wire g62450_sb;
wire TIMEBOOST_net_10321;
wire TIMEBOOST_net_15054;
wire g62451_sb;
wire TIMEBOOST_net_17093;
wire g62452_sb;
wire TIMEBOOST_net_10631;
wire g62453_sb;
wire g62454_sb;
wire TIMEBOOST_net_17515;
wire g62455_sb;
wire TIMEBOOST_net_17353;
wire TIMEBOOST_net_16053;
wire g62456_sb;
wire TIMEBOOST_net_14618;
wire g62457_sb;
wire g62458_sb;
wire TIMEBOOST_net_5685;
wire TIMEBOOST_net_23448;
wire g62459_sb;
wire TIMEBOOST_net_5686;
wire TIMEBOOST_net_15954;
wire g62460_sb;
wire TIMEBOOST_net_10988;
wire g62461_sb;
wire TIMEBOOST_net_9465;
wire TIMEBOOST_net_10890;
wire g62462_sb;
wire TIMEBOOST_net_9466;
wire TIMEBOOST_net_23441;
wire g62463_sb;
wire TIMEBOOST_net_9464;
wire g62464_sb;
wire TIMEBOOST_net_10991;
wire g62465_sb;
wire TIMEBOOST_net_9446;
wire g62466_sb;
wire TIMEBOOST_net_9451;
wire g62467_sb;
wire TIMEBOOST_net_5435;
wire g62468_sb;
wire TIMEBOOST_net_11015;
wire g62469_sb;
wire TIMEBOOST_net_9452;
wire TIMEBOOST_net_16763;
wire g62470_sb;
wire TIMEBOOST_net_9438;
wire TIMEBOOST_net_11192;
wire g62471_sb;
wire TIMEBOOST_net_14642;
wire g62472_sb;
wire TIMEBOOST_net_14641;
wire TIMEBOOST_net_17532;
wire g62473_sb;
wire TIMEBOOST_net_9439;
wire TIMEBOOST_net_11193;
wire g62474_sb;
wire TIMEBOOST_net_14640;
wire g62475_sb;
wire TIMEBOOST_net_9442;
wire TIMEBOOST_net_17402;
wire g62476_sb;
wire TIMEBOOST_net_10320;
wire TIMEBOOST_net_10632;
wire g62477_sb;
wire g62478_sb;
wire TIMEBOOST_net_10921;
wire TIMEBOOST_net_9609;
wire g62479_sb;
wire TIMEBOOST_net_21538;
wire g62480_sb;
wire TIMEBOOST_net_20302;
wire g62481_sb;
wire TIMEBOOST_net_9448;
wire g62482_sb;
wire TIMEBOOST_net_9463;
wire n_12115;
wire g62483_sb;
wire TIMEBOOST_net_10319;
wire TIMEBOOST_net_10633;
wire g62484_sb;
wire TIMEBOOST_net_9450;
wire TIMEBOOST_net_23431;
wire g62485_sb;
wire TIMEBOOST_net_10386;
wire TIMEBOOST_net_17257;
wire g62486_sb;
wire TIMEBOOST_net_9444;
wire g62487_sb;
wire TIMEBOOST_net_9443;
wire g62488_sb;
wire TIMEBOOST_net_9467;
wire g62489_sb;
wire TIMEBOOST_net_9447;
wire g62490_sb;
wire TIMEBOOST_net_13626;
wire g62491_sb;
wire TIMEBOOST_net_9440;
wire g62492_sb;
wire TIMEBOOST_net_14636;
wire g62493_sb;
wire TIMEBOOST_net_9453;
wire g62494_sb;
wire TIMEBOOST_net_16750;
wire TIMEBOOST_net_21026;
wire g62495_sb;
wire TIMEBOOST_net_9449;
wire n_12369;
wire g62496_sb;
wire TIMEBOOST_net_9441;
wire g62497_sb;
wire TIMEBOOST_net_17066;
wire g62498_sb;
wire TIMEBOOST_net_9470;
wire g62499_sb;
wire TIMEBOOST_net_9445;
wire g62500_sb;
wire TIMEBOOST_net_10318;
wire FE_RN_540_0;
wire g62501_sb;
wire TIMEBOOST_net_9437;
wire g62502_sb;
wire TIMEBOOST_net_9468;
wire n_12372;
wire g62503_sb;
wire TIMEBOOST_net_14288;
wire TIMEBOOST_net_20627;
wire g62504_sb;
wire TIMEBOOST_net_9469;
wire g62505_sb;
wire TIMEBOOST_net_9462;
wire g62506_sb;
wire TIMEBOOST_net_10923;
wire g62507_sb;
wire TIMEBOOST_net_9461;
wire g62508_sb;
wire TIMEBOOST_net_9460;
wire g62509_sb;
wire TIMEBOOST_net_9459;
wire g62510_sb;
wire TIMEBOOST_net_14647;
wire g62511_sb;
wire TIMEBOOST_net_20961;
wire TIMEBOOST_net_5504;
wire g62512_sb;
wire g62513_sb;
wire TIMEBOOST_net_9458;
wire TIMEBOOST_net_14994;
wire g62514_sb;
wire TIMEBOOST_net_9457;
wire TIMEBOOST_net_11174;
wire g62515_sb;
wire TIMEBOOST_net_10926;
wire g62516_db;
wire g62516_sb;
wire TIMEBOOST_net_9608;
wire g62517_sb;
wire TIMEBOOST_net_16615;
wire g62518_sb;
wire g62519_sb;
wire TIMEBOOST_net_8733;
wire TIMEBOOST_net_16616;
wire g62520_sb;
wire TIMEBOOST_net_9456;
wire TIMEBOOST_net_21205;
wire g62521_sb;
wire TIMEBOOST_net_9455;
wire g62522_sb;
wire TIMEBOOST_net_8732;
wire TIMEBOOST_net_16617;
wire g62523_sb;
wire TIMEBOOST_net_5720;
wire TIMEBOOST_net_11146;
wire g62524_sb;
wire TIMEBOOST_net_13514;
wire g62525_sb;
wire TIMEBOOST_net_13513;
wire g62526_sb;
wire TIMEBOOST_net_9454;
wire g62527_sb;
wire TIMEBOOST_net_10051;
wire g62528_sb;
wire TIMEBOOST_net_17489;
wire g62529_sb;
wire TIMEBOOST_net_9534;
wire g62530_sb;
wire TIMEBOOST_net_9533;
wire g62531_sb;
wire TIMEBOOST_net_17032;
wire TIMEBOOST_net_17487;
wire g62532_sb;
wire g62533_sb;
wire TIMEBOOST_net_10234;
wire g62534_sb;
wire TIMEBOOST_net_17259;
wire g62535_sb;
wire TIMEBOOST_net_9532;
wire g62536_sb;
wire TIMEBOOST_net_9531;
wire TIMEBOOST_net_16951;
wire g62537_sb;
wire TIMEBOOST_net_9510;
wire g62538_sb;
wire TIMEBOOST_net_9528;
wire g62539_sb;
wire TIMEBOOST_net_10233;
wire g62540_sb;
wire TIMEBOOST_net_9520;
wire TIMEBOOST_net_16760;
wire g62541_sb;
wire TIMEBOOST_net_9517;
wire g62542_sb;
wire TIMEBOOST_net_9514;
wire g62543_sb;
wire TIMEBOOST_net_9529;
wire g62544_sb;
wire TIMEBOOST_net_9526;
wire TIMEBOOST_net_20791;
wire g62545_sb;
wire TIMEBOOST_net_9525;
wire g62546_sb;
wire TIMEBOOST_net_16619;
wire g62547_sb;
wire TIMEBOOST_net_9522;
wire TIMEBOOST_net_11033;
wire g62548_sb;
wire TIMEBOOST_net_9518;
wire TIMEBOOST_net_17405;
wire g62549_sb;
wire TIMEBOOST_net_17286;
wire TIMEBOOST_net_17557;
wire g62550_sb;
wire g52485_da;
wire g62551_sb;
wire g62552_sb;
wire TIMEBOOST_net_10203;
wire TIMEBOOST_net_17558;
wire g62553_sb;
wire TIMEBOOST_net_9516;
wire g62554_sb;
wire TIMEBOOST_net_5739;
wire TIMEBOOST_net_17553;
wire g62555_sb;
wire TIMEBOOST_net_9511;
wire TIMEBOOST_net_10765;
wire g62556_sb;
wire TIMEBOOST_net_9543;
wire g62557_sb;
wire TIMEBOOST_net_16620;
wire g62558_sb;
wire g62559_sb;
wire TIMEBOOST_net_21204;
wire TIMEBOOST_net_16621;
wire g62560_sb;
wire TIMEBOOST_net_8725;
wire g62561_sb;
wire TIMEBOOST_net_22150;
wire g61983_db;
wire g62562_sb;
wire TIMEBOOST_net_14916;
wire g62563_sb;
wire TIMEBOOST_net_9542;
wire g62564_sb;
wire TIMEBOOST_net_9541;
wire TIMEBOOST_net_10764;
wire g62565_sb;
wire TIMEBOOST_net_9540;
wire g62566_sb;
wire TIMEBOOST_net_9539;
wire TIMEBOOST_net_17529;
wire g62567_sb;
wire TIMEBOOST_net_9524;
wire g62568_sb;
wire TIMEBOOST_net_16624;
wire g62569_sb;
wire TIMEBOOST_net_16960;
wire g62570_sb;
wire n_3932;
wire TIMEBOOST_net_16625;
wire g62571_sb;
wire TIMEBOOST_net_9513;
wire g62572_sb;
wire TIMEBOOST_net_9512;
wire g62573_sb;
wire TIMEBOOST_net_9527;
wire TIMEBOOST_net_11170;
wire g62574_sb;
wire TIMEBOOST_net_20750;
wire g62575_sb;
wire g62576_sb;
wire TIMEBOOST_net_9557;
wire TIMEBOOST_net_11101;
wire g62577_sb;
wire TIMEBOOST_net_9555;
wire TIMEBOOST_net_17401;
wire g62578_sb;
wire TIMEBOOST_net_9552;
wire TIMEBOOST_net_17409;
wire g62579_sb;
wire g62580_db;
wire g62580_sb;
wire TIMEBOOST_net_9551;
wire TIMEBOOST_net_11106;
wire g62581_sb;
wire TIMEBOOST_net_9550;
wire TIMEBOOST_net_17410;
wire g62582_sb;
wire g62583_sb;
wire TIMEBOOST_net_9549;
wire TIMEBOOST_net_17420;
wire g62584_sb;
wire TIMEBOOST_net_9547;
wire g62585_sb;
wire TIMEBOOST_net_9544;
wire TIMEBOOST_net_11114;
wire g62586_sb;
wire TIMEBOOST_net_9556;
wire g62587_sb;
wire TIMEBOOST_net_17017;
wire g62588_sb;
wire TIMEBOOST_net_9545;
wire TIMEBOOST_net_17510;
wire g62589_sb;
wire TIMEBOOST_net_9530;
wire TIMEBOOST_net_17485;
wire g62590_sb;
wire TIMEBOOST_net_9523;
wire TIMEBOOST_net_16135;
wire g62591_sb;
wire TIMEBOOST_net_10347;
wire g62592_sb;
wire TIMEBOOST_net_8720;
wire TIMEBOOST_net_16626;
wire g62593_sb;
wire TIMEBOOST_net_9554;
wire g62594_sb;
wire g62595_p;
wire TIMEBOOST_net_9553;
wire TIMEBOOST_net_11084;
wire g62596_sb;
wire TIMEBOOST_net_9515;
wire g62597_sb;
wire TIMEBOOST_net_9559;
wire TIMEBOOST_net_22209;
wire g62598_sb;
wire TIMEBOOST_net_17288;
wire g62599_sb;
wire TIMEBOOST_net_22517;
wire g62600_sb;
wire TIMEBOOST_net_17559;
wire g62601_sb;
wire TIMEBOOST_net_9558;
wire TIMEBOOST_net_23330;
wire g62602_sb;
wire TIMEBOOST_net_9548;
wire TIMEBOOST_net_11103;
wire g62603_sb;
wire TIMEBOOST_net_13535;
wire TIMEBOOST_net_17561;
wire g62604_sb;
wire TIMEBOOST_net_21187;
wire TIMEBOOST_net_5509;
wire g62605_sb;
wire TIMEBOOST_net_10182;
wire g62606_sb;
wire TIMEBOOST_net_11451;
wire g62607_sb;
wire TIMEBOOST_net_9546;
wire g62608_sb;
wire TIMEBOOST_net_9519;
wire g62609_sb;
wire TIMEBOOST_net_9538;
wire TIMEBOOST_net_10989;
wire g62610_sb;
wire TIMEBOOST_net_20793;
wire g62611_db;
wire g62611_sb;
wire g62612_sb;
wire TIMEBOOST_net_9537;
wire TIMEBOOST_net_11166;
wire g62613_sb;
wire TIMEBOOST_net_10178;
wire g62614_sb;
wire TIMEBOOST_net_9536;
wire g62615_sb;
wire TIMEBOOST_net_9535;
wire g62616_sb;
wire TIMEBOOST_net_13167;
wire g62617_sb;
wire TIMEBOOST_net_10317;
wire g62618_sb;
wire TIMEBOOST_net_10175;
wire g62619_sb;
wire TIMEBOOST_net_23166;
wire g62620_sb;
wire TIMEBOOST_net_20746;
wire g62621_sb;
wire TIMEBOOST_net_10316;
wire TIMEBOOST_net_16630;
wire g62622_sb;
wire TIMEBOOST_net_20982;
wire TIMEBOOST_net_17560;
wire g62623_sb;
wire TIMEBOOST_net_21411;
wire TIMEBOOST_net_10893;
wire g62624_sb;
wire TIMEBOOST_net_10167;
wire g62625_sb;
wire TIMEBOOST_net_10165;
wire TIMEBOOST_net_10760;
wire g62626_sb;
wire TIMEBOOST_net_16742;
wire TIMEBOOST_net_10206;
wire g62627_sb;
wire TIMEBOOST_net_15371;
wire g62628_sb;
wire TIMEBOOST_net_23082;
wire g62629_sb;
wire TIMEBOOST_net_10164;
wire TIMEBOOST_net_10788;
wire g62630_sb;
wire TIMEBOOST_net_13075;
wire g62631_sb;
wire g62632_sb;
wire TIMEBOOST_net_16631;
wire g62633_sb;
wire TIMEBOOST_net_17398;
wire g62634_sb;
wire g62635_sb;
wire TIMEBOOST_net_16633;
wire g62636_sb;
wire TIMEBOOST_net_10895;
wire g62637_sb;
wire TIMEBOOST_net_13073;
wire TIMEBOOST_net_10896;
wire g62638_sb;
wire TIMEBOOST_net_21263;
wire TIMEBOOST_net_10897;
wire g62639_sb;
wire TIMEBOOST_net_10898;
wire g62640_sb;
wire g62641_sb;
wire TIMEBOOST_net_17416;
wire TIMEBOOST_net_10899;
wire g62642_sb;
wire TIMEBOOST_net_9820;
wire g62643_sb;
wire TIMEBOOST_net_6034;
wire TIMEBOOST_net_10761;
wire g62644_sb;
wire g62645_sb;
wire g62646_sb;
wire TIMEBOOST_net_22134;
wire g62647_sb;
wire TIMEBOOST_net_11030;
wire TIMEBOOST_net_5510;
wire g62648_sb;
wire TIMEBOOST_net_11000;
wire TIMEBOOST_net_13795;
wire g62649_sb;
wire TIMEBOOST_net_17427;
wire g62650_sb;
wire TIMEBOOST_net_15874;
wire g62651_sb;
wire TIMEBOOST_net_9829;
wire TIMEBOOST_net_21062;
wire g62652_sb;
wire TIMEBOOST_net_11016;
wire g62653_sb;
wire g62654_sb;
wire g62655_sb;
wire TIMEBOOST_net_10050;
wire g62656_sb;
wire TIMEBOOST_net_21784;
wire g62657_sb;
wire TIMEBOOST_net_17301;
wire g62658_sb;
wire TIMEBOOST_net_13079;
wire TIMEBOOST_net_10885;
wire g62659_sb;
wire TIMEBOOST_net_16634;
wire g62660_sb;
wire TIMEBOOST_net_21866;
wire g62661_sb;
wire TIMEBOOST_net_17303;
wire g62662_sb;
wire TIMEBOOST_net_20981;
wire g62663_sb;
wire TIMEBOOST_net_16827;
wire n_9627;
wire g62664_sb;
wire TIMEBOOST_net_22970;
wire g62665_sb;
wire TIMEBOOST_net_10162;
wire g62666_sb;
wire g62667_sb;
wire TIMEBOOST_net_12596;
wire g62668_sb;
wire TIMEBOOST_net_13078;
wire TIMEBOOST_net_17382;
wire g62669_sb;
wire TIMEBOOST_net_13077;
wire g62670_sb;
wire TIMEBOOST_net_22025;
wire g62671_sb;
wire TIMEBOOST_net_17239;
wire TIMEBOOST_net_17518;
wire g62672_sb;
wire TIMEBOOST_net_16636;
wire g62673_sb;
wire TIMEBOOST_net_13166;
wire TIMEBOOST_net_11095;
wire g62674_sb;
wire TIMEBOOST_net_10886;
wire g62675_sb;
wire TIMEBOOST_net_11096;
wire g62676_sb;
wire TIMEBOOST_net_15115;
wire TIMEBOOST_net_11018;
wire g62677_sb;
wire TIMEBOOST_net_10891;
wire g62678_sb;
wire g62679_sb;
wire TIMEBOOST_net_21901;
wire TIMEBOOST_net_11097;
wire g62680_sb;
wire TIMEBOOST_net_17552;
wire g62681_sb;
wire TIMEBOOST_net_22586;
wire g62682_sb;
wire g62683_sb;
wire TIMEBOOST_net_10804;
wire g62684_sb;
wire TIMEBOOST_net_21811;
wire TIMEBOOST_net_10809;
wire g62685_sb;
wire TIMEBOOST_net_10029;
wire TIMEBOOST_net_17328;
wire g62688_sb;
wire TIMEBOOST_net_9916;
wire TIMEBOOST_net_17474;
wire g62689_sb;
wire TIMEBOOST_net_11031;
wire TIMEBOOST_net_16932;
wire g62690_sb;
wire g62691_sb;
wire TIMEBOOST_net_13244;
wire g62693_sb;
wire TIMEBOOST_net_10027;
wire g62697_sb;
wire TIMEBOOST_net_9913;
wire TIMEBOOST_net_10887;
wire g62698_sb;
wire g62699_p;
wire TIMEBOOST_net_10025;
wire g62701_sb;
wire g62706_sb;
wire TIMEBOOST_net_22786;
wire TIMEBOOST_net_10810;
wire g62707_sb;
wire TIMEBOOST_net_16328;
wire TIMEBOOST_net_10786;
wire g62710_sb;
wire TIMEBOOST_net_14598;
wire g62711_sb;
wire TIMEBOOST_net_16333;
wire g62712_sb;
wire g62713_sb;
wire TIMEBOOST_net_23445;
wire TIMEBOOST_net_17555;
wire g62714_sb;
wire TIMEBOOST_net_12998;
wire g62715_sb;
wire TIMEBOOST_net_13522;
wire TIMEBOOST_net_14480;
wire g62716_sb;
wire TIMEBOOST_net_11039;
wire TIMEBOOST_net_22367;
wire g62719_sb;
wire TIMEBOOST_net_16666;
wire g62720_sb;
wire g62721_sb;
wire TIMEBOOST_net_13667;
wire g62722_sb;
wire g62723_sb;
wire TIMEBOOST_net_11505;
wire g62724_db;
wire TIMEBOOST_net_21345;
wire g62725_sb;
wire TIMEBOOST_net_23322;
wire g62726_sb;
wire TIMEBOOST_net_22231;
wire g62727_sb;
wire TIMEBOOST_net_22115;
wire g62728_sb;
wire TIMEBOOST_net_23169;
wire g62729_sb;
wire n_9458;
wire g62730_sb;
wire TIMEBOOST_net_16828;
wire g62731_sb;
wire TIMEBOOST_net_16829;
wire g62732_sb;
wire TIMEBOOST_net_17411;
wire TIMEBOOST_net_14852;
wire g62733_sb;
wire TIMEBOOST_net_771;
wire g62734_db;
wire g62734_sb;
wire g62735_sb;
wire TIMEBOOST_net_23435;
wire TIMEBOOST_net_16830;
wire g62736_sb;
wire n_3789;
wire g62737_sb;
wire TIMEBOOST_net_21122;
wire g62738_sb;
wire g62739_sb;
wire TIMEBOOST_net_15500;
wire g62740_sb;
wire TIMEBOOST_net_23122;
wire g62741_sb;
wire g62742_sb;
wire TIMEBOOST_net_21392;
wire g62743_sb;
wire TIMEBOOST_net_17412;
wire g62744_sb;
wire g62745_sb;
wire TIMEBOOST_net_16968;
wire g62746_sb;
wire TIMEBOOST_net_13242;
wire TIMEBOOST_net_21496;
wire g62747_sb;
wire TIMEBOOST_net_14677;
wire g62748_sb;
wire g62749_sb;
wire TIMEBOOST_net_13241;
wire TIMEBOOST_net_21506;
wire g62750_sb;
wire TIMEBOOST_net_21488;
wire g62751_sb;
wire TIMEBOOST_net_13702;
wire g62752_sb;
wire g62753_sb;
wire TIMEBOOST_net_21156;
wire TIMEBOOST_net_17582;
wire g62754_sb;
wire TIMEBOOST_net_10024;
wire g62755_sb;
wire TIMEBOOST_net_21500;
wire g62756_sb;
wire g62757_sb;
wire TIMEBOOST_net_13898;
wire TIMEBOOST_net_16637;
wire g62758_sb;
wire TIMEBOOST_net_14588;
wire g62759_sb;
wire g62760_sb;
wire g62761_sb;
wire TIMEBOOST_net_13;
wire n_9483;
wire g62762_sb;
wire TIMEBOOST_net_10023;
wire TIMEBOOST_net_11019;
wire g62763_sb;
wire g62764_sb;
wire g62765_sb;
wire TIMEBOOST_net_13438;
wire g62766_sb;
wire g62767_sb;
wire TIMEBOOST_net_21741;
wire g62768_sb;
wire g62769_sb;
wire TIMEBOOST_net_16812;
wire g62770_sb;
wire TIMEBOOST_net_15245;
wire g62771_sb;
wire TIMEBOOST_net_15246;
wire g62772_sb;
wire g62773_db;
wire g62773_sb;
wire TIMEBOOST_net_16937;
wire g62774_sb;
wire TIMEBOOST_net_23427;
wire TIMEBOOST_net_21505;
wire g62775_sb;
wire TIMEBOOST_net_21497;
wire g62776_sb;
wire TIMEBOOST_net_22200;
wire g62777_db;
wire g62777_sb;
wire TIMEBOOST_net_23147;
wire TIMEBOOST_net_21499;
wire g62778_sb;
wire TIMEBOOST_net_21826;
wire g62779_sb;
wire TIMEBOOST_net_7919;
wire g62780_sb;
wire TIMEBOOST_net_21511;
wire g62781_sb;
wire TIMEBOOST_net_16936;
wire TIMEBOOST_net_15239;
wire g62782_sb;
wire g62783_db;
wire g62783_sb;
wire TIMEBOOST_net_15240;
wire g62784_sb;
wire TIMEBOOST_net_21486;
wire g62785_sb;
wire g62786_sb;
wire TIMEBOOST_net_23131;
wire TIMEBOOST_net_15241;
wire g62787_sb;
wire TIMEBOOST_net_14254;
wire TIMEBOOST_net_15242;
wire g62788_sb;
wire TIMEBOOST_net_7604;
wire g62789_sb;
wire TIMEBOOST_net_20166;
wire TIMEBOOST_net_21503;
wire g62790_sb;
wire TIMEBOOST_net_17413;
wire g62791_sb;
wire TIMEBOOST_net_15977;
wire TIMEBOOST_net_22309;
wire g62792_sb;
wire TIMEBOOST_net_5252;
wire TIMEBOOST_net_21513;
wire g62793_sb;
wire TIMEBOOST_net_5253;
wire TIMEBOOST_net_15243;
wire g62794_sb;
wire TIMEBOOST_net_5254;
wire g62795_sb;
wire TIMEBOOST_net_5255;
wire g62796_sb;
wire TIMEBOOST_net_5256;
wire g62797_sb;
wire TIMEBOOST_net_13629;
wire TIMEBOOST_net_21492;
wire TIMEBOOST_net_22194;
wire TIMEBOOST_net_14850;
wire g62799_sb;
wire TIMEBOOST_net_5257;
wire TIMEBOOST_net_21498;
wire g62800_sb;
wire TIMEBOOST_net_5258;
wire TIMEBOOST_net_16802;
wire g62801_sb;
wire TIMEBOOST_net_5259;
wire TIMEBOOST_net_15237;
wire g62802_sb;
wire TIMEBOOST_net_17414;
wire TIMEBOOST_net_14832;
wire g62803_sb;
wire TIMEBOOST_net_21679;
wire TIMEBOOST_net_7597;
wire g62805_sb;
wire TIMEBOOST_net_5260;
wire g62806_sb;
wire TIMEBOOST_net_17084;
wire g62807_sb;
wire TIMEBOOST_net_583;
wire g62808_db;
wire g62808_sb;
wire TIMEBOOST_net_5261;
wire g62809_sb;
wire TIMEBOOST_net_5262;
wire TIMEBOOST_net_15238;
wire g62810_sb;
wire TIMEBOOST_net_14807;
wire TIMEBOOST_net_21201;
wire g62811_sb;
wire TIMEBOOST_net_5263;
wire n_9602;
wire g62812_sb;
wire TIMEBOOST_net_5264;
wire g62813_sb;
wire TIMEBOOST_net_5265;
wire TIMEBOOST_net_11001;
wire g62814_sb;
wire TIMEBOOST_net_5266;
wire TIMEBOOST_net_16864;
wire g62815_sb;
wire TIMEBOOST_net_5267;
wire g62816_sb;
wire TIMEBOOST_net_5268;
wire g62817_sb;
wire TIMEBOOST_net_5269;
wire g62818_sb;
wire TIMEBOOST_net_5270;
wire g62819_sb;
wire TIMEBOOST_net_5271;
wire g62820_sb;
wire TIMEBOOST_net_23382;
wire TIMEBOOST_net_21123;
wire g62821_sb;
wire TIMEBOOST_net_5272;
wire g62822_sb;
wire TIMEBOOST_net_5273;
wire g62823_sb;
wire TIMEBOOST_net_5274;
wire TIMEBOOST_net_15138;
wire g62824_sb;
wire TIMEBOOST_net_5275;
wire g62825_sb;
wire TIMEBOOST_net_5276;
wire g62826_sb;
wire TIMEBOOST_net_5277;
wire TIMEBOOST_net_11793;
wire g62827_sb;
wire TIMEBOOST_net_5278;
wire TIMEBOOST_net_11794;
wire g62828_sb;
wire TIMEBOOST_net_5279;
wire g62829_sb;
wire TIMEBOOST_net_5280;
wire g62830_sb;
wire TIMEBOOST_net_5281;
wire g62831_sb;
wire TIMEBOOST_net_5282;
wire g62832_sb;
wire TIMEBOOST_net_21024;
wire g62833_sb;
wire TIMEBOOST_net_5283;
wire g62834_sb;
wire TIMEBOOST_net_625;
wire g62835_db;
wire g62835_sb;
wire TIMEBOOST_net_5284;
wire g62836_sb;
wire TIMEBOOST_net_5285;
wire g62837_sb;
wire TIMEBOOST_net_5286;
wire TIMEBOOST_net_23260;
wire g62838_sb;
wire TIMEBOOST_net_5287;
wire g62839_sb;
wire TIMEBOOST_net_5288;
wire g62840_sb;
wire TIMEBOOST_net_5289;
wire g62841_sb;
wire TIMEBOOST_net_5290;
wire g62842_sb;
wire TIMEBOOST_net_17132;
wire TIMEBOOST_net_21249;
wire g62843_sb;
wire TIMEBOOST_net_16509;
wire g62844_db;
wire g62844_sb;
wire TIMEBOOST_net_5291;
wire g62845_sb;
wire TIMEBOOST_net_5292;
wire g62846_sb;
wire TIMEBOOST_net_5293;
wire g62847_sb;
wire TIMEBOOST_net_772;
wire g62848_db;
wire g62848_sb;
wire TIMEBOOST_net_5294;
wire TIMEBOOST_net_11792;
wire g62849_sb;
wire TIMEBOOST_net_5295;
wire g62850_sb;
wire TIMEBOOST_net_7600;
wire g62851_sb;
wire TIMEBOOST_net_773;
wire TIMEBOOST_net_14756;
wire g62852_sb;
wire TIMEBOOST_net_5296;
wire g62853_sb;
wire TIMEBOOST_net_5297;
wire g62854_sb;
wire TIMEBOOST_net_5298;
wire g62855_sb;
wire TIMEBOOST_net_5299;
wire TIMEBOOST_net_23191;
wire g62856_sb;
wire TIMEBOOST_net_5300;
wire g62857_sb;
wire TIMEBOOST_net_629;
wire g62858_db;
wire g62858_sb;
wire g62859_sb;
wire TIMEBOOST_net_5301;
wire g62860_sb;
wire TIMEBOOST_net_5302;
wire TIMEBOOST_net_21793;
wire g62861_sb;
wire TIMEBOOST_net_5303;
wire g62862_sb;
wire TIMEBOOST_net_5304;
wire g62863_sb;
wire TIMEBOOST_net_5305;
wire g62864_sb;
wire TIMEBOOST_net_5306;
wire g62865_sb;
wire g62873_p;
wire g62874_p;
wire g62875_p;
wire g62876_p;
wire g62877_p;
wire g62879_p;
wire g62880_p;
wire g62881_p;
wire g62882_p;
wire TIMEBOOST_net_12987;
wire g62883_sb;
wire TIMEBOOST_net_12981;
wire TIMEBOOST_net_17378;
wire g62884_sb;
wire TIMEBOOST_net_10160;
wire g62885_sb;
wire g62886_sb;
wire TIMEBOOST_net_12978;
wire g62887_sb;
wire TIMEBOOST_net_12977;
wire TIMEBOOST_net_15804;
wire g62888_sb;
wire TIMEBOOST_net_12976;
wire TIMEBOOST_net_11070;
wire g62889_sb;
wire g62890_sb;
wire TIMEBOOST_net_23452;
wire TIMEBOOST_net_17379;
wire g62891_sb;
wire TIMEBOOST_net_23450;
wire g62892_sb;
wire TIMEBOOST_net_23428;
wire TIMEBOOST_net_17533;
wire g62893_sb;
wire g62894_sb;
wire TIMEBOOST_net_13377;
wire TIMEBOOST_net_17472;
wire g62895_sb;
wire TIMEBOOST_net_13376;
wire g62896_sb;
wire TIMEBOOST_net_21717;
wire TIMEBOOST_net_17397;
wire g62897_sb;
wire TIMEBOOST_net_10159;
wire TIMEBOOST_net_16638;
wire g62898_sb;
wire TIMEBOOST_net_9884;
wire TIMEBOOST_net_11081;
wire g62899_sb;
wire TIMEBOOST_net_9883;
wire TIMEBOOST_net_11082;
wire g62900_sb;
wire TIMEBOOST_net_10158;
wire g62901_sb;
wire TIMEBOOST_net_10157;
wire g62902_sb;
wire TIMEBOOST_net_23348;
wire TIMEBOOST_net_17588;
wire g62903_sb;
wire TIMEBOOST_net_22889;
wire TIMEBOOST_net_17514;
wire g62904_sb;
wire TIMEBOOST_net_23537;
wire TIMEBOOST_net_10770;
wire g62905_sb;
wire TIMEBOOST_net_10156;
wire TIMEBOOST_net_20915;
wire g62906_sb;
wire TIMEBOOST_net_23434;
wire TIMEBOOST_net_15918;
wire g62907_sb;
wire TIMEBOOST_net_22035;
wire g62908_sb;
wire TIMEBOOST_net_10015;
wire TIMEBOOST_net_10947;
wire g62909_sb;
wire TIMEBOOST_net_13010;
wire TIMEBOOST_net_11075;
wire g62910_sb;
wire g62911_sb;
wire TIMEBOOST_net_10155;
wire TIMEBOOST_net_14624;
wire g62912_sb;
wire TIMEBOOST_net_10889;
wire g62913_sb;
wire TIMEBOOST_net_11076;
wire g62914_sb;
wire TIMEBOOST_net_22583;
wire TIMEBOOST_net_20173;
wire g62915_sb;
wire TIMEBOOST_net_12810;
wire g62916_sb;
wire TIMEBOOST_net_11079;
wire g62917_sb;
wire TIMEBOOST_net_11080;
wire g62918_sb;
wire TIMEBOOST_net_23035;
wire g62919_sb;
wire TIMEBOOST_net_23149;
wire TIMEBOOST_net_13017;
wire g62920_sb;
wire TIMEBOOST_net_17297;
wire TIMEBOOST_net_17399;
wire g62921_sb;
wire TIMEBOOST_net_11025;
wire g62922_sb;
wire TIMEBOOST_net_22096;
wire g62923_sb;
wire TIMEBOOST_net_13608;
wire TIMEBOOST_net_10772;
wire g62924_sb;
wire g62925_db;
wire g62925_sb;
wire TIMEBOOST_net_21410;
wire g62926_sb;
wire g62927_sb;
wire TIMEBOOST_net_17003;
wire g62928_sb;
wire TIMEBOOST_net_17537;
wire g62929_sb;
wire TIMEBOOST_net_20992;
wire g62930_sb;
wire TIMEBOOST_net_21175;
wire g62931_sb;
wire TIMEBOOST_net_21715;
wire TIMEBOOST_net_10774;
wire g62932_sb;
wire TIMEBOOST_net_21695;
wire TIMEBOOST_net_10775;
wire g62933_sb;
wire TIMEBOOST_net_21690;
wire g62934_sb;
wire TIMEBOOST_net_21701;
wire TIMEBOOST_net_17473;
wire g62935_sb;
wire TIMEBOOST_net_20617;
wire TIMEBOOST_net_17580;
wire g62936_sb;
wire g62937_sb;
wire TIMEBOOST_net_14634;
wire TIMEBOOST_net_10950;
wire g62938_sb;
wire g62939_sb;
wire TIMEBOOST_net_10779;
wire g62940_sb;
wire TIMEBOOST_net_10951;
wire g62941_sb;
wire TIMEBOOST_net_12811;
wire TIMEBOOST_net_10903;
wire g62942_sb;
wire TIMEBOOST_net_13855;
wire TIMEBOOST_net_10780;
wire g62943_sb;
wire TIMEBOOST_net_22365;
wire TIMEBOOST_net_10781;
wire g62944_sb;
wire TIMEBOOST_net_10222;
wire g62945_sb;
wire TIMEBOOST_net_13895;
wire TIMEBOOST_net_10782;
wire g62946_sb;
wire TIMEBOOST_net_10154;
wire TIMEBOOST_net_20905;
wire g62947_sb;
wire TIMEBOOST_net_10153;
wire g62948_sb;
wire TIMEBOOST_net_13829;
wire g62949_sb;
wire TIMEBOOST_net_14643;
wire TIMEBOOST_net_10784;
wire g62950_sb;
wire TIMEBOOST_net_9986;
wire TIMEBOOST_net_10785;
wire g62951_sb;
wire TIMEBOOST_net_21408;
wire TIMEBOOST_net_11002;
wire g62952_sb;
wire TIMEBOOST_net_14635;
wire g62953_sb;
wire TIMEBOOST_net_13902;
wire g62954_sb;
wire TIMEBOOST_net_16952;
wire TIMEBOOST_net_16530;
wire g62955_sb;
wire TIMEBOOST_net_16531;
wire g62956_sb;
wire g62957_sb;
wire TIMEBOOST_net_13905;
wire TIMEBOOST_net_10812;
wire g62958_sb;
wire TIMEBOOST_net_9983;
wire g62959_sb;
wire TIMEBOOST_net_10150;
wire TIMEBOOST_net_16532;
wire g62960_sb;
wire TIMEBOOST_net_10149;
wire TIMEBOOST_net_16533;
wire g62961_sb;
wire TIMEBOOST_net_13903;
wire TIMEBOOST_net_10814;
wire g62962_sb;
wire TIMEBOOST_net_17556;
wire TIMEBOOST_net_5511;
wire g62963_sb;
wire TIMEBOOST_net_14646;
wire TIMEBOOST_net_16754;
wire g62964_sb;
wire TIMEBOOST_net_9970;
wire TIMEBOOST_net_10815;
wire g62965_sb;
wire TIMEBOOST_net_10119;
wire g62966_sb;
wire TIMEBOOST_net_10148;
wire TIMEBOOST_net_14577;
wire g62967_sb;
wire g64783_db;
wire TIMEBOOST_net_16534;
wire g62968_sb;
wire TIMEBOOST_net_14644;
wire g62969_sb;
wire TIMEBOOST_net_12995;
wire TIMEBOOST_net_10816;
wire g62970_sb;
wire TIMEBOOST_net_17519;
wire g62971_sb;
wire TIMEBOOST_net_10817;
wire g62972_sb;
wire TIMEBOOST_net_17041;
wire TIMEBOOST_net_17530;
wire g62973_sb;
wire TIMEBOOST_net_10818;
wire g62974_sb;
wire TIMEBOOST_net_10248;
wire TIMEBOOST_net_17523;
wire g62975_sb;
wire TIMEBOOST_net_12964;
wire g62976_sb;
wire TIMEBOOST_net_17040;
wire g62977_sb;
wire g62978_sb;
wire g62979_sb;
wire g62980_sb;
wire TIMEBOOST_net_10958;
wire g62981_sb;
wire TIMEBOOST_net_10959;
wire g62982_sb;
wire TIMEBOOST_net_20435;
wire TIMEBOOST_net_16535;
wire g62983_sb;
wire TIMEBOOST_net_13831;
wire TIMEBOOST_net_10820;
wire g62984_sb;
wire TIMEBOOST_net_10237;
wire g62985_sb;
wire TIMEBOOST_net_13901;
wire g62986_sb;
wire g62987_sb;
wire TIMEBOOST_net_16536;
wire g62988_sb;
wire TIMEBOOST_net_13904;
wire g62989_sb;
wire TIMEBOOST_net_10231;
wire TIMEBOOST_net_10803;
wire g62990_sb;
wire TIMEBOOST_net_13900;
wire TIMEBOOST_net_10823;
wire g62991_sb;
wire g62992_sb;
wire TIMEBOOST_net_13893;
wire TIMEBOOST_net_10824;
wire g62993_sb;
wire TIMEBOOST_net_21158;
wire g62994_sb;
wire TIMEBOOST_net_12957;
wire g62995_sb;
wire TIMEBOOST_net_10229;
wire g62996_sb;
wire TIMEBOOST_net_23438;
wire TIMEBOOST_net_10827;
wire g62997_sb;
wire TIMEBOOST_net_14578;
wire g62998_sb;
wire TIMEBOOST_net_12975;
wire g62999_sb;
wire TIMEBOOST_net_15296;
wire g63000_sb;
wire TIMEBOOST_net_9977;
wire g63001_sb;
wire TIMEBOOST_net_9976;
wire TIMEBOOST_net_10830;
wire g63002_sb;
wire TIMEBOOST_net_22527;
wire g63003_sb;
wire TIMEBOOST_net_16945;
wire TIMEBOOST_net_14579;
wire g63004_sb;
wire TIMEBOOST_net_21031;
wire g63005_sb;
wire TIMEBOOST_net_12966;
wire TIMEBOOST_net_10831;
wire g63006_sb;
wire g63007_sb;
wire TIMEBOOST_net_14580;
wire g63008_sb;
wire TIMEBOOST_net_10220;
wire g63009_sb;
wire TIMEBOOST_net_5307;
wire g63010_sb;
wire TIMEBOOST_net_9973;
wire TIMEBOOST_net_10833;
wire g63011_sb;
wire TIMEBOOST_net_5308;
wire TIMEBOOST_net_23130;
wire g63012_sb;
wire TIMEBOOST_net_14867;
wire g63013_sb;
wire TIMEBOOST_net_5309;
wire g63014_sb;
wire TIMEBOOST_net_5310;
wire g63015_sb;
wire TIMEBOOST_net_17549;
wire TIMEBOOST_net_14759;
wire g63016_sb;
wire TIMEBOOST_net_5311;
wire g63017_sb;
wire TIMEBOOST_net_5312;
wire TIMEBOOST_net_11821;
wire g63018_sb;
wire TIMEBOOST_net_5313;
wire g63019_sb;
wire TIMEBOOST_net_758;
wire g63020_sb;
wire TIMEBOOST_net_5314;
wire g63021_sb;
wire TIMEBOOST_net_5315;
wire TIMEBOOST_net_12781;
wire g63022_sb;
wire TIMEBOOST_net_5316;
wire g63023_sb;
wire TIMEBOOST_net_16946;
wire g63024_sb;
wire TIMEBOOST_net_759;
wire TIMEBOOST_net_21124;
wire TIMEBOOST_net_23081;
wire g63026_sb;
wire TIMEBOOST_net_11492;
wire g63027_sb;
wire TIMEBOOST_net_5319;
wire g63028_sb;
wire g63029_sb;
wire TIMEBOOST_net_5320;
wire g63030_sb;
wire TIMEBOOST_net_5321;
wire g63031_sb;
wire TIMEBOOST_net_5322;
wire g63032_sb;
wire g63033_sb;
wire TIMEBOOST_net_5324;
wire TIMEBOOST_net_9576;
wire g63034_sb;
wire TIMEBOOST_net_5325;
wire g63035_sb;
wire TIMEBOOST_net_5326;
wire g63036_sb;
wire TIMEBOOST_net_5327;
wire g63037_sb;
wire TIMEBOOST_net_5328;
wire g63038_sb;
wire TIMEBOOST_net_764;
wire TIMEBOOST_net_21125;
wire g63039_sb;
wire TIMEBOOST_net_5329;
wire g63040_sb;
wire g63041_sb;
wire TIMEBOOST_net_10218;
wire g63042_sb;
wire TIMEBOOST_net_15428;
wire g63043_sb;
wire TIMEBOOST_net_5332;
wire g63044_sb;
wire TIMEBOOST_net_760;
wire TIMEBOOST_net_13631;
wire g63045_sb;
wire g63046_sb;
wire TIMEBOOST_net_761;
wire g63047_db;
wire g63047_sb;
wire TIMEBOOST_net_762;
wire g63048_sb;
wire g63049_sb;
wire g63050_sb;
wire TIMEBOOST_net_10014;
wire g63051_sb;
wire TIMEBOOST_net_763;
wire TIMEBOOST_net_20795;
wire g63052_sb;
wire TIMEBOOST_net_5337;
wire g63053_sb;
wire TIMEBOOST_net_5338;
wire TIMEBOOST_net_15653;
wire g63054_sb;
wire TIMEBOOST_net_16955;
wire g63055_sb;
wire TIMEBOOST_net_630;
wire g63056_sb;
wire TIMEBOOST_net_631;
wire TIMEBOOST_net_7599;
wire TIMEBOOST_net_632;
wire TIMEBOOST_net_14953;
wire g63058_sb;
wire g63059_sb;
wire TIMEBOOST_net_11493;
wire g63060_sb;
wire TIMEBOOST_net_21789;
wire g63061_sb;
wire TIMEBOOST_net_15485;
wire g63062_sb;
wire TIMEBOOST_net_11494;
wire g63063_db;
wire g63063_sb;
wire TIMEBOOST_net_14283;
wire g63064_sb;
wire g63065_sb;
wire TIMEBOOST_net_5345;
wire g63066_sb;
wire TIMEBOOST_net_13511;
wire g63067_sb;
wire g63068_sb;
wire TIMEBOOST_net_5348;
wire g63069_sb;
wire g63070_sb;
wire TIMEBOOST_net_23013;
wire TIMEBOOST_net_11764;
wire g63071_sb;
wire TIMEBOOST_net_5351;
wire g63072_sb;
wire TIMEBOOST_net_21633;
wire TIMEBOOST_net_21894;
wire g63073_sb;
wire TIMEBOOST_net_5353;
wire g63074_sb;
wire TIMEBOOST_net_5354;
wire g63075_sb;
wire TIMEBOOST_net_22245;
wire TIMEBOOST_net_21721;
wire g63076_sb;
wire TIMEBOOST_net_633;
wire TIMEBOOST_net_23414;
wire g63077_sb;
wire TIMEBOOST_net_5356;
wire TIMEBOOST_net_21681;
wire g63078_sb;
wire TIMEBOOST_net_5357;
wire TIMEBOOST_net_16370;
wire g63079_sb;
wire TIMEBOOST_net_16949;
wire g63080_sb;
wire TIMEBOOST_net_5359;
wire g63081_sb;
wire TIMEBOOST_net_5360;
wire g63082_sb;
wire TIMEBOOST_net_5361;
wire g63083_sb;
wire TIMEBOOST_net_14155;
wire TIMEBOOST_net_15683;
wire g63084_sb;
wire TIMEBOOST_net_634;
wire TIMEBOOST_net_23446;
wire g63085_sb;
wire TIMEBOOST_net_635;
wire g63086_db;
wire g63086_sb;
wire TIMEBOOST_net_21657;
wire g63087_sb;
wire TIMEBOOST_net_5364;
wire g63088_sb;
wire TIMEBOOST_net_636;
wire TIMEBOOST_net_14945;
wire g63089_sb;
wire TIMEBOOST_net_12031;
wire g63090_sb;
wire TIMEBOOST_net_7342;
wire g63091_sb;
wire TIMEBOOST_net_13705;
wire g63092_sb;
wire TIMEBOOST_net_5367;
wire g63093_sb;
wire TIMEBOOST_net_10834;
wire g63094_sb;
wire g63095_db;
wire g63095_sb;
wire TIMEBOOST_net_7598;
wire g63096_sb;
wire TIMEBOOST_net_20932;
wire g63097_sb;
wire TIMEBOOST_net_21780;
wire g63098_sb;
wire TIMEBOOST_net_22313;
wire g63099_sb;
wire TIMEBOOST_net_7515;
wire TIMEBOOST_net_15417;
wire g63100_sb;
wire TIMEBOOST_net_23377;
wire g63101_db;
wire g63101_sb;
wire g63102_sb;
wire TIMEBOOST_net_5373;
wire g63103_sb;
wire TIMEBOOST_net_13560;
wire g63104_sb;
wire TIMEBOOST_net_13546;
wire g63105_sb;
wire TIMEBOOST_net_5376;
wire g63106_sb;
wire g63107_sb;
wire TIMEBOOST_net_9955;
wire g63108_sb;
wire TIMEBOOST_net_5378;
wire g63109_sb;
wire TIMEBOOST_net_13565;
wire g63110_sb;
wire TIMEBOOST_net_13558;
wire g63111_sb;
wire TIMEBOOST_net_17051;
wire g63112_sb;
wire TIMEBOOST_net_14335;
wire g63113_sb;
wire g63114_sb;
wire TIMEBOOST_net_5384;
wire g63115_sb;
wire TIMEBOOST_net_13549;
wire g63116_sb;
wire TIMEBOOST_net_21771;
wire g63117_sb;
wire TIMEBOOST_net_20716;
wire g63118_sb;
wire g63119_sb;
wire TIMEBOOST_net_14739;
wire g63120_sb;
wire TIMEBOOST_net_15399;
wire g63121_sb;
wire g63122_sb;
wire g63123_sb;
wire TIMEBOOST_net_14514;
wire g63124_db;
wire g63124_sb;
wire g63125_sb;
wire TIMEBOOST_net_637;
wire g63126_db;
wire g63126_sb;
wire TIMEBOOST_net_13630;
wire g63127_db;
wire TIMEBOOST_net_5393;
wire TIMEBOOST_net_23175;
wire g63128_sb;
wire TIMEBOOST_net_638;
wire TIMEBOOST_net_7601;
wire TIMEBOOST_net_23387;
wire g63130_sb;
wire TIMEBOOST_net_12041;
wire g63131_sb;
wire g63132_sb;
wire TIMEBOOST_net_21648;
wire TIMEBOOST_net_11652;
wire g63133_sb;
wire TIMEBOOST_net_14678;
wire g63134_sb;
wire TIMEBOOST_net_15494;
wire TIMEBOOST_net_11654;
wire g63135_sb;
wire TIMEBOOST_net_15953;
wire g63136_sb;
wire TIMEBOOST_net_5401;
wire g63137_sb;
wire TIMEBOOST_net_639;
wire TIMEBOOST_net_17031;
wire g63138_sb;
wire g63139_sb;
wire TIMEBOOST_net_14927;
wire g63140_sb;
wire TIMEBOOST_net_640;
wire g63141_db;
wire g63141_sb;
wire n_9410;
wire g63142_sb;
wire n_8998;
wire g63143_sb;
wire TIMEBOOST_net_17026;
wire g63144_sb;
wire g63145_sb;
wire TIMEBOOST_net_10837;
wire g63146_sb;
wire TIMEBOOST_net_12985;
wire TIMEBOOST_net_10838;
wire g63147_sb;
wire TIMEBOOST_net_12965;
wire g63148_sb;
wire TIMEBOOST_net_14782;
wire TIMEBOOST_net_14950;
wire g63149_sb;
wire TIMEBOOST_net_13833;
wire TIMEBOOST_net_10841;
wire g63150_sb;
wire TIMEBOOST_net_20605;
wire TIMEBOOST_net_21445;
wire g63151_sb;
wire TIMEBOOST_net_14754;
wire g63152_sb;
wire TIMEBOOST_net_21434;
wire g63153_sb;
wire g63154_db;
wire g63154_sb;
wire TIMEBOOST_net_17025;
wire g63155_sb;
wire g63156_sb;
wire TIMEBOOST_net_10238;
wire TIMEBOOST_net_8852;
wire g63157_sb;
wire TIMEBOOST_net_10236;
wire TIMEBOOST_net_10847;
wire g63158_sb;
wire TIMEBOOST_net_16931;
wire TIMEBOOST_net_16537;
wire g63159_sb;
wire TIMEBOOST_net_15410;
wire TIMEBOOST_net_16538;
wire g63160_sb;
wire TIMEBOOST_net_10134;
wire TIMEBOOST_net_16539;
wire g63161_sb;
wire TIMEBOOST_net_13896;
wire g63162_sb;
wire TIMEBOOST_net_10228;
wire g63163_sb;
wire g63164_sb;
wire TIMEBOOST_net_14523;
wire g63165_sb;
wire g63166_sb;
wire TIMEBOOST_net_17024;
wire TIMEBOOST_net_10852;
wire g63167_sb;
wire TIMEBOOST_net_10205;
wire TIMEBOOST_net_10853;
wire g63168_sb;
wire TIMEBOOST_net_14821;
wire TIMEBOOST_net_23214;
wire g63169_sb;
wire g63170_sb;
wire TIMEBOOST_net_10202;
wire TIMEBOOST_net_21438;
wire g63171_sb;
wire TIMEBOOST_net_14752;
wire g63172_sb;
wire TIMEBOOST_net_13892;
wire TIMEBOOST_net_10855;
wire g63173_sb;
wire TIMEBOOST_net_22379;
wire TIMEBOOST_net_10856;
wire g63174_sb;
wire TIMEBOOST_net_5410;
wire TIMEBOOST_net_23318;
wire g63175_sb;
wire TIMEBOOST_net_14894;
wire g63176_sb;
wire g63177_sb;
wire TIMEBOOST_net_10132;
wire TIMEBOOST_net_16540;
wire g63178_sb;
wire TIMEBOOST_net_23388;
wire g63179_db;
wire g63179_sb;
wire TIMEBOOST_net_21526;
wire g63180_sb;
wire g63181_sb;
wire TIMEBOOST_net_20733;
wire TIMEBOOST_net_20452;
wire g63182_sb;
wire TIMEBOOST_net_10858;
wire g63183_sb;
wire g54314_db;
wire g63184_sb;
wire TIMEBOOST_net_13322;
wire TIMEBOOST_net_10860;
wire g63185_sb;
wire TIMEBOOST_net_17543;
wire g63186_sb;
wire TIMEBOOST_net_17018;
wire TIMEBOOST_net_10861;
wire g63187_sb;
wire TIMEBOOST_net_14802;
wire TIMEBOOST_net_16913;
wire g63188_sb;
wire TIMEBOOST_net_17016;
wire TIMEBOOST_net_10862;
wire g63189_sb;
wire TIMEBOOST_net_17015;
wire TIMEBOOST_net_10863;
wire g63190_sb;
wire TIMEBOOST_net_14823;
wire TIMEBOOST_net_23162;
wire g63191_sb;
wire TIMEBOOST_net_10864;
wire g63192_sb;
wire TIMEBOOST_net_7614;
wire TIMEBOOST_net_21583;
wire g63193_sb;
wire TIMEBOOST_net_9328;
wire g63194_sb;
wire g63195_sb;
wire TIMEBOOST_net_14834;
wire g63196_sb;
wire TIMEBOOST_net_13852;
wire g63197_sb;
wire TIMEBOOST_net_11116;
wire g63198_db;
wire g63198_sb;
wire TIMEBOOST_net_11117;
wire g63199_db;
wire g63199_sb;
wire g63200_p;
wire g63201_p;
wire TIMEBOOST_net_9945;
wire g63202_sb;
wire TIMEBOOST_net_9946;
wire g63203_sb;
wire TIMEBOOST_net_9947;
wire g63204_sb;
wire g63206_p;
wire g63207_p;
wire g63208_p;
wire g63209_p;
wire g63215_p;
wire g63216_p;
wire g63217_p;
wire g63252_p;
wire g63253_p;
wire g63256_p;
wire g63259_p;
wire g63263_p;
wire g63268_p;
wire g63271_p;
wire g63291_p;
wire g63292_p;
wire g63293_p;
wire g63307_p;
wire g63315_p;
wire g63338_p;
wire g63340_p;
wire g63348_p;
wire g63361_p;
wire g63362_p;
wire g63364_p;
wire TIMEBOOST_net_11496;
wire TIMEBOOST_net_21126;
wire g63378_sb;
wire TIMEBOOST_net_14855;
wire g63392_sb;
wire TIMEBOOST_net_20890;
wire TIMEBOOST_net_23168;
wire g63397_sb;
wire g63409_p;
wire g63422_p;
wire g63423_p;
wire g63424_p;
wire g63426_p;
wire g63428_p;
wire g63429_p;
wire g63430_p;
wire TIMEBOOST_net_5417;
wire g63431_sb;
wire TIMEBOOST_net_14709;
wire TIMEBOOST_net_21744;
wire g63432_sb;
wire TIMEBOOST_net_23151;
wire g63433_sb;
wire TIMEBOOST_net_5420;
wire TIMEBOOST_net_20454;
wire g63434_sb;
wire TIMEBOOST_net_20876;
wire g63435_sb;
wire g63436_sb;
wire TIMEBOOST_net_16916;
wire g63437_sb;
wire TIMEBOOST_net_20892;
wire g63438_sb;
wire g63525_p;
wire TIMEBOOST_net_20340;
wire g63530_sb;
wire g63533_db;
wire g63533_sb;
wire TIMEBOOST_net_16649;
wire TIMEBOOST_net_22906;
wire g63537_sb;
wire g63538_db;
wire g63538_sb;
wire g63539_p;
wire g63542_p;
wire TIMEBOOST_net_21119;
wire g63543_db;
wire g63543_sb;
wire TIMEBOOST_net_22133;
wire g63544_db;
wire g63544_sb;
wire TIMEBOOST_net_8841;
wire TIMEBOOST_net_16400;
wire g63545_sb;
wire g63546_p;
wire g63547_db;
wire g63547_sb;
wire TIMEBOOST_net_22551;
wire g63548_db;
wire g63548_sb;
wire g63549_db;
wire g63549_sb;
wire TIMEBOOST_net_14949;
wire TIMEBOOST_net_21716;
wire g63550_sb;
wire TIMEBOOST_net_14863;
wire TIMEBOOST_net_16918;
wire g63551_sb;
wire TIMEBOOST_net_14833;
wire TIMEBOOST_net_20420;
wire g63552_sb;
wire TIMEBOOST_net_21023;
wire TIMEBOOST_net_21756;
wire g63553_sb;
wire TIMEBOOST_net_20609;
wire TIMEBOOST_net_20421;
wire g63554_sb;
wire TIMEBOOST_net_14762;
wire TIMEBOOST_net_21614;
wire g63555_sb;
wire g63556_sb;
wire TIMEBOOST_net_7998;
wire TIMEBOOST_net_11740;
wire g63557_sb;
wire TIMEBOOST_net_20391;
wire g63559_sb;
wire TIMEBOOST_net_14386;
wire g63560_sb;
wire g63561_sb;
wire TIMEBOOST_net_16005;
wire g63562_sb;
wire g63563_sb;
wire g63564_sb;
wire TIMEBOOST_net_14326;
wire g63565_db;
wire g63565_sb;
wire TIMEBOOST_net_23548;
wire g63566_sb;
wire g63567_db;
wire g63567_sb;
wire g63568_db;
wire g63568_sb;
wire TIMEBOOST_net_15176;
wire TIMEBOOST_net_12035;
wire g63569_sb;
wire TIMEBOOST_net_22827;
wire g63570_db;
wire g63570_sb;
wire TIMEBOOST_net_21128;
wire g63571_sb;
wire TIMEBOOST_net_645;
wire g63572_sb;
wire TIMEBOOST_net_646;
wire g63573_sb;
wire TIMEBOOST_net_21129;
wire g63574_sb;
wire TIMEBOOST_net_10264;
wire TIMEBOOST_net_11588;
wire g63576_sb;
wire g63577_sb;
wire g63578_p;
wire g63579_p;
wire g63580_p;
wire g63581_p;
wire TIMEBOOST_net_21457;
wire g63582_db;
wire g63582_sb;
wire TIMEBOOST_net_9321;
wire TIMEBOOST_net_13962;
wire g63584_db;
wire g63584_sb;
wire g63585_db;
wire TIMEBOOST_net_338;
wire g63586_db;
wire g63586_sb;
wire TIMEBOOST_net_20657;
wire g63587_db;
wire TIMEBOOST_net_16510;
wire g63588_db;
wire g63588_sb;
wire TIMEBOOST_net_17022;
wire g63589_sb;
wire g63590_db;
wire g63590_sb;
wire TIMEBOOST_net_9487;
wire TIMEBOOST_net_562;
wire g63591_sb;
wire TIMEBOOST_net_23442;
wire g63592_sb;
wire g63593_sb;
wire TIMEBOOST_net_9488;
wire g63594_sb;
wire g65905_db;
wire g63595_sb;
wire TIMEBOOST_net_16843;
wire TIMEBOOST_net_23413;
wire g63596_sb;
wire g63597_sb;
wire TIMEBOOST_net_9489;
wire g63598_sb;
wire TIMEBOOST_net_11424;
wire g63599_db;
wire g63599_sb;
wire TIMEBOOST_net_9490;
wire TIMEBOOST_net_565;
wire g63600_sb;
wire TIMEBOOST_net_16845;
wire g63601_db;
wire g63601_sb;
wire g63602_db;
wire g63602_sb;
wire g63603_db;
wire g63603_sb;
wire TIMEBOOST_net_9491;
wire TIMEBOOST_net_566;
wire g63604_sb;
wire g63605_db;
wire g63605_sb;
wire TIMEBOOST_net_16355;
wire g63606_sb;
wire g63607_db;
wire g63607_sb;
wire TIMEBOOST_net_9492;
wire TIMEBOOST_net_13229;
wire g63608_sb;
wire g65920_db;
wire g63609_sb;
wire TIMEBOOST_net_9493;
wire TIMEBOOST_net_20749;
wire g63610_sb;
wire TIMEBOOST_net_21302;
wire g63611_db;
wire g63611_sb;
wire g63612_sb;
wire TIMEBOOST_net_476;
wire g63613_db;
wire g63613_sb;
wire TIMEBOOST_net_477;
wire g63614_db;
wire g63614_sb;
wire TIMEBOOST_net_9494;
wire TIMEBOOST_net_569;
wire g63615_sb;
wire g63616_sb;
wire TIMEBOOST_net_9495;
wire g63617_sb;
wire TIMEBOOST_net_17135;
wire g63618_db;
wire g63618_sb;
wire TIMEBOOST_net_478;
wire g63619_db;
wire g63619_sb;
wire TIMEBOOST_net_9496;
wire g63620_sb;
wire TIMEBOOST_net_9497;
wire TIMEBOOST_net_13222;
wire g63621_sb;
wire g63891_p;
wire g63892_p;
wire g63895_p;
wire g63902_p;
wire g63916_p;
wire g63922_p;
wire g63925_p;
wire g63935_p;
wire g63939_p;
wire TIMEBOOST_net_20536;
wire TIMEBOOST_net_13700;
wire g63943_p;
wire g63989_p;
wire g64022_p;
wire TIMEBOOST_net_14962;
wire g64078_db;
wire g64078_sb;
wire g64079_db;
wire g64079_sb;
wire TIMEBOOST_net_14835;
wire TIMEBOOST_net_23373;
wire g64080_sb;
wire TIMEBOOST_net_20336;
wire g64081_sb;
wire g64082_sb;
wire g64083_db;
wire g64083_sb;
wire TIMEBOOST_net_21884;
wire g64084_sb;
wire TIMEBOOST_net_14628;
wire g64085_db;
wire g64085_sb;
wire g64086_sb;
wire TIMEBOOST_net_16651;
wire TIMEBOOST_net_17053;
wire g64087_sb;
wire TIMEBOOST_net_16671;
wire g64088_sb;
wire TIMEBOOST_net_20878;
wire g64089_sb;
wire TIMEBOOST_net_14470;
wire g64090_db;
wire g64090_sb;
wire TIMEBOOST_net_16950;
wire g64091_sb;
wire TIMEBOOST_net_20611;
wire g64092_sb;
wire TIMEBOOST_net_15339;
wire TIMEBOOST_net_22561;
wire g64093_sb;
wire TIMEBOOST_net_21032;
wire g64094_sb;
wire TIMEBOOST_net_14141;
wire g64095_sb;
wire TIMEBOOST_net_14631;
wire TIMEBOOST_net_7603;
wire g64096_sb;
wire TIMEBOOST_net_8590;
wire g64097_sb;
wire TIMEBOOST_net_22053;
wire g64098_sb;
wire TIMEBOOST_net_21732;
wire TIMEBOOST_net_14639;
wire g64099_sb;
wire g64100_sb;
wire TIMEBOOST_net_9423;
wire TIMEBOOST_net_15455;
wire g64102_sb;
wire TIMEBOOST_net_14520;
wire g64103_sb;
wire TIMEBOOST_net_9413;
wire TIMEBOOST_net_14460;
wire g64105_sb;
wire TIMEBOOST_net_21667;
wire g64106_db;
wire g64106_sb;
wire TIMEBOOST_net_21686;
wire TIMEBOOST_net_12911;
wire g64107_sb;
wire g64108_sb;
wire TIMEBOOST_net_20385;
wire g64109_sb;
wire TIMEBOOST_net_21639;
wire TIMEBOOST_net_12912;
wire g64110_sb;
wire TIMEBOOST_net_21033;
wire g64111_sb;
wire TIMEBOOST_net_20615;
wire g64112_sb;
wire g64113_sb;
wire g62789_db;
wire g64114_sb;
wire TIMEBOOST_net_21461;
wire g64115_sb;
wire g64116_db;
wire g64116_sb;
wire TIMEBOOST_net_14488;
wire TIMEBOOST_net_23490;
wire g64117_sb;
wire TIMEBOOST_net_8842;
wire g64118_sb;
wire TIMEBOOST_net_9425;
wire g64119_sb;
wire TIMEBOOST_net_9424;
wire g64120_sb;
wire TIMEBOOST_net_9430;
wire TIMEBOOST_net_21723;
wire g64122_sb;
wire TIMEBOOST_net_9431;
wire TIMEBOOST_net_7606;
wire g64123_sb;
wire g64124_p;
wire TIMEBOOST_net_21034;
wire g64125_sb;
wire TIMEBOOST_net_9432;
wire TIMEBOOST_net_21570;
wire g64126_sb;
wire TIMEBOOST_net_21607;
wire g64127_sb;
wire TIMEBOOST_net_9433;
wire g64128_sb;
wire TIMEBOOST_net_8843;
wire TIMEBOOST_net_20752;
wire g64129_sb;
wire TIMEBOOST_net_8844;
wire TIMEBOOST_net_11183;
wire g64130_sb;
wire g64131_sb;
wire TIMEBOOST_net_20325;
wire g64132_sb;
wire TIMEBOOST_net_15809;
wire g64133_sb;
wire TIMEBOOST_net_22521;
wire g64134_db;
wire g64134_sb;
wire TIMEBOOST_net_9434;
wire g64135_db;
wire g64135_sb;
wire TIMEBOOST_net_14922;
wire TIMEBOOST_net_21035;
wire g64136_sb;
wire TIMEBOOST_net_21566;
wire g64137_sb;
wire TIMEBOOST_net_9435;
wire TIMEBOOST_net_22921;
wire g64138_sb;
wire g64139_db;
wire g64139_sb;
wire TIMEBOOST_net_14923;
wire g64140_sb;
wire TIMEBOOST_net_23146;
wire TIMEBOOST_net_21569;
wire g64141_sb;
wire TIMEBOOST_net_14479;
wire g64142_sb;
wire TIMEBOOST_net_13976;
wire g64143_sb;
wire TIMEBOOST_net_8846;
wire g64144_sb;
wire TIMEBOOST_net_21433;
wire g64145_sb;
wire TIMEBOOST_net_13977;
wire g64146_sb;
wire TIMEBOOST_net_22225;
wire TIMEBOOST_net_22552;
wire g64147_sb;
wire TIMEBOOST_net_9407;
wire TIMEBOOST_net_15516;
wire g64148_sb;
wire TIMEBOOST_net_14910;
wire TIMEBOOST_net_13201;
wire g64149_sb;
wire TIMEBOOST_net_13978;
wire TIMEBOOST_net_12428;
wire g64150_sb;
wire g64151_db;
wire g64151_sb;
wire g64152_sb;
wire TIMEBOOST_net_8849;
wire TIMEBOOST_net_12429;
wire g64153_sb;
wire TIMEBOOST_net_13248;
wire g64154_sb;
wire TIMEBOOST_net_14939;
wire g64155_sb;
wire TIMEBOOST_net_22423;
wire TIMEBOOST_net_20327;
wire g64156_sb;
wire TIMEBOOST_net_20364;
wire TIMEBOOST_net_22169;
wire g64157_sb;
wire TIMEBOOST_net_16432;
wire TIMEBOOST_net_12430;
wire g64158_sb;
wire TIMEBOOST_net_13243;
wire TIMEBOOST_net_21867;
wire g64159_sb;
wire TIMEBOOST_net_13072;
wire g64160_db;
wire g64160_sb;
wire TIMEBOOST_net_23439;
wire g64161_sb;
wire TIMEBOOST_net_22779;
wire TIMEBOOST_net_21890;
wire g64162_sb;
wire TIMEBOOST_net_22784;
wire g64163_sb;
wire TIMEBOOST_net_13985;
wire TIMEBOOST_net_12431;
wire g64164_sb;
wire TIMEBOOST_net_15944;
wire g64165_sb;
wire TIMEBOOST_net_13944;
wire TIMEBOOST_net_12432;
wire g64166_sb;
wire g64167_db;
wire g64167_sb;
wire TIMEBOOST_net_13945;
wire TIMEBOOST_net_22640;
wire g64168_sb;
wire TIMEBOOST_net_9408;
wire g64169_sb;
wire TIMEBOOST_net_20977;
wire g64170_sb;
wire TIMEBOOST_net_13951;
wire TIMEBOOST_net_23372;
wire g64171_sb;
wire g58434_db;
wire g64172_sb;
wire TIMEBOOST_net_21760;
wire TIMEBOOST_net_17501;
wire g64173_sb;
wire TIMEBOOST_net_13854;
wire g64175_sb;
wire TIMEBOOST_net_13791;
wire g64176_sb;
wire TIMEBOOST_net_22227;
wire TIMEBOOST_net_22485;
wire g64177_sb;
wire TIMEBOOST_net_13799;
wire g64178_sb;
wire g64179_sb;
wire TIMEBOOST_net_21905;
wire g64180_sb;
wire TIMEBOOST_net_13807;
wire n_9775;
wire g64181_sb;
wire TIMEBOOST_net_12433;
wire g64182_sb;
wire TIMEBOOST_net_22700;
wire g64183_sb;
wire TIMEBOOST_net_13804;
wire g64184_db;
wire g64184_sb;
wire TIMEBOOST_net_8877;
wire g64185_sb;
wire g64186_sb;
wire TIMEBOOST_net_21685;
wire g64187_db;
wire g64187_sb;
wire g58421_db;
wire TIMEBOOST_net_17054;
wire g64188_sb;
wire TIMEBOOST_net_9409;
wire g54207_da;
wire g64189_sb;
wire TIMEBOOST_net_9429;
wire g64190_sb;
wire TIMEBOOST_net_9410;
wire TIMEBOOST_net_16239;
wire g64191_sb;
wire TIMEBOOST_net_22580;
wire g64192_sb;
wire TIMEBOOST_net_14102;
wire g64193_sb;
wire g64194_p;
wire TIMEBOOST_net_21528;
wire g64195_sb;
wire TIMEBOOST_net_7607;
wire g64196_sb;
wire TIMEBOOST_net_9411;
wire g64197_sb;
wire TIMEBOOST_net_13828;
wire TIMEBOOST_net_21917;
wire g64198_sb;
wire g64199_db;
wire g64199_sb;
wire TIMEBOOST_net_21646;
wire g64200_db;
wire g64200_sb;
wire g58377_db;
wire g66399_db;
wire g64201_sb;
wire TIMEBOOST_net_9412;
wire g64202_sb;
wire TIMEBOOST_net_9436;
wire TIMEBOOST_net_21776;
wire g64203_sb;
wire TIMEBOOST_net_20455;
wire TIMEBOOST_net_12914;
wire g64204_sb;
wire g64205_sb;
wire TIMEBOOST_net_21609;
wire g64206_db;
wire g64206_sb;
wire TIMEBOOST_net_9330;
wire TIMEBOOST_net_7608;
wire g64207_sb;
wire TIMEBOOST_net_22059;
wire TIMEBOOST_net_22371;
wire g64208_sb;
wire TIMEBOOST_net_14493;
wire g64209_sb;
wire TIMEBOOST_net_13994;
wire g64210_sb;
wire TIMEBOOST_net_23437;
wire TIMEBOOST_net_13202;
wire g64211_sb;
wire TIMEBOOST_net_21036;
wire g64212_sb;
wire TIMEBOOST_net_21575;
wire TIMEBOOST_net_8596;
wire g64213_sb;
wire g64214_sb;
wire TIMEBOOST_net_12915;
wire g64215_sb;
wire TIMEBOOST_net_9426;
wire TIMEBOOST_net_15905;
wire g64216_sb;
wire TIMEBOOST_net_16610;
wire g64217_sb;
wire g64218_sb;
wire TIMEBOOST_net_9427;
wire TIMEBOOST_net_7609;
wire g64219_sb;
wire g64220_sb;
wire g64221_sb;
wire TIMEBOOST_net_6804;
wire g64222_sb;
wire TIMEBOOST_net_14103;
wire TIMEBOOST_net_15802;
wire g64223_sb;
wire g64224_sb;
wire TIMEBOOST_net_17134;
wire g64225_sb;
wire g64226_sb;
wire g64227_sb;
wire TIMEBOOST_net_15398;
wire TIMEBOOST_net_17491;
wire g64228_sb;
wire g64229_sb;
wire g64230_sb;
wire TIMEBOOST_net_503;
wire TIMEBOOST_net_13876;
wire g64231_sb;
wire g64232_sb;
wire TIMEBOOST_net_22027;
wire g64233_sb;
wire g64234_sb;
wire TIMEBOOST_net_22193;
wire TIMEBOOST_net_23551;
wire g64235_sb;
wire TIMEBOOST_net_21341;
wire TIMEBOOST_net_21562;
wire g64236_sb;
wire TIMEBOOST_net_21745;
wire g64237_db;
wire g64237_sb;
wire TIMEBOOST_net_21611;
wire TIMEBOOST_net_675;
wire g64238_sb;
wire TIMEBOOST_net_16496;
wire TIMEBOOST_net_23552;
wire g64239_sb;
wire TIMEBOOST_net_17492;
wire g64240_sb;
wire TIMEBOOST_net_17344;
wire TIMEBOOST_net_20220;
wire g64241_sb;
wire TIMEBOOST_net_8209;
wire g64242_db;
wire g64242_sb;
wire TIMEBOOST_net_13696;
wire g64243_sb;
wire g64244_db;
wire g64244_sb;
wire TIMEBOOST_net_14069;
wire TIMEBOOST_net_17493;
wire g64245_sb;
wire TIMEBOOST_net_21430;
wire TIMEBOOST_net_22029;
wire g64246_sb;
wire TIMEBOOST_net_16497;
wire g64247_sb;
wire TIMEBOOST_net_22043;
wire g64248_sb;
wire TIMEBOOST_net_17033;
wire g64250_db;
wire g64250_sb;
wire TIMEBOOST_net_21725;
wire g64251_sb;
wire TIMEBOOST_net_8201;
wire g64252_db;
wire g64252_sb;
wire TIMEBOOST_net_21431;
wire TIMEBOOST_net_22918;
wire g64253_sb;
wire TIMEBOOST_net_22369;
wire TIMEBOOST_net_15565;
wire g64254_sb;
wire g64255_sb;
wire TIMEBOOST_net_21757;
wire TIMEBOOST_net_23417;
wire g64256_sb;
wire TIMEBOOST_net_16477;
wire g64257_sb;
wire TIMEBOOST_net_13931;
wire TIMEBOOST_net_17539;
wire g64258_sb;
wire TIMEBOOST_net_8199;
wire g64259_sb;
wire g64260_sb;
wire TIMEBOOST_net_8197;
wire g64261_db;
wire g64261_sb;
wire g64262_sb;
wire TIMEBOOST_net_21563;
wire g64263_sb;
wire TIMEBOOST_net_8194;
wire TIMEBOOST_net_22019;
wire g64264_sb;
wire TIMEBOOST_net_22055;
wire g64265_sb;
wire TIMEBOOST_net_21224;
wire g64266_sb;
wire TIMEBOOST_net_21347;
wire TIMEBOOST_net_17540;
wire g64267_sb;
wire TIMEBOOST_net_8679;
wire TIMEBOOST_net_20355;
wire g64268_sb;
wire TIMEBOOST_net_23444;
wire g64269_sb;
wire TIMEBOOST_net_22098;
wire TIMEBOOST_net_12436;
wire g64270_sb;
wire TIMEBOOST_net_8754;
wire g64271_sb;
wire TIMEBOOST_net_13932;
wire g64272_sb;
wire g64273_db;
wire g64273_sb;
wire g64274_sb;
wire TIMEBOOST_net_16413;
wire TIMEBOOST_net_12437;
wire g64275_sb;
wire TIMEBOOST_net_21624;
wire g64276_db;
wire g64276_sb;
wire g64277_da;
wire g64277_db;
wire g64277_sb;
wire TIMEBOOST_net_21895;
wire g64278_sb;
wire g64279_sb;
wire TIMEBOOST_net_15523;
wire g64280_db;
wire g64280_sb;
wire TIMEBOOST_net_13887;
wire TIMEBOOST_net_15100;
wire g64281_sb;
wire TIMEBOOST_net_20373;
wire g64282_sb;
wire TIMEBOOST_net_21252;
wire g64283_db;
wire g64283_sb;
wire TIMEBOOST_net_21560;
wire TIMEBOOST_net_21856;
wire g64284_sb;
wire TIMEBOOST_net_22984;
wire g64285_sb;
wire TIMEBOOST_net_21749;
wire TIMEBOOST_net_23535;
wire g64286_sb;
wire TIMEBOOST_net_23539;
wire g64287_sb;
wire TIMEBOOST_net_22117;
wire g64288_db;
wire g64288_sb;
wire TIMEBOOST_net_23534;
wire g64289_sb;
wire TIMEBOOST_net_21637;
wire g64290_sb;
wire g64291_sb;
wire g64292_sb;
wire g64293_sb;
wire TIMEBOOST_net_153;
wire g64295_sb;
wire TIMEBOOST_net_14178;
wire TIMEBOOST_net_12280;
wire g64296_sb;
wire g64297_sb;
wire TIMEBOOST_net_21777;
wire g64298_sb;
wire TIMEBOOST_net_20993;
wire g64300_sb;
wire TIMEBOOST_net_21663;
wire TIMEBOOST_net_12439;
wire g64301_sb;
wire TIMEBOOST_net_11893;
wire g64302_db;
wire g64302_sb;
wire TIMEBOOST_net_154;
wire TIMEBOOST_net_12034;
wire TIMEBOOST_net_16948;
wire g64304_sb;
wire TIMEBOOST_net_21863;
wire TIMEBOOST_net_17281;
wire g64306_sb;
wire TIMEBOOST_net_21255;
wire g64307_sb;
wire TIMEBOOST_net_21082;
wire g64308_sb;
wire TIMEBOOST_net_13933;
wire TIMEBOOST_net_17334;
wire g64309_sb;
wire TIMEBOOST_net_16498;
wire TIMEBOOST_net_23553;
wire g64310_sb;
wire TIMEBOOST_net_22093;
wire g64311_sb;
wire g64312_db;
wire g64312_sb;
wire TIMEBOOST_net_15166;
wire TIMEBOOST_net_12945;
wire g64313_sb;
wire TIMEBOOST_net_22185;
wire g64314_sb;
wire TIMEBOOST_net_9332;
wire TIMEBOOST_net_21750;
wire g64315_sb;
wire TIMEBOOST_net_15212;
wire g64316_sb;
wire g64317_sb;
wire TIMEBOOST_net_13934;
wire g64318_sb;
wire g64319_sb;
wire TIMEBOOST_net_16808;
wire g64320_sb;
wire TIMEBOOST_net_16807;
wire g64321_sb;
wire TIMEBOOST_net_15113;
wire TIMEBOOST_net_23555;
wire g64322_sb;
wire TIMEBOOST_net_15136;
wire g64323_sb;
wire TIMEBOOST_net_22625;
wire g64324_sb;
wire TIMEBOOST_net_21321;
wire g64325_sb;
wire TIMEBOOST_net_22105;
wire g64326_sb;
wire TIMEBOOST_net_17196;
wire g64327_sb;
wire TIMEBOOST_net_22815;
wire g64328_db;
wire g64328_sb;
wire g64329_sb;
wire TIMEBOOST_net_13777;
wire g64330_db;
wire g64330_sb;
wire TIMEBOOST_net_13778;
wire TIMEBOOST_net_21704;
wire g64331_sb;
wire g64332_sb;
wire TIMEBOOST_net_13779;
wire g64333_sb;
wire TIMEBOOST_net_22376;
wire TIMEBOOST_net_21980;
wire g64334_sb;
wire TIMEBOOST_net_15571;
wire g64335_sb;
wire TIMEBOOST_net_13780;
wire TIMEBOOST_net_17197;
wire g64336_sb;
wire TIMEBOOST_net_8191;
wire g64337_db;
wire g64337_sb;
wire TIMEBOOST_net_8190;
wire TIMEBOOST_net_17494;
wire g64339_sb;
wire TIMEBOOST_net_13781;
wire g64340_sb;
wire TIMEBOOST_net_16788;
wire TIMEBOOST_net_23419;
wire g64341_sb;
wire TIMEBOOST_net_21676;
wire TIMEBOOST_net_22046;
wire g64342_sb;
wire g64343_sb;
wire TIMEBOOST_net_13247;
wire g64344_sb;
wire TIMEBOOST_net_16781;
wire g64345_sb;
wire g64346_sb;
wire TIMEBOOST_net_17495;
wire g64347_sb;
wire TIMEBOOST_net_17198;
wire g64348_sb;
wire g64349_db;
wire g64349_sb;
wire TIMEBOOST_net_16453;
wire TIMEBOOST_net_17282;
wire g64350_sb;
wire TIMEBOOST_net_14864;
wire g64351_sb;
wire g64352_db;
wire g64352_sb;
wire TIMEBOOST_net_21413;
wire TIMEBOOST_net_15573;
wire g64353_sb;
wire TIMEBOOST_net_13939;
wire g64354_db;
wire g64354_sb;
wire TIMEBOOST_net_9368;
wire TIMEBOOST_net_22448;
wire g64355_sb;
wire TIMEBOOST_net_15574;
wire g64356_sb;
wire TIMEBOOST_net_13940;
wire TIMEBOOST_net_22730;
wire g64357_sb;
wire TIMEBOOST_net_13941;
wire g64358_db;
wire g64358_sb;
wire g54203_db;
wire TIMEBOOST_net_12281;
wire g64359_sb;
wire TIMEBOOST_net_17200;
wire g64360_sb;
wire TIMEBOOST_net_16501;
wire TIMEBOOST_net_17201;
wire g64361_sb;
wire TIMEBOOST_net_13942;
wire TIMEBOOST_net_17202;
wire g64362_sb;
wire TIMEBOOST_net_13943;
wire TIMEBOOST_net_17203;
wire g64363_sb;
wire TIMEBOOST_net_17366;
wire TIMEBOOST_net_7533;
wire TIMEBOOST_net_21422;
wire g64366_sb;
wire TIMEBOOST_net_13927;
wire TIMEBOOST_net_15575;
wire g64367_sb;
wire g64368_p;
wire g64369_p;
wire g64370_p;
wire g64371_p;
wire g64375_p;
wire g64376_p;
wire g64377_p;
wire g64378_p;
wire g64379_p;
wire g64380_p;
wire TIMEBOOST_net_17007;
wire g64382_p;
wire g64383_p;
wire g64384_p;
wire g64385_p;
wire g64454_p;
wire g64461_p;
wire g64465_p;
wire g64466_p;
wire g64577_p;
wire g64578_p;
wire g64581_p;
wire g64582_p;
wire g64585_p;
wire g64587_p;
wire g64595_p;
wire g64596_p;
wire g64597_p;
wire g64610_p;
wire TIMEBOOST_net_686;
wire g64630_p;
wire g64631_p;
wire g64632_p;
wire g64633_p;
wire g64639_p;
wire g64643_p;
wire g64646_p;
wire g64671_p;
wire g64678_p;
wire g64687_p;
wire g64694_p;
wire g64697_p;
wire g64700_p;
wire g64701_p;
wire g64702_p;
wire g64704_p;
wire g64705_p;
wire g64707_p;
wire g64712_p;
wire g64727_p;
wire g64736_p;
wire g64740_p;
wire g64746_p;
wire g64747_p;
wire TIMEBOOST_net_14633;
wire g64748_sb;
wire TIMEBOOST_net_12282;
wire g64749_sb;
wire g64750_sb;
wire TIMEBOOST_net_21620;
wire TIMEBOOST_net_20714;
wire g64751_sb;
wire TIMEBOOST_net_14080;
wire g64752_db;
wire g64752_sb;
wire TIMEBOOST_net_13234;
wire TIMEBOOST_net_12392;
wire g64753_sb;
wire TIMEBOOST_net_9373;
wire g64754_sb;
wire TIMEBOOST_net_9369;
wire TIMEBOOST_net_14650;
wire g64755_sb;
wire TIMEBOOST_net_17564;
wire TIMEBOOST_net_12393;
wire g64756_sb;
wire TIMEBOOST_net_22016;
wire TIMEBOOST_net_22034;
wire g64757_sb;
wire TIMEBOOST_net_16526;
wire g64758_db;
wire g64758_sb;
wire TIMEBOOST_net_9374;
wire g64759_sb;
wire g64760_sb;
wire TIMEBOOST_net_228;
wire TIMEBOOST_net_7657;
wire g64761_sb;
wire TIMEBOOST_net_13865;
wire TIMEBOOST_net_21927;
wire g64762_sb;
wire TIMEBOOST_net_15374;
wire g64763_sb;
wire TIMEBOOST_net_13857;
wire g64764_sb;
wire TIMEBOOST_net_13861;
wire g64765_sb;
wire TIMEBOOST_net_17565;
wire TIMEBOOST_net_17584;
wire g64766_sb;
wire TIMEBOOST_net_16655;
wire TIMEBOOST_net_20719;
wire g64767_sb;
wire TIMEBOOST_net_13869;
wire g64768_sb;
wire TIMEBOOST_net_9375;
wire TIMEBOOST_net_22710;
wire g64769_sb;
wire g64770_sb;
wire TIMEBOOST_net_9370;
wire g64771_sb;
wire TIMEBOOST_net_9376;
wire g64772_sb;
wire TIMEBOOST_net_185;
wire TIMEBOOST_net_13573;
wire g64773_sb;
wire g58354_da;
wire g64774_db;
wire g64774_sb;
wire TIMEBOOST_net_9371;
wire g64775_db;
wire g64775_sb;
wire TIMEBOOST_net_9377;
wire g64776_db;
wire g64776_sb;
wire TIMEBOOST_net_17566;
wire TIMEBOOST_net_12497;
wire g64777_sb;
wire TIMEBOOST_net_9372;
wire n_15731;
wire g64778_sb;
wire TIMEBOOST_net_9360;
wire TIMEBOOST_net_7660;
wire g64779_sb;
wire TIMEBOOST_net_13018;
wire g64780_db;
wire g64780_sb;
wire TIMEBOOST_net_9378;
wire g64781_db;
wire g64781_sb;
wire TIMEBOOST_net_9379;
wire g64782_sb;
wire TIMEBOOST_net_9380;
wire TIMEBOOST_net_10147;
wire g64783_sb;
wire g64784_sb;
wire TIMEBOOST_net_9381;
wire g64785_sb;
wire g64786_db;
wire g64786_sb;
wire TIMEBOOST_net_22076;
wire g64787_sb;
wire TIMEBOOST_net_16591;
wire g64788_sb;
wire TIMEBOOST_net_13982;
wire g64789_sb;
wire TIMEBOOST_net_22422;
wire g64790_sb;
wire TIMEBOOST_net_12968;
wire g64791_sb;
wire g64792_sb;
wire TIMEBOOST_net_16506;
wire g64793_sb;
wire g61840_db;
wire TIMEBOOST_net_22497;
wire g64794_sb;
wire TIMEBOOST_net_16507;
wire g64795_db;
wire g64795_sb;
wire TIMEBOOST_net_17568;
wire g64796_sb;
wire TIMEBOOST_net_20743;
wire TIMEBOOST_net_7661;
wire g64797_sb;
wire TIMEBOOST_net_12969;
wire g64798_sb;
wire TIMEBOOST_net_14499;
wire TIMEBOOST_net_17114;
wire g64799_sb;
wire TIMEBOOST_net_14025;
wire g64800_sb;
wire g64801_db;
wire g64801_sb;
wire TIMEBOOST_net_16612;
wire g64802_sb;
wire TIMEBOOST_net_17226;
wire g64803_db;
wire g64803_sb;
wire TIMEBOOST_net_9483;
wire TIMEBOOST_net_9482;
wire g64804_sb;
wire TIMEBOOST_net_14872;
wire g64805_sb;
wire TIMEBOOST_net_9382;
wire TIMEBOOST_net_15529;
wire g64806_sb;
wire TIMEBOOST_net_8838;
wire TIMEBOOST_net_13785;
wire g64807_sb;
wire TIMEBOOST_net_14478;
wire TIMEBOOST_net_15270;
wire g64808_sb;
wire g64809_sb;
wire g64810_db;
wire g64810_sb;
wire TIMEBOOST_net_22758;
wire g64811_sb;
wire TIMEBOOST_net_13988;
wire TIMEBOOST_net_12283;
wire g64812_sb;
wire TIMEBOOST_net_142;
wire g64813_sb;
wire TIMEBOOST_net_186;
wire g64814_db;
wire g64814_sb;
wire TIMEBOOST_net_264;
wire g64815_db;
wire g64815_sb;
wire TIMEBOOST_net_9361;
wire g64816_db;
wire g64816_sb;
wire TIMEBOOST_net_22626;
wire TIMEBOOST_net_20225;
wire g64817_sb;
wire TIMEBOOST_net_23527;
wire TIMEBOOST_net_15869;
wire g64818_sb;
wire TIMEBOOST_net_20610;
wire g64819_db;
wire g64819_sb;
wire n_4354;
wire TIMEBOOST_net_12285;
wire g64820_sb;
wire TIMEBOOST_net_265;
wire TIMEBOOST_net_10454;
wire g64821_sb;
wire TIMEBOOST_net_8781;
wire g64822_db;
wire g64822_sb;
wire TIMEBOOST_net_15577;
wire g64823_sb;
wire TIMEBOOST_net_16487;
wire TIMEBOOST_net_12286;
wire g64824_sb;
wire TIMEBOOST_net_14075;
wire TIMEBOOST_net_12287;
wire g64825_sb;
wire g64826_sb;
wire TIMEBOOST_net_17475;
wire g64827_sb;
wire TIMEBOOST_net_17091;
wire g64828_sb;
wire TIMEBOOST_net_20269;
wire g64829_sb;
wire TIMEBOOST_net_21382;
wire g64830_sb;
wire g64831_sb;
wire TIMEBOOST_net_17476;
wire g64832_sb;
wire TIMEBOOST_net_14485;
wire g64833_db;
wire g64833_sb;
wire TIMEBOOST_net_21820;
wire g64834_sb;
wire g64835_db;
wire g64835_sb;
wire TIMEBOOST_net_23529;
wire g64836_sb;
wire TIMEBOOST_net_17570;
wire g64837_sb;
wire TIMEBOOST_net_16343;
wire g64838_sb;
wire g64323_db;
wire g64839_sb;
wire TIMEBOOST_net_12144;
wire g64840_sb;
wire TIMEBOOST_net_9474;
wire g64841_sb;
wire TIMEBOOST_net_219;
wire TIMEBOOST_net_12288;
wire g64842_sb;
wire TIMEBOOST_net_14093;
wire g64843_db;
wire g64843_sb;
wire TIMEBOOST_net_17571;
wire TIMEBOOST_net_17204;
wire g64844_sb;
wire TIMEBOOST_net_5383;
wire g64845_sb;
wire TIMEBOOST_net_23486;
wire TIMEBOOST_net_15863;
wire g64846_sb;
wire TIMEBOOST_net_13906;
wire g64847_sb;
wire TIMEBOOST_net_13980;
wire TIMEBOOST_net_12292;
wire g64848_sb;
wire TIMEBOOST_net_22724;
wire g64849_db;
wire g64849_sb;
wire TIMEBOOST_net_12916;
wire g64850_sb;
wire TIMEBOOST_net_17572;
wire TIMEBOOST_net_12293;
wire g64851_sb;
wire TIMEBOOST_net_8275;
wire g64852_sb;
wire TIMEBOOST_net_20741;
wire TIMEBOOST_net_12294;
wire g64853_sb;
wire TIMEBOOST_net_21371;
wire TIMEBOOST_net_12295;
wire g64854_sb;
wire TIMEBOOST_net_21547;
wire g64855_sb;
wire TIMEBOOST_net_13969;
wire g64856_sb;
wire TIMEBOOST_net_14096;
wire TIMEBOOST_net_12296;
wire g64857_sb;
wire g64858_sb;
wire TIMEBOOST_net_14611;
wire TIMEBOOST_net_12458;
wire g64859_sb;
wire TIMEBOOST_net_22063;
wire g64860_sb;
wire TIMEBOOST_net_22012;
wire g64861_sb;
wire TIMEBOOST_net_14091;
wire TIMEBOOST_net_17262;
wire g64862_sb;
wire TIMEBOOST_net_13965;
wire TIMEBOOST_net_10773;
wire g64863_sb;
wire TIMEBOOST_net_21764;
wire g64864_db;
wire g64864_sb;
wire TIMEBOOST_net_12401;
wire g64865_sb;
wire TIMEBOOST_net_21909;
wire TIMEBOOST_net_23231;
wire g64866_sb;
wire TIMEBOOST_net_15684;
wire g64867_sb;
wire TIMEBOOST_net_13853;
wire TIMEBOOST_net_12402;
wire g64868_sb;
wire TIMEBOOST_net_21782;
wire TIMEBOOST_net_13050;
wire g64869_sb;
wire TIMEBOOST_net_21692;
wire TIMEBOOST_net_23510;
wire g64870_sb;
wire TIMEBOOST_net_14831;
wire g64871_sb;
wire TIMEBOOST_net_22107;
wire g64872_sb;
wire TIMEBOOST_net_535;
wire TIMEBOOST_net_14859;
wire g64873_sb;
wire TIMEBOOST_net_22781;
wire g64874_db;
wire g64874_sb;
wire TIMEBOOST_net_22535;
wire TIMEBOOST_net_17115;
wire g64875_sb;
wire TIMEBOOST_net_23451;
wire TIMEBOOST_net_14948;
wire g64876_sb;
wire TIMEBOOST_net_13975;
wire g52471_da;
wire g64877_sb;
wire TIMEBOOST_net_13291;
wire g64878_sb;
wire TIMEBOOST_net_14095;
wire TIMEBOOST_net_12297;
wire g64879_sb;
wire TIMEBOOST_net_22543;
wire TIMEBOOST_net_12298;
wire g64880_sb;
wire TIMEBOOST_net_13753;
wire TIMEBOOST_net_17206;
wire g64881_sb;
wire TIMEBOOST_net_16345;
wire TIMEBOOST_net_12299;
wire g64882_sb;
wire TIMEBOOST_net_13937;
wire g64883_sb;
wire TIMEBOOST_net_14094;
wire TIMEBOOST_net_12301;
wire g64884_sb;
wire TIMEBOOST_net_22167;
wire TIMEBOOST_net_12302;
wire g64885_sb;
wire TIMEBOOST_net_17577;
wire g64886_sb;
wire TIMEBOOST_net_14101;
wire TIMEBOOST_net_22455;
wire g64887_sb;
wire g64253_da;
wire g64888_db;
wire g64888_sb;
wire TIMEBOOST_net_8799;
wire g64889_sb;
wire TIMEBOOST_net_12304;
wire g64890_sb;
wire TIMEBOOST_net_22569;
wire TIMEBOOST_net_12305;
wire g64891_sb;
wire TIMEBOOST_net_14099;
wire TIMEBOOST_net_22077;
wire g64892_sb;
wire TIMEBOOST_net_13717;
wire TIMEBOOST_net_17208;
wire g64893_sb;
wire TIMEBOOST_net_12306;
wire g64894_sb;
wire TIMEBOOST_net_12307;
wire g64895_sb;
wire TIMEBOOST_net_21590;
wire g64896_db;
wire g64896_sb;
wire g63569_da;
wire g64897_sb;
wire g64898_sb;
wire TIMEBOOST_net_14504;
wire TIMEBOOST_net_12145;
wire g64899_sb;
wire TIMEBOOST_net_20360;
wire TIMEBOOST_net_16458;
wire g64900_sb;
wire TIMEBOOST_net_16335;
wire g64901_db;
wire g64901_sb;
wire TIMEBOOST_net_13990;
wire g64902_sb;
wire TIMEBOOST_net_14503;
wire g64903_db;
wire g64903_sb;
wire TIMEBOOST_net_22244;
wire g64904_sb;
wire TIMEBOOST_net_10448;
wire g64905_sb;
wire TIMEBOOST_net_14506;
wire g64906_sb;
wire TIMEBOOST_net_14507;
wire g64907_db;
wire g64907_sb;
wire TIMEBOOST_net_23533;
wire g64908_sb;
wire TIMEBOOST_net_13178;
wire g64909_db;
wire g64909_sb;
wire TIMEBOOST_net_21436;
wire g64910_sb;
wire g64911_sb;
wire TIMEBOOST_net_8276;
wire g64912_sb;
wire TIMEBOOST_net_21440;
wire g64913_sb;
wire TIMEBOOST_net_14032;
wire g64914_sb;
wire TIMEBOOST_net_14508;
wire g64915_sb;
wire g64916_sb;
wire TIMEBOOST_net_13798;
wire TIMEBOOST_net_23238;
wire g64917_sb;
wire TIMEBOOST_net_9122;
wire TIMEBOOST_net_12309;
wire g64918_sb;
wire TIMEBOOST_net_21731;
wire TIMEBOOST_net_12821;
wire g64919_sb;
wire TIMEBOOST_net_15163;
wire TIMEBOOST_net_323;
wire g64920_sb;
wire g64921_sb;
wire TIMEBOOST_net_14033;
wire g64922_sb;
wire TIMEBOOST_net_17290;
wire TIMEBOOST_net_15699;
wire g64923_sb;
wire g64924_sb;
wire TIMEBOOST_net_22562;
wire g64925_sb;
wire g64926_db;
wire g64926_sb;
wire g64927_sb;
wire TIMEBOOST_net_12314;
wire g64928_sb;
wire TIMEBOOST_net_21117;
wire g64929_db;
wire g64929_sb;
wire g64930_sb;
wire TIMEBOOST_net_14035;
wire TIMEBOOST_net_17287;
wire g64931_sb;
wire TIMEBOOST_net_14036;
wire g64932_db;
wire g64932_sb;
wire TIMEBOOST_net_14037;
wire g64933_db;
wire g64933_sb;
wire TIMEBOOST_net_16611;
wire g64934_sb;
wire g64935_sb;
wire TIMEBOOST_net_9127;
wire g64936_sb;
wire TIMEBOOST_net_16423;
wire TIMEBOOST_net_12319;
wire g64937_sb;
wire TIMEBOOST_net_9128;
wire TIMEBOOST_net_6769;
wire g64938_sb;
wire g64939_db;
wire g64939_sb;
wire g64940_sb;
wire TIMEBOOST_net_12854;
wire TIMEBOOST_net_17345;
wire g64941_sb;
wire TIMEBOOST_net_12853;
wire TIMEBOOST_net_17346;
wire g64942_sb;
wire TIMEBOOST_net_22044;
wire g64943_sb;
wire TIMEBOOST_net_20448;
wire g64944_sb;
wire TIMEBOOST_net_14303;
wire g64945_db;
wire g64945_sb;
wire TIMEBOOST_net_22006;
wire TIMEBOOST_net_12559;
wire g64946_sb;
wire g64947_db;
wire g64947_sb;
wire TIMEBOOST_net_22036;
wire TIMEBOOST_net_20449;
wire g64948_sb;
wire TIMEBOOST_net_20669;
wire g64949_sb;
wire g64950_db;
wire g64950_sb;
wire g64951_sb;
wire TIMEBOOST_net_20440;
wire g64952_db;
wire g64952_sb;
wire TIMEBOOST_net_9362;
wire g64953_sb;
wire TIMEBOOST_net_20170;
wire g64954_sb;
wire g64955_sb;
wire TIMEBOOST_net_12872;
wire TIMEBOOST_net_22420;
wire g64956_sb;
wire TIMEBOOST_net_12871;
wire TIMEBOOST_net_17218;
wire g64957_sb;
wire TIMEBOOST_net_12870;
wire g64958_sb;
wire TIMEBOOST_net_12404;
wire g64959_sb;
wire TIMEBOOST_net_13805;
wire g64960_sb;
wire TIMEBOOST_net_13802;
wire g64961_sb;
wire TIMEBOOST_net_22747;
wire g64962_db;
wire g64962_sb;
wire TIMEBOOST_net_8878;
wire TIMEBOOST_net_23232;
wire g64963_sb;
wire TIMEBOOST_net_13155;
wire TIMEBOOST_net_12320;
wire TIMEBOOST_net_21565;
wire g64965_sb;
wire g64966_db;
wire g64966_sb;
wire TIMEBOOST_net_13859;
wire g64967_sb;
wire TIMEBOOST_net_8839;
wire TIMEBOOST_net_21483;
wire g64968_sb;
wire TIMEBOOST_net_13858;
wire TIMEBOOST_net_12407;
wire g64969_sb;
wire TIMEBOOST_net_21274;
wire TIMEBOOST_net_17116;
wire g64970_sb;
wire TIMEBOOST_net_13860;
wire TIMEBOOST_net_12408;
wire g64971_sb;
wire TIMEBOOST_net_13051;
wire g64972_sb;
wire TIMEBOOST_net_21640;
wire g64973_db;
wire g64973_sb;
wire TIMEBOOST_net_12869;
wire TIMEBOOST_net_20282;
wire g64974_sb;
wire g64975_sb;
wire TIMEBOOST_net_13081;
wire TIMEBOOST_net_12409;
wire g64976_sb;
wire g64977_db;
wire g64977_sb;
wire TIMEBOOST_net_22567;
wire g64978_sb;
wire TIMEBOOST_net_13864;
wire TIMEBOOST_net_12410;
wire g64979_sb;
wire TIMEBOOST_net_16486;
wire TIMEBOOST_net_20226;
wire g64980_sb;
wire TIMEBOOST_net_14106;
wire TIMEBOOST_net_14078;
wire TIMEBOOST_net_22493;
wire g64982_sb;
wire TIMEBOOST_net_12868;
wire g64983_db;
wire g64983_sb;
wire TIMEBOOST_net_12867;
wire TIMEBOOST_net_10843;
wire g64984_sb;
wire g64985_sb;
wire g64986_db;
wire g64986_sb;
wire TIMEBOOST_net_15316;
wire g64987_sb;
wire TIMEBOOST_net_14306;
wire TIMEBOOST_net_20451;
wire g64988_sb;
wire TIMEBOOST_net_14016;
wire g64989_sb;
wire TIMEBOOST_net_21186;
wire TIMEBOOST_net_17213;
wire g64990_sb;
wire TIMEBOOST_net_12918;
wire g64991_sb;
wire TIMEBOOST_net_13237;
wire g64992_sb;
wire TIMEBOOST_net_16488;
wire g64993_sb;
wire TIMEBOOST_net_12324;
wire g64994_sb;
wire TIMEBOOST_net_22491;
wire g64995_db;
wire g64995_sb;
wire TIMEBOOST_net_14053;
wire TIMEBOOST_net_17214;
wire g64996_sb;
wire TIMEBOOST_net_13872;
wire g64997_sb;
wire TIMEBOOST_net_14347;
wire g64998_db;
wire g64998_sb;
wire TIMEBOOST_net_22869;
wire g64999_sb;
wire TIMEBOOST_net_16963;
wire g65000_sb;
wire TIMEBOOST_net_21846;
wire TIMEBOOST_net_12326;
wire g65001_sb;
wire g65002_db;
wire g65002_sb;
wire TIMEBOOST_net_13871;
wire g65003_db;
wire g65003_sb;
wire n_3894;
wire g65004_db;
wire g65004_sb;
wire TIMEBOOST_net_22466;
wire g65005_sb;
wire TIMEBOOST_net_23473;
wire TIMEBOOST_net_12327;
wire g65006_sb;
wire TIMEBOOST_net_13022;
wire TIMEBOOST_net_12328;
wire g65007_sb;
wire TIMEBOOST_net_12329;
wire g65008_sb;
wire TIMEBOOST_net_16482;
wire TIMEBOOST_net_22741;
wire g65009_sb;
wire TIMEBOOST_net_20376;
wire TIMEBOOST_net_7672;
wire g65010_sb;
wire TIMEBOOST_net_9383;
wire g65011_sb;
wire TIMEBOOST_net_23456;
wire TIMEBOOST_net_22860;
wire g65012_sb;
wire TIMEBOOST_net_21654;
wire TIMEBOOST_net_15404;
wire g65013_sb;
wire g65014_sb;
wire TIMEBOOST_net_17502;
wire g65015_sb;
wire g65016_sb;
wire TIMEBOOST_net_14319;
wire g65017_sb;
wire TIMEBOOST_net_20213;
wire TIMEBOOST_net_12330;
wire g65018_sb;
wire g65019_da;
wire g65019_db;
wire g65019_sb;
wire g65020_sb;
wire TIMEBOOST_net_14502;
wire g65021_sb;
wire g65022_sb;
wire TIMEBOOST_net_21391;
wire g65023_sb;
wire TIMEBOOST_net_14501;
wire TIMEBOOST_net_16194;
wire g65024_sb;
wire g65025_sb;
wire g65026_sb;
wire g65027_sb;
wire TIMEBOOST_net_15689;
wire g65028_sb;
wire TIMEBOOST_net_12332;
wire g65029_sb;
wire g65030_sb;
wire TIMEBOOST_net_12333;
wire g65031_sb;
wire g58284_da;
wire TIMEBOOST_net_12368;
wire g65032_sb;
wire TIMEBOOST_net_16720;
wire g65033_db;
wire g65033_sb;
wire TIMEBOOST_net_16456;
wire g65034_sb;
wire TIMEBOOST_net_10880;
wire g65035_sb;
wire TIMEBOOST_net_22114;
wire TIMEBOOST_net_21824;
wire g65036_sb;
wire TIMEBOOST_net_12346;
wire TIMEBOOST_net_22859;
wire g65037_sb;
wire TIMEBOOST_net_22787;
wire g65038_sb;
wire TIMEBOOST_net_22727;
wire g65039_sb;
wire g65040_sb;
wire TIMEBOOST_net_14601;
wire g65041_sb;
wire TIMEBOOST_net_16481;
wire TIMEBOOST_net_12567;
wire g65042_sb;
wire TIMEBOOST_net_8106;
wire g65043_sb;
wire g65044_sb;
wire TIMEBOOST_net_21251;
wire TIMEBOOST_net_12823;
wire g65045_sb;
wire TIMEBOOST_net_16428;
wire g65046_sb;
wire n_4283;
wire g65047_sb;
wire TIMEBOOST_net_16480;
wire TIMEBOOST_net_22068;
wire g65048_sb;
wire g65049_sb;
wire TIMEBOOST_net_22890;
wire TIMEBOOST_net_12335;
wire g65050_sb;
wire TIMEBOOST_net_14318;
wire TIMEBOOST_net_20453;
wire g65051_sb;
wire TIMEBOOST_net_14048;
wire g65052_sb;
wire TIMEBOOST_net_17578;
wire g65053_sb;
wire TIMEBOOST_net_13830;
wire TIMEBOOST_net_17265;
wire g65054_sb;
wire TIMEBOOST_net_21674;
wire g65055_sb;
wire TIMEBOOST_net_7130;
wire g65056_sb;
wire g65057_db;
wire g65057_sb;
wire TIMEBOOST_net_13866;
wire g65058_db;
wire g65058_sb;
wire TIMEBOOST_net_13868;
wire g65059_sb;
wire TIMEBOOST_net_22777;
wire g65060_sb;
wire TIMEBOOST_net_21883;
wire g65061_sb;
wire TIMEBOOST_net_23235;
wire g65062_sb;
wire TIMEBOOST_net_16424;
wire g65063_db;
wire g65063_sb;
wire TIMEBOOST_net_15661;
wire g65064_sb;
wire TIMEBOOST_net_10232;
wire g65065_db;
wire g65065_sb;
wire TIMEBOOST_net_14024;
wire g65066_sb;
wire TIMEBOOST_net_261;
wire TIMEBOOST_net_22486;
wire g65067_sb;
wire TIMEBOOST_net_262;
wire TIMEBOOST_net_14951;
wire g65068_sb;
wire TIMEBOOST_net_22425;
wire g65069_db;
wire g65069_sb;
wire TIMEBOOST_net_21553;
wire g65070_sb;
wire g54317_db;
wire g65071_sb;
wire g65072_db;
wire g65072_sb;
wire TIMEBOOST_net_21550;
wire TIMEBOOST_net_12336;
wire g65073_sb;
wire TIMEBOOST_net_13039;
wire TIMEBOOST_net_12337;
wire g65074_sb;
wire TIMEBOOST_net_20986;
wire g65075_sb;
wire TIMEBOOST_net_16525;
wire TIMEBOOST_net_12338;
wire g65076_sb;
wire TIMEBOOST_net_16990;
wire g65077_db;
wire g65077_sb;
wire TIMEBOOST_net_13911;
wire TIMEBOOST_net_12339;
wire g65078_sb;
wire TIMEBOOST_net_17567;
wire g65079_db;
wire g65079_sb;
wire TIMEBOOST_net_13912;
wire TIMEBOOST_net_12340;
wire g65080_sb;
wire g65081_sb;
wire TIMEBOOST_net_13913;
wire TIMEBOOST_net_17215;
wire g65082_sb;
wire g65083_sb;
wire TIMEBOOST_net_13914;
wire TIMEBOOST_net_17216;
wire g65084_sb;
wire TIMEBOOST_net_20209;
wire g65085_sb;
wire TIMEBOOST_net_16523;
wire TIMEBOOST_net_12341;
wire g65086_sb;
wire TIMEBOOST_net_22857;
wire g65087_sb;
wire TIMEBOOST_net_13919;
wire TIMEBOOST_net_12342;
wire g65088_sb;
wire TIMEBOOST_net_13591;
wire g65089_sb;
wire TIMEBOOST_net_13918;
wire g65090_sb;
wire TIMEBOOST_net_15325;
wire g65091_sb;
wire TIMEBOOST_net_263;
wire TIMEBOOST_net_21481;
wire g65092_sb;
wire g65093_db;
wire g65093_sb;
wire TIMEBOOST_net_13040;
wire g65094_sb;
wire TIMEBOOST_net_13920;
wire g65095_sb;
wire g65096_db;
wire g65096_sb;
wire TIMEBOOST_net_13921;
wire g67069_db;
wire g65097_sb;
wire TIMEBOOST_net_13878;
wire g65098_sb;
wire g65099_db;
wire g65099_sb;
wire TIMEBOOST_net_13360;
wire TIMEBOOST_net_188;
wire g65210_sb;
wire TIMEBOOST_net_12866;
wire TIMEBOOST_net_189;
wire g65211_sb;
wire g58360_db;
wire g65212_db;
wire TIMEBOOST_net_13361;
wire TIMEBOOST_net_190;
wire g65213_sb;
wire TIMEBOOST_net_13616;
wire TIMEBOOST_net_15496;
wire g65214_sb;
wire TIMEBOOST_net_16604;
wire g65215_sb;
wire TIMEBOOST_net_9359;
wire g65216_sb;
wire TIMEBOOST_net_23408;
wire TIMEBOOST_net_193;
wire g65217_sb;
wire TIMEBOOST_net_14982;
wire TIMEBOOST_net_12584;
wire g65218_sb;
wire TIMEBOOST_net_20978;
wire TIMEBOOST_net_195;
wire g65219_sb;
wire TIMEBOOST_net_21188;
wire g65220_sb;
wire g65221_sb;
wire TIMEBOOST_net_198;
wire g65222_sb;
wire TIMEBOOST_net_14783;
wire TIMEBOOST_net_199;
wire g65223_sb;
wire TIMEBOOST_net_200;
wire g65224_sb;
wire TIMEBOOST_net_23375;
wire TIMEBOOST_net_22310;
wire g65225_sb;
wire TIMEBOOST_net_22116;
wire TIMEBOOST_net_202;
wire g65226_sb;
wire TIMEBOOST_net_8560;
wire g65227_sb;
wire g65228_sb;
wire TIMEBOOST_net_8563;
wire g65229_sb;
wire TIMEBOOST_net_17306;
wire g65230_sb;
wire TIMEBOOST_net_14334;
wire TIMEBOOST_net_206;
wire g65231_sb;
wire TIMEBOOST_net_9363;
wire g65232_sb;
wire g65233_sb;
wire g65235_sb;
wire TIMEBOOST_net_16609;
wire TIMEBOOST_net_14921;
wire g65236_sb;
wire TIMEBOOST_net_16775;
wire TIMEBOOST_net_211;
wire g65237_sb;
wire TIMEBOOST_net_8552;
wire g65238_sb;
wire g65240_sb;
wire g65241_sb;
wire TIMEBOOST_net_13359;
wire g65242_sb;
wire TIMEBOOST_net_12928;
wire TIMEBOOST_net_216;
wire g65243_sb;
wire g63616_db;
wire TIMEBOOST_net_217;
wire g65244_sb;
wire TIMEBOOST_net_9502;
wire g65245_sb;
wire TIMEBOOST_net_22574;
wire g65246_sb;
wire TIMEBOOST_net_22442;
wire g65247_sb;
wire TIMEBOOST_net_20606;
wire TIMEBOOST_net_9364;
wire g65248_sb;
wire TIMEBOOST_net_12816;
wire TIMEBOOST_net_9365;
wire g65249_sb;
wire TIMEBOOST_net_307;
wire TIMEBOOST_net_23407;
wire g65250_sb;
wire TIMEBOOST_net_22135;
wire g65251_sb;
wire g65252_sb;
wire g65254_p;
wire g65255_p;
wire g58355_db;
wire g65257_p;
wire g65258_p;
wire g65259_p;
wire g65260_p;
wire g65261_p;
wire TIMEBOOST_net_13085;
wire g65262_sb;
wire g65263_p;
wire g65264_p;
wire g65265_p;
wire g65266_p;
wire g65267_p;
wire g65268_da;
wire g65268_db;
wire g65268_sb;
wire TIMEBOOST_net_17021;
wire TIMEBOOST_net_16002;
wire g65269_sb;
wire TIMEBOOST_net_31;
wire g65270_sb;
wire TIMEBOOST_net_13922;
wire g65271_sb;
wire TIMEBOOST_net_13391;
wire TIMEBOOST_net_16436;
wire g65272_sb;
wire TIMEBOOST_net_12828;
wire TIMEBOOST_net_13923;
wire g65273_sb;
wire TIMEBOOST_net_12687;
wire TIMEBOOST_net_13924;
wire g65274_sb;
wire TIMEBOOST_net_12829;
wire TIMEBOOST_net_8227;
wire g65275_sb;
wire TIMEBOOST_net_21071;
wire g65276_sb;
wire TIMEBOOST_net_12818;
wire TIMEBOOST_net_14000;
wire g65277_sb;
wire TIMEBOOST_net_12832;
wire TIMEBOOST_net_13925;
wire g65278_sb;
wire TIMEBOOST_net_12833;
wire g65279_sb;
wire TIMEBOOST_net_12834;
wire TIMEBOOST_net_20399;
wire g65280_sb;
wire TIMEBOOST_net_12808;
wire g65281_sb;
wire TIMEBOOST_net_13926;
wire g65282_sb;
wire TIMEBOOST_net_17417;
wire g65283_sb;
wire g65284_sb;
wire TIMEBOOST_net_12838;
wire TIMEBOOST_net_16416;
wire g65285_sb;
wire TIMEBOOST_net_13974;
wire g65286_sb;
wire TIMEBOOST_net_14307;
wire TIMEBOOST_net_12380;
wire g65287_sb;
wire g65288_db;
wire g65288_sb;
wire TIMEBOOST_net_12837;
wire TIMEBOOST_net_22651;
wire g65289_sb;
wire TIMEBOOST_net_9485;
wire TIMEBOOST_net_13536;
wire g65291_sb;
wire TIMEBOOST_net_16443;
wire g65292_sb;
wire TIMEBOOST_net_12839;
wire TIMEBOOST_net_13907;
wire g65293_sb;
wire TIMEBOOST_net_12688;
wire TIMEBOOST_net_16444;
wire g65294_sb;
wire TIMEBOOST_net_20974;
wire g65295_sb;
wire TIMEBOOST_net_22531;
wire g65296_sb;
wire TIMEBOOST_net_12689;
wire TIMEBOOST_net_16414;
wire g65297_sb;
wire g65298_db;
wire g65298_sb;
wire TIMEBOOST_net_22199;
wire g65299_sb;
wire TIMEBOOST_net_16433;
wire g65300_sb;
wire TIMEBOOST_net_13086;
wire g65301_sb;
wire TIMEBOOST_net_13967;
wire TIMEBOOST_net_12412;
wire g65302_sb;
wire TIMEBOOST_net_12840;
wire TIMEBOOST_net_13910;
wire g65303_sb;
wire g65304_sb;
wire TIMEBOOST_net_14008;
wire TIMEBOOST_net_13908;
wire g65305_sb;
wire TIMEBOOST_net_13909;
wire g65306_sb;
wire TIMEBOOST_net_22048;
wire g65307_sb;
wire TIMEBOOST_net_12693;
wire TIMEBOOST_net_16415;
wire g65308_sb;
wire g65309_da;
wire g65309_sb;
wire g65310_sb;
wire TIMEBOOST_net_20541;
wire g65311_sb;
wire TIMEBOOST_net_10423;
wire TIMEBOOST_net_14932;
wire g65312_sb;
wire TIMEBOOST_net_8807;
wire TIMEBOOST_net_14937;
wire g65313_sb;
wire TIMEBOOST_net_8808;
wire g65314_sb;
wire TIMEBOOST_net_13038;
wire TIMEBOOST_net_14944;
wire g65315_sb;
wire TIMEBOOST_net_12696;
wire g65316_sb;
wire TIMEBOOST_net_8810;
wire TIMEBOOST_net_17428;
wire g65317_sb;
wire TIMEBOOST_net_13369;
wire g65318_sb;
wire TIMEBOOST_net_8788;
wire TIMEBOOST_net_17266;
wire g65319_sb;
wire TIMEBOOST_net_12699;
wire TIMEBOOST_net_13916;
wire g65320_sb;
wire g65321_sb;
wire TIMEBOOST_net_13917;
wire g65322_sb;
wire g65323_sb;
wire g65324_da;
wire TIMEBOOST_net_15931;
wire g65324_sb;
wire g65325_da;
wire TIMEBOOST_net_147;
wire g65325_sb;
wire g58449_db;
wire g65326_sb;
wire TIMEBOOST_net_20877;
wire g65327_sb;
wire TIMEBOOST_net_13371;
wire TIMEBOOST_net_22015;
wire g65328_sb;
wire TIMEBOOST_net_12703;
wire g58445_db;
wire g65329_sb;
wire TIMEBOOST_net_12704;
wire TIMEBOOST_net_21482;
wire g65330_sb;
wire TIMEBOOST_net_12705;
wire g65331_sb;
wire TIMEBOOST_net_8789;
wire g65332_db;
wire g65332_sb;
wire TIMEBOOST_net_15182;
wire g65333_sb;
wire g65334_sb;
wire TIMEBOOST_net_14668;
wire g65335_db;
wire g65335_sb;
wire TIMEBOOST_net_13955;
wire g65336_sb;
wire TIMEBOOST_net_12708;
wire g65337_sb;
wire g65338_db;
wire g65338_sb;
wire TIMEBOOST_net_12835;
wire TIMEBOOST_net_14890;
wire g65339_sb;
wire g65340_sb;
wire TIMEBOOST_net_16643;
wire g65341_sb;
wire TIMEBOOST_net_8797;
wire g65342_sb;
wire TIMEBOOST_net_12710;
wire g65343_sb;
wire TIMEBOOST_net_8800;
wire g65345_sb;
wire TIMEBOOST_net_8786;
wire g65346_sb;
wire TIMEBOOST_net_13052;
wire g65347_sb;
wire TIMEBOOST_net_13997;
wire TIMEBOOST_net_16454;
wire g65348_sb;
wire TIMEBOOST_net_17454;
wire g65349_sb;
wire TIMEBOOST_net_13053;
wire TIMEBOOST_net_8225;
wire g65350_sb;
wire TIMEBOOST_net_23374;
wire TIMEBOOST_net_21738;
wire g65351_sb;
wire TIMEBOOST_net_14045;
wire TIMEBOOST_net_12791;
wire g65352_sb;
wire TIMEBOOST_net_17274;
wire g65353_sb;
wire TIMEBOOST_net_12738;
wire TIMEBOOST_net_16455;
wire g65354_sb;
wire g65355_sb;
wire TIMEBOOST_net_13748;
wire TIMEBOOST_net_15817;
wire g65356_sb;
wire TIMEBOOST_net_13055;
wire TIMEBOOST_net_21687;
wire g65357_sb;
wire TIMEBOOST_net_13056;
wire g65858_db;
wire g65358_sb;
wire TIMEBOOST_net_13057;
wire g65359_sb;
wire TIMEBOOST_net_12734;
wire g65360_sb;
wire TIMEBOOST_net_13058;
wire g65361_sb;
wire TIMEBOOST_net_12724;
wire TIMEBOOST_net_12792;
wire g65362_sb;
wire TIMEBOOST_net_22062;
wire TIMEBOOST_net_21432;
wire g65363_sb;
wire TIMEBOOST_net_13059;
wire TIMEBOOST_net_8632;
wire g65364_sb;
wire TIMEBOOST_net_12720;
wire TIMEBOOST_net_16511;
wire g65365_sb;
wire TIMEBOOST_net_12711;
wire TIMEBOOST_net_22148;
wire g65366_sb;
wire TIMEBOOST_net_22208;
wire g65367_sb;
wire TIMEBOOST_net_12831;
wire TIMEBOOST_net_20794;
wire g65368_sb;
wire TIMEBOOST_net_22102;
wire TIMEBOOST_net_14938;
wire g65369_sb;
wire TIMEBOOST_net_12712;
wire g65370_sb;
wire g65371_da;
wire g62805_db;
wire TIMEBOOST_net_12842;
wire g65372_sb;
wire g65373_sb;
wire TIMEBOOST_net_8787;
wire TIMEBOOST_net_14930;
wire g65374_sb;
wire TIMEBOOST_net_14013;
wire g58419_db;
wire g65375_sb;
wire g65376_sb;
wire TIMEBOOST_net_9484;
wire g65377_sb;
wire TIMEBOOST_net_12714;
wire g58409_db;
wire g65378_sb;
wire g58408_db;
wire g65379_sb;
wire TIMEBOOST_net_23405;
wire g65380_sb;
wire TIMEBOOST_net_13060;
wire g65381_sb;
wire TIMEBOOST_net_8634;
wire g65382_sb;
wire TIMEBOOST_net_13062;
wire TIMEBOOST_net_21678;
wire g65383_sb;
wire TIMEBOOST_net_22144;
wire TIMEBOOST_net_21655;
wire g65384_sb;
wire TIMEBOOST_net_12793;
wire g65385_sb;
wire TIMEBOOST_net_155;
wire TIMEBOOST_net_13063;
wire TIMEBOOST_net_21748;
wire g65387_sb;
wire TIMEBOOST_net_12955;
wire TIMEBOOST_net_21049;
wire g65388_sb;
wire TIMEBOOST_net_13064;
wire TIMEBOOST_net_21682;
wire g65389_sb;
wire TIMEBOOST_net_80;
wire g65390_db;
wire g65390_sb;
wire TIMEBOOST_net_21441;
wire g65391_sb;
wire TIMEBOOST_net_13065;
wire TIMEBOOST_net_21806;
wire g65392_sb;
wire TIMEBOOST_net_12758;
wire g65393_sb;
wire TIMEBOOST_net_13747;
wire TIMEBOOST_net_21596;
wire g65394_sb;
wire TIMEBOOST_net_17371;
wire g65395_sb;
wire TIMEBOOST_net_13066;
wire g65396_sb;
wire TIMEBOOST_net_22145;
wire g65397_sb;
wire TIMEBOOST_net_12830;
wire TIMEBOOST_net_21085;
wire g65398_sb;
wire TIMEBOOST_net_12716;
wire g65399_sb;
wire TIMEBOOST_net_12717;
wire g65400_sb;
wire TIMEBOOST_net_13067;
wire TIMEBOOST_net_21763;
wire g65401_sb;
wire TIMEBOOST_net_12718;
wire g58364_db;
wire g65402_sb;
wire g58363_db;
wire g65403_sb;
wire TIMEBOOST_net_12719;
wire g58361_db;
wire g65404_sb;
wire TIMEBOOST_net_20717;
wire g65405_sb;
wire TIMEBOOST_net_12721;
wire g65406_sb;
wire g65407_sb;
wire TIMEBOOST_net_13068;
wire g65408_sb;
wire TIMEBOOST_net_12722;
wire g58352_db;
wire g65409_sb;
wire TIMEBOOST_net_14893;
wire g65410_sb;
wire TIMEBOOST_net_9561;
wire TIMEBOOST_net_12723;
wire g58345_db;
wire g65412_sb;
wire TIMEBOOST_net_13485;
wire g65413_sb;
wire TIMEBOOST_net_22067;
wire TIMEBOOST_net_8277;
wire g65414_sb;
wire TIMEBOOST_net_12725;
wire TIMEBOOST_net_16642;
wire g65415_sb;
wire TIMEBOOST_net_12726;
wire g58328_db;
wire g65416_sb;
wire TIMEBOOST_net_12727;
wire g65417_sb;
wire TIMEBOOST_net_12728;
wire g58327_db;
wire g65418_sb;
wire TIMEBOOST_net_9428;
wire TIMEBOOST_net_21999;
wire TIMEBOOST_net_20359;
wire g65421_sb;
wire TIMEBOOST_net_22040;
wire g58311_db;
wire g65422_sb;
wire TIMEBOOST_net_21998;
wire g58305_db;
wire g65423_sb;
wire TIMEBOOST_net_12730;
wire TIMEBOOST_net_21829;
wire g65424_sb;
wire TIMEBOOST_net_9486;
wire g65425_db;
wire g65425_sb;
wire TIMEBOOST_net_22002;
wire g65426_sb;
wire TIMEBOOST_net_22010;
wire g65427_sb;
wire TIMEBOOST_net_22215;
wire g65428_sb;
wire TIMEBOOST_net_12731;
wire TIMEBOOST_net_21804;
wire g65429_sb;
wire TIMEBOOST_net_12732;
wire g58265_db;
wire g65430_sb;
wire TIMEBOOST_net_21414;
wire g65431_sb;
wire g65432_sb;
wire TIMEBOOST_net_12733;
wire TIMEBOOST_net_22454;
wire g65433_sb;
wire TIMEBOOST_net_22091;
wire g65434_sb;
wire TIMEBOOST_net_12735;
wire TIMEBOOST_net_16524;
wire g65435_sb;
wire g65436_p;
wire g65437_p;
wire g65439_p;
wire g65486_p;
wire g65488_p;
wire g65489_p;
wire g65490_p;
wire g65491_p;
wire g65493_p;
wire g65495_p;
wire g65497_p;
wire g65498_p;
wire g65510_p;
wire g65511_p;
wire g65513_p;
wire g65514_p;
wire g65515_p;
wire g65517_p;
wire g65518_p;
wire g65520_p;
wire g65522_p1;
wire g65522_p2;
wire g65523_p;
wire g65530_p;
wire g65533_p;
wire g65543_p;
wire g65549_p;
wire g65550_p;
wire g65555_p;
wire g65557_p;
wire g65559_p;
wire g65562_p;
wire g65567_p;
wire g65568_p;
wire g65569_p;
wire g65570_p;
wire g65571_p;
wire g65572_p1;
wire g65572_p2;
wire g65573_p;
wire g65583_p;
wire g65588_p;
wire g65590_p;
wire g65595_p;
wire g65614_p;
wire g65617_p;
wire g65626_p;
wire TIMEBOOST_net_9384;
wire g65668_sb;
wire TIMEBOOST_net_23212;
wire g65669_sb;
wire TIMEBOOST_net_16479;
wire TIMEBOOST_net_21466;
wire g65670_sb;
wire TIMEBOOST_net_14474;
wire g65671_db;
wire g65671_sb;
wire g65672_sb;
wire g65673_sb;
wire g62757_db;
wire g65674_sb;
wire g65675_sb;
wire TIMEBOOST_net_23406;
wire g65676_sb;
wire TIMEBOOST_net_9562;
wire g65677_sb;
wire TIMEBOOST_net_15999;
wire g65678_sb;
wire TIMEBOOST_net_9385;
wire TIMEBOOST_net_22443;
wire g65679_sb;
wire TIMEBOOST_net_16606;
wire TIMEBOOST_net_23453;
wire g65680_sb;
wire g65681_db;
wire g65681_sb;
wire TIMEBOOST_net_9190;
wire TIMEBOOST_net_21911;
wire g65682_sb;
wire TIMEBOOST_net_8598;
wire g65683_sb;
wire TIMEBOOST_net_9386;
wire g65684_sb;
wire TIMEBOOST_net_16001;
wire g65685_sb;
wire TIMEBOOST_net_16000;
wire TIMEBOOST_net_17008;
wire g65686_sb;
wire TIMEBOOST_net_9563;
wire g65687_sb;
wire g65688_sb;
wire TIMEBOOST_net_16585;
wire TIMEBOOST_net_17009;
wire g65689_sb;
wire TIMEBOOST_net_21412;
wire TIMEBOOST_net_12490;
wire g65690_sb;
wire TIMEBOOST_net_9387;
wire g65691_db;
wire g65691_sb;
wire TIMEBOOST_net_16527;
wire g65692_sb;
wire TIMEBOOST_net_22555;
wire TIMEBOOST_net_12491;
wire g65693_sb;
wire TIMEBOOST_net_12347;
wire g65694_sb;
wire TIMEBOOST_net_9505;
wire g65695_sb;
wire g65696_sb;
wire TIMEBOOST_net_15989;
wire g65697_db;
wire g65697_sb;
wire TIMEBOOST_net_16324;
wire TIMEBOOST_net_22519;
wire g65698_sb;
wire TIMEBOOST_net_22953;
wire g65699_sb;
wire TIMEBOOST_net_9506;
wire g65700_sb;
wire TIMEBOOST_net_16650;
wire g65701_db;
wire g65701_sb;
wire TIMEBOOST_net_8600;
wire TIMEBOOST_net_17322;
wire g65702_sb;
wire TIMEBOOST_net_16586;
wire TIMEBOOST_net_17010;
wire g65703_sb;
wire TIMEBOOST_net_21376;
wire TIMEBOOST_net_12472;
wire g65704_sb;
wire TIMEBOOST_net_21523;
wire g65705_db;
wire g65705_sb;
wire g65706_sb;
wire TIMEBOOST_net_20924;
wire g65707_sb;
wire g65708_sb;
wire TIMEBOOST_net_20415;
wire g65709_sb;
wire g65710_sb;
wire TIMEBOOST_net_9508;
wire g65711_sb;
wire TIMEBOOST_net_15988;
wire TIMEBOOST_net_23512;
wire g65712_sb;
wire g58326_db;
wire g65713_db;
wire g65713_sb;
wire TIMEBOOST_net_9388;
wire g65714_db;
wire g65714_sb;
wire TIMEBOOST_net_9389;
wire g65715_sb;
wire g65716_db;
wire TIMEBOOST_net_22236;
wire g65717_db;
wire g65717_sb;
wire TIMEBOOST_net_16437;
wire TIMEBOOST_net_14428;
wire g65718_sb;
wire TIMEBOOST_net_21543;
wire g65719_sb;
wire TIMEBOOST_net_17323;
wire g65720_sb;
wire g65721_sb;
wire TIMEBOOST_net_21470;
wire g65722_sb;
wire TIMEBOOST_net_22217;
wire TIMEBOOST_net_20265;
wire g65723_sb;
wire TIMEBOOST_net_22432;
wire g65724_db;
wire g65724_sb;
wire g65725_sb;
wire TIMEBOOST_net_16656;
wire g65726_sb;
wire TIMEBOOST_net_12851;
wire g65727_sb;
wire TIMEBOOST_net_14349;
wire g65728_sb;
wire g65729_p;
wire TIMEBOOST_net_21012;
wire g65730_sb;
wire TIMEBOOST_net_21288;
wire TIMEBOOST_net_17221;
wire g65731_sb;
wire TIMEBOOST_net_8602;
wire g65732_sb;
wire TIMEBOOST_net_16339;
wire g65733_db;
wire g65733_sb;
wire TIMEBOOST_net_9390;
wire g65734_db;
wire g65734_sb;
wire TIMEBOOST_net_16207;
wire TIMEBOOST_net_17307;
wire g65735_sb;
wire TIMEBOOST_net_8538;
wire TIMEBOOST_net_17308;
wire g65736_sb;
wire TIMEBOOST_net_9391;
wire g65737_db;
wire g65737_sb;
wire TIMEBOOST_net_16503;
wire g65738_sb;
wire g65739_sb;
wire TIMEBOOST_net_16504;
wire TIMEBOOST_net_21912;
wire g65740_sb;
wire TIMEBOOST_net_16722;
wire g65741_db;
wire g65741_sb;
wire TIMEBOOST_net_16505;
wire g65742_sb;
wire TIMEBOOST_net_20277;
wire TIMEBOOST_net_21951;
wire g65743_sb;
wire TIMEBOOST_net_16425;
wire g65744_sb;
wire g65745_sb;
wire TIMEBOOST_net_16502;
wire TIMEBOOST_net_12354;
wire g65746_sb;
wire TIMEBOOST_net_8603;
wire TIMEBOOST_net_23053;
wire g65747_sb;
wire TIMEBOOST_net_12850;
wire TIMEBOOST_net_10857;
wire g65748_sb;
wire g65749_db;
wire g65749_sb;
wire TIMEBOOST_net_9333;
wire TIMEBOOST_net_17055;
wire g65750_sb;
wire TIMEBOOST_net_8604;
wire TIMEBOOST_net_17324;
wire g65751_sb;
wire g65752_sb;
wire TIMEBOOST_net_9392;
wire g65753_db;
wire g65753_sb;
wire TIMEBOOST_net_20457;
wire g65754_db;
wire g65754_sb;
wire TIMEBOOST_net_22235;
wire TIMEBOOST_net_17056;
wire g65755_sb;
wire g58309_db;
wire g65756_db;
wire g65756_sb;
wire TIMEBOOST_net_22214;
wire TIMEBOOST_net_23167;
wire TIMEBOOST_net_14865;
wire g65758_sb;
wire TIMEBOOST_net_16442;
wire TIMEBOOST_net_22463;
wire g65759_sb;
wire TIMEBOOST_net_9334;
wire g65760_db;
wire g65760_sb;
wire TIMEBOOST_net_9331;
wire g65761_sb;
wire TIMEBOOST_net_14358;
wire g65762_sb;
wire TIMEBOOST_net_9393;
wire g65763_db;
wire TIMEBOOST_net_9394;
wire g65764_db;
wire g65764_sb;
wire TIMEBOOST_net_13394;
wire g65765_db;
wire TIMEBOOST_net_12849;
wire TIMEBOOST_net_12475;
wire g65766_sb;
wire TIMEBOOST_net_14378;
wire g65767_sb;
wire TIMEBOOST_net_8539;
wire TIMEBOOST_net_12476;
wire g65768_sb;
wire TIMEBOOST_net_9395;
wire TIMEBOOST_net_22888;
wire g65769_sb;
wire TIMEBOOST_net_9396;
wire g65770_db;
wire g65770_sb;
wire TIMEBOOST_net_8540;
wire TIMEBOOST_net_17309;
wire g65771_sb;
wire TIMEBOOST_net_16340;
wire TIMEBOOST_net_17011;
wire g65772_sb;
wire TIMEBOOST_net_8605;
wire TIMEBOOST_net_21937;
wire g65773_sb;
wire g65774_sb;
wire TIMEBOOST_net_22513;
wire g65775_sb;
wire TIMEBOOST_net_22370;
wire TIMEBOOST_net_13347;
wire g65776_sb;
wire TIMEBOOST_net_9335;
wire g65777_db;
wire g65777_sb;
wire g58291_db;
wire TIMEBOOST_net_21625;
wire g65778_sb;
wire TIMEBOOST_net_14375;
wire g65779_sb;
wire TIMEBOOST_net_22362;
wire g65780_db;
wire g65780_sb;
wire TIMEBOOST_net_16658;
wire g65781_db;
wire g65781_sb;
wire g58286_db;
wire g65782_db;
wire g65782_sb;
wire TIMEBOOST_net_8541;
wire g65783_sb;
wire TIMEBOOST_net_22440;
wire g65784_sb;
wire TIMEBOOST_net_9397;
wire TIMEBOOST_net_15480;
wire TIMEBOOST_net_8542;
wire TIMEBOOST_net_12477;
wire g65786_sb;
wire g65787_sb;
wire TIMEBOOST_net_8543;
wire g65788_db;
wire g65788_sb;
wire TIMEBOOST_net_22363;
wire TIMEBOOST_net_15520;
wire g65789_sb;
wire TIMEBOOST_net_17057;
wire g65790_sb;
wire TIMEBOOST_net_17310;
wire g65791_sb;
wire TIMEBOOST_net_9336;
wire g65792_sb;
wire TIMEBOOST_net_13364;
wire g65793_sb;
wire g58280_db;
wire TIMEBOOST_net_14575;
wire g65794_sb;
wire g65795_db;
wire g65795_sb;
wire TIMEBOOST_net_9398;
wire TIMEBOOST_net_9509;
wire g65797_sb;
wire TIMEBOOST_net_17312;
wire g65798_sb;
wire TIMEBOOST_net_13372;
wire g65799_sb;
wire TIMEBOOST_net_22259;
wire TIMEBOOST_net_20236;
wire g65800_sb;
wire g65801_p;
wire TIMEBOOST_net_16692;
wire g65802_sb;
wire TIMEBOOST_net_15983;
wire TIMEBOOST_net_15525;
wire g65803_sb;
wire TIMEBOOST_net_14259;
wire g65804_sb;
wire TIMEBOOST_net_9337;
wire g59797_db;
wire g65805_sb;
wire TIMEBOOST_net_9338;
wire TIMEBOOST_net_15978;
wire g65806_sb;
wire TIMEBOOST_net_8606;
wire g65807_db;
wire g65807_sb;
wire TIMEBOOST_net_13699;
wire TIMEBOOST_net_15663;
wire g65808_p;
wire TIMEBOOST_net_21579;
wire g65809_db;
wire g65809_sb;
wire g65810_sb;
wire g65811_sb;
wire g65812_db;
wire g65812_sb;
wire TIMEBOOST_net_14311;
wire g65813_sb;
wire g65814_db;
wire g65814_sb;
wire TIMEBOOST_net_23460;
wire g65815_db;
wire g65815_sb;
wire g65816_db;
wire g65816_sb;
wire g65817_db;
wire TIMEBOOST_net_22051;
wire g65818_db;
wire g65818_sb;
wire TIMEBOOST_net_16771;
wire TIMEBOOST_net_21923;
wire g65819_sb;
wire g65820_db;
wire g65820_sb;
wire TIMEBOOST_net_12923;
wire TIMEBOOST_net_22413;
wire g65821_sb;
wire TIMEBOOST_net_13697;
wire g65822_db;
wire g65822_sb;
wire TIMEBOOST_net_12895;
wire TIMEBOOST_net_21746;
wire g65823_sb;
wire TIMEBOOST_net_22714;
wire g65824_sb;
wire TIMEBOOST_net_22049;
wire TIMEBOOST_net_17460;
wire g65825_sb;
wire TIMEBOOST_net_12796;
wire g65826_sb;
wire TIMEBOOST_net_22039;
wire TIMEBOOST_net_22073;
wire g65827_sb;
wire TIMEBOOST_net_13489;
wire g65828_db;
wire g65828_sb;
wire TIMEBOOST_net_12709;
wire g65829_sb;
wire TIMEBOOST_net_22028;
wire g65830_sb;
wire TIMEBOOST_net_13888;
wire TIMEBOOST_net_12799;
wire g65831_sb;
wire TIMEBOOST_net_22482;
wire TIMEBOOST_net_12800;
wire g65832_sb;
wire TIMEBOOST_net_12707;
wire TIMEBOOST_net_17550;
wire g65833_sb;
wire g65834_sb;
wire TIMEBOOST_net_93;
wire g65835_sb;
wire TIMEBOOST_net_12702;
wire g65836_db;
wire g65836_sb;
wire TIMEBOOST_net_22022;
wire TIMEBOOST_net_12803;
wire g65837_sb;
wire g65838_sb;
wire TIMEBOOST_net_14029;
wire g65839_db;
wire g65839_sb;
wire g65840_sb;
wire TIMEBOOST_net_21304;
wire g65841_sb;
wire TIMEBOOST_net_17461;
wire g65842_sb;
wire g65843_db;
wire g65843_sb;
wire TIMEBOOST_net_23128;
wire TIMEBOOST_net_17462;
wire g65844_sb;
wire TIMEBOOST_net_12697;
wire g65845_db;
wire g65845_sb;
wire TIMEBOOST_net_22013;
wire TIMEBOOST_net_12804;
wire g65846_sb;
wire g65847_db;
wire g65847_sb;
wire g65848_sb;
wire TIMEBOOST_net_21919;
wire g65849_db;
wire g65849_sb;
wire TIMEBOOST_net_13666;
wire g65850_sb;
wire TIMEBOOST_net_9339;
wire g65851_db;
wire g65851_sb;
wire TIMEBOOST_net_16018;
wire g65852_sb;
wire TIMEBOOST_net_17029;
wire g65853_db;
wire g65853_sb;
wire g65854_db;
wire g65854_sb;
wire g65855_sb;
wire TIMEBOOST_net_13995;
wire g65856_sb;
wire TIMEBOOST_net_121;
wire TIMEBOOST_net_7524;
wire g65857_sb;
wire TIMEBOOST_net_23161;
wire TIMEBOOST_net_20433;
wire g65858_sb;
wire g65859_sb;
wire g65860_db;
wire g65860_sb;
wire TIMEBOOST_net_94;
wire g65861_sb;
wire g65862_da;
wire g65862_db;
wire g65862_sb;
wire TIMEBOOST_net_122;
wire TIMEBOOST_net_13567;
wire g65863_sb;
wire TIMEBOOST_net_16508;
wire TIMEBOOST_net_123;
wire g65865_db;
wire g65865_sb;
wire g65866_db;
wire g65866_sb;
wire g65867_db;
wire g65867_sb;
wire TIMEBOOST_net_13698;
wire g65868_db;
wire g65868_sb;
wire TIMEBOOST_net_22023;
wire g65869_sb;
wire n_15457;
wire g65870_db;
wire g65870_sb;
wire TIMEBOOST_net_12852;
wire g65871_sb;
wire TIMEBOOST_net_23165;
wire TIMEBOOST_net_17463;
wire g65872_sb;
wire g65873_db;
wire g65873_sb;
wire g65874_db;
wire g65874_sb;
wire g65875_db;
wire g65875_sb;
wire TIMEBOOST_net_13806;
wire TIMEBOOST_net_17284;
wire g65876_sb;
wire TIMEBOOST_net_21162;
wire g65877_sb;
wire TIMEBOOST_net_9340;
wire g65878_db;
wire g65878_sb;
wire TIMEBOOST_net_15515;
wire g65879_sb;
wire g65880_db;
wire g65880_sb;
wire TIMEBOOST_net_21181;
wire g65881_sb;
wire g65882_db;
wire g65882_sb;
wire g65883_sb;
wire TIMEBOOST_net_23491;
wire g65884_db;
wire g65884_sb;
wire TIMEBOOST_net_124;
wire g65885_db;
wire TIMEBOOST_net_125;
wire g65887_sb;
wire TIMEBOOST_net_16421;
wire g65888_sb;
wire g65889_sb;
wire g65890_sb;
wire g65891_sb;
wire TIMEBOOST_net_15320;
wire TIMEBOOST_net_12841;
wire g65892_sb;
wire TIMEBOOST_net_14662;
wire g65893_sb;
wire TIMEBOOST_net_12694;
wire TIMEBOOST_net_17464;
wire g65894_sb;
wire TIMEBOOST_net_126;
wire TIMEBOOST_net_7526;
wire TIMEBOOST_net_301;
wire g65896_db;
wire g65896_sb;
wire TIMEBOOST_net_15730;
wire TIMEBOOST_net_12805;
wire g65897_sb;
wire TIMEBOOST_net_14314;
wire g65899_da;
wire g65899_db;
wire g65899_sb;
wire TIMEBOOST_net_13996;
wire TIMEBOOST_net_12919;
wire g65900_sb;
wire g65901_sb;
wire g65902_da;
wire g65902_db;
wire g65902_sb;
wire TIMEBOOST_net_9341;
wire TIMEBOOST_net_17060;
wire g65903_sb;
wire TIMEBOOST_net_9342;
wire g65904_db;
wire g65904_sb;
wire g65905_da;
wire g65905_sb;
wire g65906_da;
wire g65906_sb;
wire g65907_db;
wire g65907_sb;
wire TIMEBOOST_net_20668;
wire g65908_sb;
wire g65909_sb;
wire TIMEBOOST_net_22381;
wire g65910_db;
wire g65910_sb;
wire TIMEBOOST_net_20198;
wire TIMEBOOST_net_15459;
wire g65912_db;
wire TIMEBOOST_net_8576;
wire TIMEBOOST_net_17285;
wire g65913_sb;
wire TIMEBOOST_net_21778;
wire TIMEBOOST_net_17503;
wire g65914_sb;
wire g65915_db;
wire g65915_sb;
wire TIMEBOOST_net_8790;
wire g65916_sb;
wire TIMEBOOST_net_16680;
wire TIMEBOOST_net_22956;
wire TIMEBOOST_net_13367;
wire g65919_db;
wire g65919_sb;
wire TIMEBOOST_net_13963;
wire g65920_sb;
wire TIMEBOOST_net_22265;
wire g65921_db;
wire g65921_sb;
wire TIMEBOOST_net_16071;
wire TIMEBOOST_net_22276;
wire g65923_db;
wire g65923_sb;
wire TIMEBOOST_net_16672;
wire TIMEBOOST_net_17465;
wire g65924_sb;
wire TIMEBOOST_net_14277;
wire TIMEBOOST_net_22478;
wire TIMEBOOST_net_14278;
wire TIMEBOOST_net_13886;
wire TIMEBOOST_net_14279;
wire TIMEBOOST_net_513;
wire TIMEBOOST_net_14055;
wire TIMEBOOST_net_16495;
wire TIMEBOOST_net_12413;
wire g65931_sb;
wire g65932_p;
wire TIMEBOOST_net_17030;
wire TIMEBOOST_net_7527;
wire TIMEBOOST_net_9343;
wire g65934_db;
wire g65934_sb;
wire TIMEBOOST_net_9344;
wire g65935_sb;
wire g65936_da;
wire g65936_db;
wire g65936_sb;
wire g65937_p;
wire g65938_p;
wire g65939_p;
wire TIMEBOOST_net_11426;
wire g65940_db;
wire g65940_sb;
wire g65942_db;
wire g65942_sb;
wire TIMEBOOST_net_12691;
wire TIMEBOOST_net_12807;
wire g65943_sb;
wire TIMEBOOST_net_515;
wire TIMEBOOST_net_22474;
wire TIMEBOOST_net_16956;
wire TIMEBOOST_net_21572;
wire g65946_db;
wire TIMEBOOST_net_517;
wire TIMEBOOST_net_13883;
wire TIMEBOOST_net_13966;
wire g65949_sb;
wire TIMEBOOST_net_21340;
wire TIMEBOOST_net_7534;
wire g65951_db;
wire g65951_sb;
wire TIMEBOOST_net_302;
wire g65952_db;
wire g65952_sb;
wire TIMEBOOST_net_15197;
wire TIMEBOOST_net_21475;
wire g65953_sb;
wire TIMEBOOST_net_303;
wire TIMEBOOST_net_22988;
wire g65954_sb;
wire TIMEBOOST_net_77;
wire TIMEBOOST_net_16494;
wire n_13467;
wire g65957_db;
wire g65957_sb;
wire TIMEBOOST_net_22299;
wire g65958_db;
wire g65958_sb;
wire TIMEBOOST_net_96;
wire g65959_db;
wire TIMEBOOST_net_22320;
wire g65960_db;
wire g65960_sb;
wire TIMEBOOST_net_97;
wire g65961_db;
wire TIMEBOOST_net_9345;
wire g65962_db;
wire g65962_sb;
wire TIMEBOOST_net_12038;
wire TIMEBOOST_net_13882;
wire TIMEBOOST_net_15330;
wire g65964_sb;
wire TIMEBOOST_net_8609;
wire g65965_sb;
wire TIMEBOOST_net_22118;
wire TIMEBOOST_net_21132;
wire g65966_sb;
wire TIMEBOOST_net_15169;
wire g65967_db;
wire g65967_sb;
wire g65968_db;
wire g65969_sb;
wire TIMEBOOST_net_17355;
wire g65970_sb;
wire TIMEBOOST_net_21783;
wire TIMEBOOST_net_21353;
wire g65971_sb;
wire TIMEBOOST_net_21642;
wire TIMEBOOST_net_21598;
wire g65972_sb;
wire TIMEBOOST_net_98;
wire TIMEBOOST_net_99;
wire TIMEBOOST_net_13880;
wire TIMEBOOST_net_8578;
wire g65976_sb;
wire TIMEBOOST_net_8577;
wire g65977_sb;
wire TIMEBOOST_net_13363;
wire g65978_sb;
wire g65983_p;
wire g65984_p;
wire TIMEBOOST_net_14540;
wire TIMEBOOST_net_9;
wire g65992_p;
wire g65993_p;
wire TIMEBOOST_net_7595;
wire g65994_sb;
wire g65995_da;
wire TIMEBOOST_net_21766;
wire g65996_da;
wire g65996_db;
wire TIMEBOOST_net_15502;
wire TIMEBOOST_net_22290;
wire TIMEBOOST_net_16013;
wire TIMEBOOST_net_9560;
wire g66001_db;
wire g66002_p;
wire g66003_p;
wire g66004_p;
wire g66005_p;
wire g66006_p;
wire g66007_p;
wire g66008_p;
wire g66009_p;
wire g66010_p;
wire g66011_p;
wire g66012_p;
wire g66013_p;
wire g66014_p;
wire g66015_p;
wire g66016_p;
wire g66066_p;
wire g66068_p;
wire g66072_p;
wire g66074_p;
wire g66075_p;
wire g66076_p;
wire g66077_p;
wire g66078_p;
wire g66079_p;
wire g66080_p;
wire g66081_p;
wire g66082_p;
wire g66083_p;
wire g66084_p;
wire g66085_p;
wire g66086_p;
wire g66087_p;
wire g66089_p;
wire g66090_p;
wire g66093_p;
wire g66094_p;
wire g66095_p;
wire g66096_p;
wire g66097_p;
wire g66098_p;
wire g66099_p;
wire g66100_p;
wire g66107_p;
wire g66108_p;
wire g66110_p;
wire g66113_p;
wire g66118_p;
wire g66121_p;
wire g66122_p;
wire g66124_p;
wire g66125_p;
wire g66127_p;
wire g66128_p;
wire g66129_p;
wire g66130_p;
wire g66132_p;
wire g66133_p;
wire g66134_p;
wire g66136_p;
wire g66138_p;
wire g66143_p;
wire g66145_p;
wire g66147_p;
wire g66153_p;
wire g66155_p;
wire g66160_p;
wire g66165_p;
wire g66176_p;
wire g66178_p;
wire g66184_p;
wire g66190_p;
wire g66194_p;
wire g66195_p;
wire g66197_p;
wire g66202_p;
wire g66215_p;
wire g66223_p;
wire g66232_p;
wire g66234_p;
wire g66237_p;
wire g66239_p;
wire g66248_p;
wire g66267_p;
wire g66269_p;
wire g66278_p;
wire g66286_p;
wire g66287_p;
wire g66290_dup_p;
wire g66291_p;
wire g66298_p;
wire g66299_p;
wire g66302_p;
wire g66303_p;
wire g66310_p;
wire g66315_p;
wire g66322_p;
wire g66323_p;
wire g66327_p;
wire g66336_p;
wire g66338_p;
wire g66357_p;
wire g66358_p;
wire TIMEBOOST_net_9399;
wire TIMEBOOST_net_22439;
wire g66397_sb;
wire TIMEBOOST_net_16346;
wire g66398_db;
wire g66398_sb;
wire TIMEBOOST_net_22611;
wire g66399_sb;
wire TIMEBOOST_net_17233;
wire g66400_db;
wire TIMEBOOST_net_9400;
wire TIMEBOOST_net_14115;
wire TIMEBOOST_net_17230;
wire g66402_db;
wire g66402_sb;
wire g66403_db;
wire g66403_sb;
wire TIMEBOOST_net_166;
wire g66404_db;
wire g66405_db;
wire TIMEBOOST_net_9401;
wire g66406_db;
wire g66406_sb;
wire TIMEBOOST_net_168;
wire g66407_db;
wire TIMEBOOST_net_169;
wire g66408_db;
wire TIMEBOOST_net_21516;
wire g66409_db;
wire TIMEBOOST_net_171;
wire g66410_db;
wire TIMEBOOST_net_22306;
wire g66411_db;
wire TIMEBOOST_net_22304;
wire g66412_db;
wire TIMEBOOST_net_17367;
wire g66413_db;
wire TIMEBOOST_net_22273;
wire g66414_db;
wire TIMEBOOST_net_7590;
wire g66415_db;
wire g66415_sb;
wire TIMEBOOST_net_9402;
wire g66416_db;
wire g66417_db;
wire TIMEBOOST_net_9403;
wire g66418_db;
wire TIMEBOOST_net_21631;
wire g66419_db;
wire TIMEBOOST_net_12037;
wire g66420_db;
wire g66421_db;
wire TIMEBOOST_net_16648;
wire g66422_db;
wire TIMEBOOST_net_14627;
wire TIMEBOOST_net_23026;
wire TIMEBOOST_net_20935;
wire g66424_db;
wire g66425_db;
wire TIMEBOOST_net_22294;
wire g66426_db;
wire g66427_db;
wire g66428_db;
wire g66429_db;
wire TIMEBOOST_net_13365;
wire g66430_db;
wire TIMEBOOST_net_14281;
wire g66433_db;
wire g66433_sb;
wire TIMEBOOST_net_17126;
wire g66456_db;
wire g66456_sb;
wire g66457_sb;
wire g66458_p;
wire g66458_p0;
wire g66459_p0;
wire g66464_p;
wire g66464_p0;
wire g66465_p;
wire g66465_p0;
wire g66473_p;
wire g66475_p;
wire g66544_p;
wire g66547_p;
wire g66550_p;
wire g66577_p;
wire g66583_p;
wire g66584_p;
wire g66607_p;
wire g66620_p;
wire g66627_p;
wire g66628_p;
wire g66646_p;
wire g66649_p;
wire g66650_p;
wire g66652_p;
wire g66658_p;
wire g66662_p;
wire g66663_p;
wire g66669_p;
wire g66672_p;
wire g66714_p;
wire g66726_p;
wire g66728_p;
wire g66737_p;
wire g66738_p;
wire g66742_p;
wire g66752_p;
wire g66753_p;
wire g66759_p;
wire g66773_p;
wire g66777_p;
wire g66789_p;
wire g66805_p;
wire g66813_p;
wire g66825_p;
wire g66827_p;
wire g66854_p;
wire g66856_p;
wire g66866_p;
wire g66875_p;
wire g66876_p;
wire g66888_p;
wire g66889_p;
wire g66902_p;
wire g66911_p;
wire g66912_p;
wire g66913_p;
wire g66915_p;
wire g66917_p;
wire g66918_p;
wire g66921_p;
wire g66922_p;
wire g66923_p;
wire g66924_p;
wire g66925_p;
wire g66927_p;
wire g66929_p;
wire g66930_p;
wire g66931_p;
wire g66932_p;
wire g66933_p;
wire g66934_p;
wire g66935_p;
wire g66936_p;
wire g66937_p;
wire g66940_p;
wire g66941_p;
wire g66942_p;
wire g66944_p;
wire g66945_p;
wire g66946_p;
wire g66947_p;
wire g66948_p;
wire g66949_p;
wire g66951_p;
wire g66952_p;
wire g66953_p;
wire g66954_p;
wire g66955_p;
wire g66957_p;
wire g66959_p;
wire g66960_p;
wire g66963_p;
wire g66964_p;
wire g66965_p;
wire g66966_p;
wire g66968_p;
wire g66975_p;
wire g66978_p;
wire g66984_p;
wire g66985_p;
wire g66986_p;
wire g66987_p;
wire g66988_p;
wire g66989_p;
wire g66990_p;
wire g66997_p;
wire g67001_p;
wire g67003_p;
wire g67005_p;
wire g67006_p;
wire g67008_p;
wire g67010_p;
wire g67011_p;
wire g67014_p;
wire g67015_p;
wire g67017_p;
wire g67018_p;
wire g67019_p;
wire g67020_p;
wire g67021_p;
wire g67022_p;
wire g67023_p;
wire g67024_p;
wire g67025_p;
wire g67026_p;
wire g67029_p;
wire g67030_p;
wire g67031_p;
wire g67032_p;
wire g67033_p;
wire g67036_p;
wire TIMEBOOST_net_22483;
wire g67040_sb;
wire TIMEBOOST_net_100;
wire TIMEBOOST_net_7387;
wire TIMEBOOST_net_13992;
wire g67042_db;
wire g67042_sb;
wire TIMEBOOST_net_12;
wire g67043_db;
wire g67044_sb;
wire g67045_da;
wire TIMEBOOST_net_15533;
wire TIMEBOOST_net_16728;
wire g67046_sb;
wire g67048_sb;
wire g67049_db;
wire g67049_sb;
wire TIMEBOOST_net_7359;
wire g67050_db;
wire g67051_sb;
wire TIMEBOOST_net_10434;
wire TIMEBOOST_net_22907;
wire TIMEBOOST_net_22713;
wire TIMEBOOST_net_14521;
wire TIMEBOOST_net_14666;
wire TIMEBOOST_net_85;
wire TIMEBOOST_net_17450;
wire TIMEBOOST_net_21208;
wire TIMEBOOST_net_20439;
wire TIMEBOOST_net_21152;
wire TIMEBOOST_net_22342;
wire g67057_sb;
wire TIMEBOOST_net_43;
wire TIMEBOOST_net_14284;
wire TIMEBOOST_net_101;
wire TIMEBOOST_net_12685;
wire TIMEBOOST_net_22696;
wire TIMEBOOST_net_44;
wire TIMEBOOST_net_40;
wire TIMEBOOST_net_22707;
wire g67070_sb;
wire TIMEBOOST_net_86;
wire TIMEBOOST_net_21698;
wire TIMEBOOST_net_87;
wire TIMEBOOST_net_13676;
wire TIMEBOOST_net_35;
wire g67074_db;
wire g67075_db;
wire TIMEBOOST_net_21670;
wire TIMEBOOST_net_16689;
wire g67082_sb;
wire g67083_db;
wire TIMEBOOST_net_88;
wire g67085_db;
wire TIMEBOOST_net_41;
wire TIMEBOOST_net_89;
wire TIMEBOOST_net_13681;
wire TIMEBOOST_net_102;
wire TIMEBOOST_net_46;
wire TIMEBOOST_net_9769;
wire TIMEBOOST_net_14282;
wire TIMEBOOST_net_16691;
wire TIMEBOOST_net_47;
wire g67095_p;
wire g67096_p;
wire g67097_p;
wire g67098_p;
wire g67099_p;
wire g67100_p;
wire g67102_p;
wire g67103_p;
wire g67104_p;
wire g67105_p;
wire g67106_p;
wire g67107_p;
wire g67108_p;
wire g67109_p;
wire g67110_p;
wire g67111_p;
wire g67112_p;
wire g67113_p;
wire g67114_p;
wire g67115_p;
wire g67116_p;
wire g67117_p;
wire g67118_p;
wire g67119_p;
wire g67120_p;
wire g67122_p;
wire g67123_p;
wire g67125_p;
wire g67126_p;
wire g67127_p;
wire g67128_p;
wire g67129_p;
wire g67130_p;
wire g67131_p;
wire g67132_p;
wire g67133_p;
wire g67134_p;
wire g67135_p;
wire g67136_p;
wire g67138_p;
wire g67139_p;
wire g67140_p;
wire g67141_p;
wire g67142_p;
wire g67143_p;
wire TIMEBOOST_net_22582;
wire g67145_p;
wire g67146_p;
wire g67148_p;
wire g67149_p;
wire g67150_p;
wire g67151_p;
wire g67152_p;
wire g67153_p;
wire g67154_p;
wire g67155_p;
wire g67156_p;
wire g67157_p;
wire g67311_p;
wire g67313_p;
wire g67324_p;
wire g67327_p;
wire g67329_p;
wire g67340_p;
wire g67353_p;
wire g67355_p;
wire g67360_p;
wire g67364_p;
wire g67369_p;
wire g67371_p;
wire g67386_p;
wire g67389_p;
wire g67390_p;
wire g67392_p;
wire g67394_p;
wire g67396_p;
wire g67397_p;
wire g67403_p;
wire g67405_p;
wire g67411_p;
wire g67421_p;
wire g67425_p;
wire g67430_p;
wire g67432_p;
wire g67434_p;
wire g67437_p;
wire g67446_p;
wire g67453_p;
wire g67457_p;
wire g67459_p;
wire g67463_p;
wire g67468_p;
wire g67489_p;
wire g67493_p;
wire g67495_p;
wire g67498_p;
wire g67502_p;
wire g67505_p;
wire g67506_p;
wire g67507_p;
wire g67514_p;
wire g67519_p;
wire g67523_p;
wire g67531_p;
wire g67534_p;
wire g67535_p;
wire g67536_p;
wire g67537_p;
wire g67538_p;
wire g67544_p;
wire g67545_p;
wire g67549_p;
wire g67559_p;
wire g67581_p;
wire g67582_p;
wire g67583_p;
wire g67592_p;
wire g67596_p;
wire g67600_p;
wire g67603_p;
wire g67605_p;
wire g67610_p;
wire g67613_p;
wire g67624_p;
wire g67625_p;
wire g67626_p;
wire g67631_p;
wire g67671_p;
wire g67672_p;
wire g67675_p;
wire g67680_p;
wire g67688_p;
wire g67689_p;
wire g67699_p;
wire g67707_p;
wire g67709_p;
wire g67712_p;
wire g67721_p;
wire g67722_p;
wire g67725_p;
wire g67731_p;
wire g67735_p;
wire g67739_p;
wire g67745_p;
wire g67746_p;
wire g67747_p;
wire g67754_p;
wire g67757_p;
wire g67758_p;
wire g67763_p;
wire g67765_p;
wire g67778_p;
wire g67783_p;
wire g67791_p;
wire g67799_p;
wire g67802_p;
wire g67804_p;
wire g67806_p;
wire g67807_p;
wire g67814_p;
wire g67828_p;
wire g68_p;
wire g70_p;
wire g73989_p;
wire g74028_p;
wire g74140_p;
wire g74153_p;
wire g74154_p;
wire g74162_dup_p;
wire g74174_p;
wire g74243_p;
wire g74245_p;
wire g74270_p;
wire g74283_p;
wire g74363_p;
wire g74408_p;
wire g74429_p;
wire g74434_sb;
wire g74470_p;
wire g74475_p;
wire g74553_p;
wire g74563_p;
wire g74576_p;
wire g74580_p;
wire g74628_p;
wire g74644_p;
wire g74660_p;
wire g74661_p;
wire g74689_p;
wire g74739_p;
wire g74749_p;
wire g74787_p;
wire g74859_p;
wire g74872_p;
wire g74879_p;
wire g74886_p;
wire g74920_p;
wire g74930_p;
wire g74961_p;
wire g74967_p;
wire g74981_p;
wire g74996_p;
wire g75024_sb;
wire g75059_p;
wire g75061_p;
wire g75067_p;
wire TIMEBOOST_net_15815;
wire g75072_db;
wire g75072_sb;
wire g75081_p;
wire g75084_p;
wire g75088_p;
wire g75126_p;
wire TIMEBOOST_net_17247;
wire g75160_db;
wire g75160_sb;
wire g75162_db;
wire g75162_sb;
wire g75165_p;
wire g75174_p;
wire TIMEBOOST_net_15062;
wire g75181_db;
wire g75200_p;
wire g75332_p;
wire g75413_db;
wire TIMEBOOST_net_21306;
wire g75416_db;
wire g75418_da;
wire g75418_db;
wire g75_p;
wire i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q;
wire i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid;
wire n_0;
wire n_10002;
wire n_10007;
wire n_10010;
wire n_10014;
wire n_10017;
wire n_10020;
wire n_10023;
wire n_10026;
wire n_10029;
wire n_10032;
wire n_10035;
wire n_10038;
wire n_1004;
wire n_10041;
wire n_10048;
wire n_1005;
wire n_10051;
wire n_10054;
wire n_10057;
wire n_10060;
wire n_10063;
wire n_10066;
wire n_10069;
wire n_1007;
wire n_10075;
wire n_10078;
wire n_1008;
wire n_10081;
wire n_10084;
wire n_10087;
wire n_1009;
wire n_10090;
wire n_10093;
wire n_10096;
wire n_10099;
wire n_10102;
wire n_10105;
wire n_10106;
wire n_10109;
wire n_1011;
wire n_10112;
wire n_10116;
wire n_1012;
wire n_10120;
wire n_10124;
wire n_10127;
wire n_1013;
wire n_10131;
wire n_10134;
wire TIMEBOOST_net_16772;
wire TIMEBOOST_net_16774;
wire n_1014;
wire n_10141;
wire n_10143;
wire n_10144;
wire n_10147;
wire TIMEBOOST_net_15440;
wire n_1015;
wire n_10151;
wire n_10154;
wire n_10155;
wire n_10157;
wire n_1016;
wire n_10160;
wire n_10163;
wire TIMEBOOST_net_23546;
wire n_1017;
wire n_10170;
wire n_10173;
wire n_10176;
wire n_10179;
wire n_10183;
wire n_10185;
wire n_10188;
wire n_1019;
wire n_10193;
wire n_10195;
wire n_10198;
wire TIMEBOOST_net_16779;
wire n_10202;
wire n_10205;
wire n_10216;
wire n_10221;
wire n_1023;
wire n_10230;
wire n_10232;
wire n_10235;
wire n_10244;
wire n_10252;
wire n_10254;
wire n_10256;
wire TIMEBOOST_net_16778;
wire n_10258;
wire n_10259;
wire n_10261;
wire n_10268;
wire n_1027;
wire n_10270;
wire TIMEBOOST_net_17061;
wire n_10273;
wire TIMEBOOST_net_16773;
wire n_1028;
wire n_10281;
wire n_10285;
wire n_10286;
wire n_10288;
wire n_10289;
wire n_10290;
wire n_10291;
wire n_10292;
wire n_10294;
wire n_10296;
wire n_10297;
wire n_10298;
wire n_10300;
wire n_10302;
wire n_10304;
wire n_10306;
wire n_10308;
wire n_1031;
wire n_10310;
wire n_10311;
wire n_10312;
wire n_10314;
wire n_10316;
wire n_10317;
wire n_10319;
wire n_10321;
wire n_10323;
wire n_10325;
wire n_10327;
wire n_10329;
wire n_1033;
wire n_10331;
wire n_10332;
wire n_10334;
wire n_10336;
wire n_10338;
wire n_1034;
wire n_10340;
wire n_10342;
wire n_10343;
wire n_10344;
wire n_10346;
wire n_10348;
wire n_10349;
wire n_1035;
wire n_10351;
wire n_10353;
wire n_10355;
wire n_10357;
wire n_10359;
wire n_1036;
wire n_10361;
wire n_10362;
wire n_10363;
wire n_10365;
wire n_10366;
wire n_10368;
wire n_1037;
wire n_10370;
wire n_10372;
wire n_10374;
wire n_10376;
wire n_10377;
wire n_10378;
wire n_1038;
wire n_10380;
wire n_10381;
wire n_10383;
wire n_10384;
wire n_10385;
wire n_10386;
wire n_10388;
wire n_1039;
wire n_10390;
wire n_10391;
wire n_10393;
wire n_10394;
wire n_10396;
wire n_10397;
wire n_10399;
wire n_104;
wire n_10400;
wire n_10401;
wire n_10402;
wire n_10404;
wire n_10405;
wire n_10407;
wire n_10408;
wire n_1041;
wire n_10410;
wire n_10411;
wire n_10412;
wire n_10413;
wire n_10414;
wire n_10416;
wire n_10417;
wire n_10418;
wire n_10419;
wire n_10421;
wire n_10423;
wire n_10424;
wire n_10426;
wire n_10428;
wire n_10430;
wire n_10432;
wire n_10433;
wire n_10434;
wire n_10436;
wire n_10438;
wire n_10439;
wire n_10440;
wire n_10441;
wire n_10443;
wire n_10444;
wire n_10445;
wire n_10446;
wire n_10447;
wire n_10449;
wire n_10450;
wire n_10451;
wire n_10453;
wire n_10455;
wire n_10457;
wire n_10459;
wire n_10460;
wire n_10462;
wire n_10463;
wire n_10464;
wire n_10465;
wire n_10467;
wire n_10469;
wire n_10470;
wire n_10473;
wire n_10474;
wire n_10476;
wire n_10477;
wire n_10478;
wire n_10479;
wire n_10481;
wire n_10483;
wire n_10485;
wire n_10487;
wire n_10489;
wire n_10491;
wire n_10493;
wire n_10495;
wire n_10497;
wire n_10499;
wire n_10501;
wire n_10503;
wire n_10506;
wire n_10508;
wire n_10509;
wire n_10511;
wire n_10513;
wire n_10515;
wire n_10518;
wire n_10521;
wire n_10524;
wire n_10527;
wire n_10530;
wire n_10533;
wire n_10541;
wire n_10544;
wire n_10547;
wire n_10553;
wire n_10554;
wire n_10556;
wire n_10559;
wire n_10560;
wire n_10561;
wire n_10564;
wire n_10566;
wire n_10569;
wire n_1057;
wire n_10572;
wire n_10575;
wire n_10576;
wire n_10577;
wire n_10579;
wire n_10584;
wire n_10588;
wire n_10592;
wire n_10595;
wire n_10596;
wire n_10599;
wire n_10602;
wire n_10605;
wire n_10608;
wire n_1061;
wire n_10611;
wire n_10614;
wire n_10617;
wire n_10622;
wire n_10624;
wire n_10627;
wire n_10630;
wire n_10631;
wire n_10634;
wire n_10637;
wire n_10638;
wire n_1064;
wire n_10641;
wire n_10644;
wire n_10647;
wire n_10650;
wire n_10653;
wire n_10656;
wire n_10659;
wire n_10660;
wire n_10661;
wire n_10662;
wire n_10669;
wire n_10672;
wire n_10675;
wire n_10676;
wire n_10679;
wire n_10680;
wire n_10681;
wire n_10682;
wire n_10685;
wire n_10688;
wire n_1069;
wire n_10691;
wire n_10693;
wire n_10696;
wire n_10699;
wire n_10702;
wire n_10705;
wire n_10708;
wire n_10711;
wire n_10715;
wire n_1072;
wire n_10728;
wire n_1073;
wire n_10731;
wire n_10734;
wire n_10738;
wire n_1074;
wire n_10741;
wire n_10744;
wire n_10747;
wire n_10750;
wire n_10753;
wire n_10754;
wire n_10755;
wire n_10758;
wire n_10763;
wire n_10764;
wire n_10765;
wire n_10768;
wire n_1077;
wire n_10771;
wire n_10774;
wire n_10777;
wire n_10780;
wire n_10781;
wire n_10782;
wire n_10784;
wire n_10785;
wire n_10787;
wire n_10788;
wire n_10789;
wire n_1079;
wire n_10791;
wire n_10792;
wire n_10793;
wire n_10795;
wire n_10797;
wire n_10799;
wire n_1080;
wire n_10800;
wire n_10802;
wire n_10803;
wire n_10804;
wire n_10806;
wire n_10807;
wire n_1081;
wire n_10810;
wire n_10812;
wire n_10813;
wire n_10815;
wire n_10817;
wire n_10819;
wire n_10820;
wire n_10821;
wire n_10823;
wire n_10825;
wire n_10828;
wire n_10829;
wire n_1083;
wire n_10832;
wire n_10833;
wire n_10834;
wire n_10835;
wire n_10836;
wire n_10838;
wire n_10839;
wire n_1084;
wire n_10841;
wire n_10843;
wire n_10845;
wire n_10847;
wire n_10848;
wire n_1085;
wire n_10851;
wire n_10853;
wire n_10855;
wire n_10856;
wire n_10859;
wire n_1086;
wire n_10860;
wire n_10864;
wire n_10865;
wire n_10866;
wire n_10867;
wire n_10870;
wire n_10873;
wire n_10875;
wire n_10876;
wire n_10877;
wire n_1088;
wire n_10880;
wire n_10881;
wire n_10882;
wire n_10885;
wire n_10889;
wire n_1089;
wire n_10890;
wire n_10891;
wire n_10892;
wire n_10895;
wire n_10898;
wire n_10901;
wire n_10902;
wire n_10903;
wire n_10904;
wire n_10905;
wire n_10906;
wire n_10907;
wire n_10908;
wire n_10909;
wire n_1091;
wire n_10912;
wire n_10913;
wire n_10916;
wire n_10917;
wire n_10918;
wire n_10919;
wire n_10922;
wire n_10923;
wire n_10927;
wire n_1093;
wire n_10930;
wire n_10931;
wire n_10932;
wire n_10939;
wire n_1094;
wire n_10942;
wire n_10943;
wire n_10944;
wire n_10947;
wire n_1095;
wire n_10951;
wire n_10952;
wire n_10956;
wire n_1096;
wire n_10961;
wire n_10962;
wire n_10963;
wire n_10967;
wire n_10970;
wire n_10971;
wire n_10974;
wire n_10975;
wire n_10976;
wire n_10977;
wire n_10978;
wire n_1098;
wire n_10981;
wire n_10985;
wire n_10986;
wire n_10987;
wire n_1099;
wire n_10991;
wire n_10994;
wire n_11;
wire n_1100;
wire n_11002;
wire n_11005;
wire n_11008;
wire n_1101;
wire n_11013;
wire n_11014;
wire n_11019;
wire n_1103;
wire n_11034;
wire n_11036;
wire n_11037;
wire n_11038;
wire n_11039;
wire n_1104;
wire n_11040;
wire n_11041;
wire n_11042;
wire n_11043;
wire n_11044;
wire n_11046;
wire n_11047;
wire n_11048;
wire n_11049;
wire n_1105;
wire n_11050;
wire n_11051;
wire n_11053;
wire n_11054;
wire n_11055;
wire n_11056;
wire n_11057;
wire n_11058;
wire n_11059;
wire n_1106;
wire n_11060;
wire n_11061;
wire n_11062;
wire n_11063;
wire n_11064;
wire n_11065;
wire n_11066;
wire n_11067;
wire n_11069;
wire n_1107;
wire n_11070;
wire n_11071;
wire n_11072;
wire n_11073;
wire n_11075;
wire n_11076;
wire n_11077;
wire n_11078;
wire n_11079;
wire n_1108;
wire n_11081;
wire n_11083;
wire n_11084;
wire n_11085;
wire n_11086;
wire n_11087;
wire n_11088;
wire n_11089;
wire n_1109;
wire n_11090;
wire n_11091;
wire n_11092;
wire n_11093;
wire n_11094;
wire n_11095;
wire n_11096;
wire n_11097;
wire n_11099;
wire n_1110;
wire n_11100;
wire n_11101;
wire n_11102;
wire n_11104;
wire n_11106;
wire n_11107;
wire n_11108;
wire n_11109;
wire n_1111;
wire n_11110;
wire n_11111;
wire n_11113;
wire n_11115;
wire n_11118;
wire n_11119;
wire n_1112;
wire n_11120;
wire n_11121;
wire n_11122;
wire n_11123;
wire n_11124;
wire n_11125;
wire n_11126;
wire n_11129;
wire n_1113;
wire n_11130;
wire n_11131;
wire n_11132;
wire n_11134;
wire n_11135;
wire n_11136;
wire n_11137;
wire n_11138;
wire n_11139;
wire n_11140;
wire n_11142;
wire n_11143;
wire n_11144;
wire n_11145;
wire n_11146;
wire n_11147;
wire n_11148;
wire n_11149;
wire n_1115;
wire n_11152;
wire n_11153;
wire n_11155;
wire n_11157;
wire n_11158;
wire n_11159;
wire n_1116;
wire n_11161;
wire n_11162;
wire n_11164;
wire n_11165;
wire n_11167;
wire n_11169;
wire n_1117;
wire n_11171;
wire n_11173;
wire n_11174;
wire n_11175;
wire n_11177;
wire n_11178;
wire n_11179;
wire n_1118;
wire n_11180;
wire n_11181;
wire n_11182;
wire n_11184;
wire n_11186;
wire n_11187;
wire n_11188;
wire n_1119;
wire n_11190;
wire n_11191;
wire n_11193;
wire n_11194;
wire n_11196;
wire n_11198;
wire n_112;
wire n_1120;
wire n_11200;
wire n_11202;
wire n_11203;
wire n_11205;
wire n_11206;
wire n_11207;
wire n_11208;
wire n_11209;
wire n_11211;
wire n_11212;
wire n_11213;
wire n_11214;
wire n_11215;
wire n_11216;
wire n_11217;
wire n_11218;
wire n_11219;
wire n_1122;
wire n_11220;
wire n_11222;
wire n_11223;
wire n_11224;
wire n_11226;
wire n_11228;
wire n_11229;
wire n_1123;
wire n_11230;
wire n_11232;
wire n_11234;
wire n_11235;
wire n_11236;
wire n_11238;
wire n_11239;
wire n_1124;
wire n_11240;
wire n_11241;
wire n_11242;
wire n_11243;
wire n_11244;
wire n_11245;
wire n_11246;
wire n_11247;
wire n_11249;
wire n_1125;
wire n_11250;
wire n_11251;
wire n_11252;
wire n_11254;
wire n_11255;
wire n_11256;
wire n_11258;
wire n_11259;
wire n_1126;
wire n_11260;
wire n_11261;
wire n_11262;
wire n_11264;
wire n_11265;
wire n_11266;
wire n_11268;
wire n_11270;
wire n_11271;
wire n_11273;
wire n_11274;
wire n_11276;
wire n_11277;
wire n_11279;
wire n_11280;
wire n_11281;
wire n_11282;
wire n_11283;
wire n_11284;
wire n_11285;
wire n_11286;
wire n_11287;
wire n_11289;
wire n_11290;
wire n_11293;
wire n_11295;
wire n_11297;
wire n_11300;
wire n_11302;
wire n_11303;
wire n_11305;
wire n_11306;
wire n_11307;
wire n_11309;
wire n_11311;
wire n_11314;
wire n_11316;
wire n_11318;
wire n_11320;
wire n_11322;
wire n_11324;
wire n_11326;
wire n_11327;
wire n_11328;
wire n_1133;
wire n_11330;
wire n_11332;
wire n_11334;
wire n_11336;
wire n_11337;
wire n_11338;
wire n_1134;
wire n_11340;
wire n_11342;
wire n_11344;
wire n_11345;
wire n_11347;
wire n_11349;
wire n_11350;
wire n_11352;
wire n_11353;
wire n_11355;
wire n_11357;
wire n_11359;
wire n_11361;
wire n_11362;
wire n_11363;
wire n_11365;
wire n_11367;
wire n_11369;
wire n_11370;
wire n_11372;
wire n_11373;
wire n_11375;
wire n_11377;
wire n_11379;
wire n_11380;
wire n_11381;
wire n_11382;
wire n_11383;
wire n_11384;
wire n_11385;
wire n_11386;
wire n_11388;
wire n_11390;
wire n_11391;
wire n_11393;
wire n_11394;
wire n_11396;
wire n_11398;
wire n_11399;
wire n_11401;
wire n_11402;
wire n_11403;
wire n_11405;
wire n_11406;
wire n_11408;
wire n_11410;
wire n_11411;
wire n_11413;
wire n_11414;
wire n_11415;
wire n_11417;
wire n_11418;
wire n_11419;
wire n_11420;
wire n_11421;
wire n_11423;
wire n_11424;
wire n_11425;
wire n_11427;
wire n_11429;
wire n_11431;
wire n_11432;
wire n_11433;
wire n_11434;
wire n_11435;
wire n_11436;
wire n_11437;
wire n_11438;
wire n_11440;
wire n_11441;
wire n_11442;
wire n_11443;
wire n_11445;
wire n_11446;
wire n_11448;
wire n_11449;
wire n_11450;
wire n_11451;
wire n_11452;
wire n_11454;
wire n_11456;
wire n_11457;
wire n_11458;
wire n_11460;
wire n_11462;
wire n_11463;
wire n_11464;
wire n_11466;
wire n_11467;
wire n_11468;
wire n_11470;
wire n_11472;
wire n_11473;
wire n_11474;
wire n_11476;
wire n_11477;
wire n_11478;
wire n_11479;
wire n_11480;
wire n_11482;
wire n_11483;
wire n_11484;
wire n_11485;
wire n_11487;
wire n_11489;
wire n_11490;
wire n_11492;
wire n_11493;
wire n_11495;
wire n_11496;
wire n_11497;
wire n_11499;
wire n_11500;
wire n_11502;
wire n_11503;
wire n_11505;
wire n_11507;
wire n_11509;
wire n_11510;
wire n_11512;
wire n_11513;
wire n_11515;
wire n_11516;
wire n_11517;
wire n_11519;
wire n_11521;
wire n_11523;
wire n_11524;
wire n_11526;
wire n_11528;
wire n_11530;
wire n_11531;
wire n_11532;
wire n_11533;
wire n_11534;
wire n_11535;
wire n_11536;
wire n_11538;
wire n_11540;
wire n_11542;
wire n_11543;
wire n_11544;
wire n_11545;
wire n_11546;
wire n_11547;
wire n_11548;
wire n_11549;
wire n_11551;
wire n_11553;
wire n_11555;
wire n_11556;
wire n_11557;
wire n_11559;
wire n_11560;
wire n_11561;
wire n_11562;
wire n_11564;
wire n_11565;
wire n_11566;
wire n_11568;
wire n_11570;
wire n_11571;
wire n_11572;
wire n_11573;
wire n_11575;
wire n_11577;
wire n_11579;
wire n_11580;
wire n_11582;
wire n_11583;
wire n_11584;
wire n_11585;
wire n_11586;
wire n_11587;
wire n_11588;
wire n_11589;
wire n_1159;
wire n_11590;
wire n_11592;
wire n_11593;
wire n_11595;
wire n_11597;
wire n_11598;
wire n_11599;
wire n_1160;
wire n_11600;
wire n_11601;
wire n_11602;
wire n_11603;
wire n_11604;
wire n_11605;
wire n_11606;
wire n_11607;
wire n_11609;
wire n_1161;
wire n_11610;
wire n_11611;
wire n_11613;
wire n_11614;
wire n_11616;
wire n_11617;
wire n_11618;
wire n_1162;
wire n_11620;
wire n_11622;
wire n_11623;
wire n_11624;
wire n_11625;
wire n_11626;
wire n_11628;
wire n_11630;
wire n_11631;
wire n_11632;
wire n_11633;
wire n_11634;
wire n_11635;
wire n_11637;
wire n_11638;
wire n_11639;
wire n_1164;
wire n_11640;
wire n_11641;
wire n_11642;
wire n_11644;
wire n_11645;
wire n_11647;
wire n_11648;
wire n_1165;
wire n_11650;
wire n_11651;
wire n_11652;
wire n_11653;
wire n_11655;
wire n_11657;
wire n_11659;
wire n_1166;
wire n_11660;
wire n_11661;
wire n_11662;
wire n_11663;
wire n_11665;
wire n_11666;
wire n_11667;
wire n_11668;
wire n_11669;
wire n_1167;
wire n_11670;
wire n_11671;
wire n_11672;
wire n_11674;
wire n_11675;
wire n_11676;
wire n_11677;
wire n_11679;
wire n_1168;
wire n_11680;
wire n_11681;
wire n_11682;
wire n_11683;
wire n_11684;
wire n_11685;
wire n_11686;
wire n_11687;
wire n_11688;
wire n_11689;
wire n_1169;
wire n_11690;
wire n_11691;
wire n_11692;
wire n_11693;
wire n_11694;
wire n_11695;
wire n_11696;
wire n_11697;
wire n_11698;
wire n_11699;
wire n_1170;
wire n_11700;
wire n_11701;
wire n_11702;
wire n_11703;
wire n_11705;
wire n_11706;
wire n_11707;
wire n_11708;
wire n_11710;
wire n_11712;
wire n_11715;
wire n_11716;
wire n_11717;
wire n_11718;
wire n_11719;
wire n_11720;
wire n_11723;
wire n_11724;
wire n_11725;
wire n_11726;
wire n_11727;
wire n_11728;
wire n_1173;
wire n_11730;
wire n_11731;
wire n_11732;
wire n_11733;
wire n_11734;
wire n_11735;
wire n_11736;
wire n_11738;
wire n_11739;
wire n_1174;
wire n_11740;
wire n_11741;
wire n_1175;
wire n_1176;
wire n_11762;
wire n_11767;
wire n_1177;
wire n_11773;
wire n_11774;
wire n_11775;
wire n_11776;
wire n_11777;
wire n_11778;
wire n_1178;
wire n_11780;
wire n_11781;
wire n_11782;
wire n_11783;
wire n_11784;
wire n_11786;
wire n_11788;
wire n_11790;
wire n_11791;
wire n_11792;
wire n_11793;
wire n_11795;
wire n_11796;
wire TIMEBOOST_net_21207;
wire n_1180;
wire TIMEBOOST_net_21206;
wire TIMEBOOST_net_12775;
wire TIMEBOOST_net_13316;
wire n_11805;
wire n_11806;
wire TIMEBOOST_net_13783;
wire TIMEBOOST_net_23311;
wire n_11814;
wire TIMEBOOST_net_14548;
wire n_11818;
wire n_11819;
wire TIMEBOOST_net_16295;
wire n_11823;
wire TIMEBOOST_net_23316;
wire TIMEBOOST_net_21515;
wire TIMEBOOST_net_12763;
wire n_1183;
wire TIMEBOOST_net_17320;
wire n_11831;
wire TIMEBOOST_net_23412;
wire TIMEBOOST_net_23336;
wire TIMEBOOST_net_12757;
wire TIMEBOOST_net_22354;
wire n_11841;
wire TIMEBOOST_net_12606;
wire n_11844;
wire n_11845;
wire n_11846;
wire n_11847;
wire n_11848;
wire n_11849;
wire n_1185;
wire n_11850;
wire n_11851;
wire n_11852;
wire n_11853;
wire n_11854;
wire n_11855;
wire n_11856;
wire n_11857;
wire n_11858;
wire n_11859;
wire n_1186;
wire n_11860;
wire n_11861;
wire n_11862;
wire n_11863;
wire n_11864;
wire n_11865;
wire n_11866;
wire n_11867;
wire n_11868;
wire n_11869;
wire n_1187;
wire n_11870;
wire n_11871;
wire n_11872;
wire n_11873;
wire n_11874;
wire n_11875;
wire n_11876;
wire n_11877;
wire n_11878;
wire n_1188;
wire n_11880;
wire n_11881;
wire n_11884;
wire n_11885;
wire n_11887;
wire TIMEBOOST_net_22009;
wire TIMEBOOST_net_21348;
wire n_1189;
wire TIMEBOOST_net_22086;
wire n_11891;
wire n_119;
wire n_1190;
wire TIMEBOOST_net_15158;
wire TIMEBOOST_net_23401;
wire n_11903;
wire TIMEBOOST_net_7027;
wire n_11908;
wire n_1191;
wire TIMEBOOST_net_20613;
wire TIMEBOOST_net_16165;
wire n_11912;
wire n_11913;
wire n_11914;
wire n_11915;
wire TIMEBOOST_net_23378;
wire TIMEBOOST_net_22041;
wire n_1192;
wire TIMEBOOST_net_21364;
wire TIMEBOOST_net_12787;
wire TIMEBOOST_net_21358;
wire TIMEBOOST_net_7283;
wire TIMEBOOST_net_21518;
wire TIMEBOOST_net_12786;
wire TIMEBOOST_net_16801;
wire n_1193;
wire TIMEBOOST_net_21724;
wire TIMEBOOST_net_13250;
wire TIMEBOOST_net_21189;
wire TIMEBOOST_net_20942;
wire TIMEBOOST_net_17372;
wire n_11937;
wire n_11938;
wire n_1194;
wire TIMEBOOST_net_16823;
wire TIMEBOOST_net_14911;
wire TIMEBOOST_net_17449;
wire TIMEBOOST_net_16814;
wire n_1195;
wire TIMEBOOST_net_21352;
wire TIMEBOOST_net_21343;
wire TIMEBOOST_net_23319;
wire TIMEBOOST_net_17511;
wire n_11956;
wire n_11957;
wire TIMEBOOST_net_14533;
wire n_1196;
wire n_11960;
wire n_11961;
wire n_11962;
wire n_11964;
wire TIMEBOOST_net_23502;
wire TIMEBOOST_net_12761;
wire TIMEBOOST_net_15152;
wire n_1197;
wire TIMEBOOST_net_15151;
wire TIMEBOOST_net_14301;
wire TIMEBOOST_net_15133;
wire n_11975;
wire n_11977;
wire n_1198;
wire TIMEBOOST_net_12774;
wire TIMEBOOST_net_21530;
wire n_1199;
wire n_11990;
wire n_11991;
wire n_11992;
wire TIMEBOOST_net_21540;
wire TIMEBOOST_net_10872;
wire TIMEBOOST_net_7275;
wire TIMEBOOST_net_15131;
wire n_12;
wire n_1200;
wire TIMEBOOST_net_11571;
wire n_12001;
wire n_12002;
wire n_12003;
wire n_12004;
wire TIMEBOOST_net_7143;
wire TIMEBOOST_net_15147;
wire TIMEBOOST_net_15293;
wire TIMEBOOST_net_20522;
wire n_1201;
wire n_12010;
wire TIMEBOOST_net_12593;
wire TIMEBOOST_net_17373;
wire TIMEBOOST_net_21386;
wire n_1202;
wire TIMEBOOST_net_15144;
wire TIMEBOOST_net_13782;
wire TIMEBOOST_net_21785;
wire n_12028;
wire TIMEBOOST_net_22104;
wire n_12031;
wire n_12032;
wire n_12036;
wire n_12037;
wire n_12038;
wire n_1204;
wire TIMEBOOST_net_17237;
wire TIMEBOOST_net_12613;
wire n_12044;
wire TIMEBOOST_net_23325;
wire n_12052;
wire n_12053;
wire n_12054;
wire n_12055;
wire TIMEBOOST_net_15142;
wire TIMEBOOST_net_21510;
wire TIMEBOOST_net_11642;
wire TIMEBOOST_net_21578;
wire n_12066;
wire TIMEBOOST_net_13048;
wire n_12068;
wire TIMEBOOST_net_20914;
wire n_1207;
wire TIMEBOOST_net_13047;
wire n_12072;
wire n_12073;
wire n_12075;
wire n_1208;
wire TIMEBOOST_net_22926;
wire n_12084;
wire TIMEBOOST_net_23333;
wire n_12088;
wire TIMEBOOST_net_13045;
wire n_1209;
wire TIMEBOOST_net_15847;
wire TIMEBOOST_net_13044;
wire TIMEBOOST_net_13043;
wire TIMEBOOST_net_22112;
wire n_12099;
wire n_1210;
wire TIMEBOOST_net_17508;
wire TIMEBOOST_net_22108;
wire n_12104;
wire TIMEBOOST_net_17507;
wire TIMEBOOST_net_13042;
wire TIMEBOOST_net_22109;
wire n_1211;
wire TIMEBOOST_net_21199;
wire n_12112;
wire TIMEBOOST_net_21418;
wire TIMEBOOST_net_23454;
wire TIMEBOOST_net_22316;
wire TIMEBOOST_net_22315;
wire n_12117;
wire TIMEBOOST_net_16834;
wire n_12122;
wire TIMEBOOST_net_20973;
wire TIMEBOOST_net_7313;
wire n_12128;
wire n_12129;
wire n_1213;
wire n_12130;
wire n_12132;
wire n_12133;
wire n_12134;
wire n_12135;
wire n_12137;
wire n_12139;
wire n_12140;
wire n_12141;
wire n_12143;
wire n_12144;
wire n_12145;
wire n_12146;
wire n_12147;
wire n_12148;
wire n_1215;
wire n_12151;
wire n_12153;
wire n_12154;
wire n_12155;
wire n_12156;
wire n_12158;
wire n_12159;
wire n_1216;
wire n_12160;
wire n_12161;
wire n_12162;
wire n_12163;
wire n_12164;
wire n_12165;
wire n_12166;
wire n_12167;
wire n_12168;
wire n_12169;
wire n_1217;
wire n_12170;
wire n_12179;
wire n_1218;
wire TIMEBOOST_net_22312;
wire TIMEBOOST_net_21549;
wire TIMEBOOST_net_16800;
wire n_12186;
wire TIMEBOOST_net_16826;
wire n_1219;
wire TIMEBOOST_net_23361;
wire TIMEBOOST_net_7162;
wire TIMEBOOST_net_13317;
wire TIMEBOOST_net_15101;
wire n_12195;
wire n_12196;
wire TIMEBOOST_net_22639;
wire n_1220;
wire TIMEBOOST_net_7160;
wire TIMEBOOST_net_7159;
wire TIMEBOOST_net_16806;
wire n_12203;
wire TIMEBOOST_net_21546;
wire TIMEBOOST_net_16825;
wire n_12206;
wire TIMEBOOST_net_7158;
wire TIMEBOOST_net_16805;
wire n_1221;
wire TIMEBOOST_net_15128;
wire TIMEBOOST_net_16824;
wire n_12212;
wire TIMEBOOST_net_7157;
wire TIMEBOOST_net_7285;
wire TIMEBOOST_net_21509;
wire TIMEBOOST_net_7156;
wire TIMEBOOST_net_22120;
wire TIMEBOOST_net_12461;
wire TIMEBOOST_net_21491;
wire TIMEBOOST_net_22181;
wire TIMEBOOST_net_7154;
wire TIMEBOOST_net_15301;
wire TIMEBOOST_net_21490;
wire n_12228;
wire TIMEBOOST_net_16804;
wire TIMEBOOST_net_7153;
wire TIMEBOOST_net_13145;
wire TIMEBOOST_net_15124;
wire TIMEBOOST_net_22642;
wire TIMEBOOST_net_7152;
wire n_12238;
wire TIMEBOOST_net_7151;
wire n_1224;
wire TIMEBOOST_net_21525;
wire n_12243;
wire n_12244;
wire TIMEBOOST_net_7150;
wire n_12246;
wire n_12248;
wire n_1225;
wire TIMEBOOST_net_16813;
wire TIMEBOOST_net_14286;
wire TIMEBOOST_net_16822;
wire n_12257;
wire n_12258;
wire TIMEBOOST_net_20988;
wire n_1226;
wire TIMEBOOST_net_16821;
wire TIMEBOOST_net_7147;
wire n_12264;
wire n_12266;
wire TIMEBOOST_net_21709;
wire TIMEBOOST_net_22446;
wire n_1227;
wire n_12271;
wire TIMEBOOST_net_11529;
wire TIMEBOOST_net_7309;
wire n_12274;
wire n_12275;
wire n_12276;
wire TIMEBOOST_net_21494;
wire TIMEBOOST_net_12459;
wire n_1228;
wire n_12280;
wire TIMEBOOST_net_7274;
wire TIMEBOOST_net_21493;
wire TIMEBOOST_net_7164;
wire TIMEBOOST_net_21191;
wire n_1229;
wire TIMEBOOST_net_21487;
wire TIMEBOOST_net_15122;
wire n_12293;
wire n_12294;
wire TIMEBOOST_net_12460;
wire TIMEBOOST_net_21226;
wire n_123;
wire n_1230;
wire n_12300;
wire TIMEBOOST_net_7140;
wire TIMEBOOST_net_21521;
wire TIMEBOOST_net_15290;
wire TIMEBOOST_net_7139;
wire n_1231;
wire n_12310;
wire TIMEBOOST_net_21527;
wire n_12313;
wire TIMEBOOST_net_22103;
wire TIMEBOOST_net_14511;
wire TIMEBOOST_net_20527;
wire TIMEBOOST_net_16816;
wire TIMEBOOST_net_16799;
wire TIMEBOOST_net_16841;
wire TIMEBOOST_net_17513;
wire TIMEBOOST_net_12457;
wire TIMEBOOST_net_16803;
wire TIMEBOOST_net_16815;
wire TIMEBOOST_net_21450;
wire TIMEBOOST_net_21534;
wire TIMEBOOST_net_21524;
wire TIMEBOOST_net_17512;
wire TIMEBOOST_net_15236;
wire TIMEBOOST_net_7265;
wire TIMEBOOST_net_15235;
wire n_12341;
wire TIMEBOOST_net_22189;
wire TIMEBOOST_net_15234;
wire TIMEBOOST_net_16811;
wire n_12345;
wire TIMEBOOST_net_23230;
wire n_12349;
wire TIMEBOOST_net_13231;
wire TIMEBOOST_net_23339;
wire TIMEBOOST_net_15233;
wire TIMEBOOST_net_15232;
wire TIMEBOOST_net_15231;
wire n_12357;
wire TIMEBOOST_net_15230;
wire TIMEBOOST_net_23363;
wire n_12362;
wire TIMEBOOST_net_17329;
wire TIMEBOOST_net_21442;
wire TIMEBOOST_net_22253;
wire TIMEBOOST_net_22285;
wire TIMEBOOST_net_16579;
wire TIMEBOOST_net_17374;
wire TIMEBOOST_net_22284;
wire TIMEBOOST_net_7136;
wire TIMEBOOST_net_15228;
wire n_12378;
wire n_12379;
wire n_1238;
wire n_12381;
wire n_12382;
wire TIMEBOOST_net_15559;
wire TIMEBOOST_net_10660;
wire TIMEBOOST_net_15225;
wire TIMEBOOST_net_15224;
wire TIMEBOOST_net_21478;
wire n_12393;
wire TIMEBOOST_net_21728;
wire TIMEBOOST_net_21477;
wire TIMEBOOST_net_13732;
wire TIMEBOOST_net_14652;
wire n_1241;
wire TIMEBOOST_net_13016;
wire TIMEBOOST_net_15217;
wire n_12417;
wire TIMEBOOST_net_15215;
wire TIMEBOOST_net_15214;
wire n_12423;
wire TIMEBOOST_net_16836;
wire n_12425;
wire TIMEBOOST_net_16838;
wire TIMEBOOST_net_16835;
wire n_12429;
wire n_12430;
wire TIMEBOOST_net_16833;
wire TIMEBOOST_net_16832;
wire TIMEBOOST_net_16831;
wire n_12439;
wire n_12440;
wire n_12441;
wire n_12442;
wire TIMEBOOST_net_21991;
wire n_12447;
wire n_12448;
wire n_12449;
wire n_12450;
wire n_12451;
wire n_12452;
wire n_12453;
wire TIMEBOOST_net_23134;
wire n_12455;
wire n_12459;
wire TIMEBOOST_net_14258;
wire n_12461;
wire TIMEBOOST_net_12592;
wire TIMEBOOST_net_15226;
wire TIMEBOOST_net_15218;
wire TIMEBOOST_net_7259;
wire TIMEBOOST_net_16839;
wire n_12474;
wire n_12475;
wire n_12476;
wire n_12478;
wire n_12479;
wire n_1248;
wire n_12480;
wire n_12481;
wire n_12483;
wire n_12484;
wire n_12485;
wire n_12486;
wire n_12487;
wire n_12488;
wire n_12489;
wire n_12490;
wire n_12491;
wire n_12492;
wire n_12493;
wire n_12494;
wire n_12495;
wire n_12496;
wire n_12498;
wire n_12499;
wire n_12500;
wire n_12501;
wire n_12502;
wire n_12503;
wire n_12504;
wire n_12505;
wire n_12506;
wire n_12507;
wire n_12508;
wire n_12509;
wire n_1251;
wire n_12510;
wire n_12511;
wire n_12512;
wire n_12513;
wire n_12514;
wire n_12515;
wire n_12516;
wire n_12517;
wire n_12518;
wire n_12519;
wire n_1252;
wire n_12520;
wire n_12521;
wire n_12522;
wire n_12523;
wire n_12524;
wire n_12525;
wire n_12526;
wire n_12527;
wire n_12528;
wire n_12529;
wire n_1253;
wire n_12530;
wire n_12531;
wire n_12532;
wire n_12533;
wire n_12534;
wire n_12535;
wire n_12536;
wire n_12537;
wire n_12538;
wire n_12539;
wire n_12540;
wire n_12541;
wire n_12542;
wire n_12543;
wire n_12544;
wire n_12545;
wire n_12546;
wire n_12547;
wire n_12548;
wire n_12549;
wire n_12550;
wire n_12551;
wire n_12552;
wire n_12553;
wire n_12554;
wire n_12555;
wire n_12556;
wire n_12557;
wire n_12558;
wire n_12559;
wire n_12560;
wire n_12561;
wire n_12562;
wire n_12563;
wire n_12564;
wire n_12565;
wire n_12566;
wire n_12567;
wire n_12568;
wire n_12569;
wire n_12570;
wire n_12571;
wire n_12572;
wire n_12573;
wire n_12574;
wire n_12575;
wire n_12577;
wire n_12578;
wire n_12579;
wire n_1258;
wire n_12580;
wire n_12581;
wire n_12583;
wire n_12584;
wire n_12585;
wire n_12586;
wire n_12587;
wire n_12588;
wire n_12589;
wire n_1259;
wire n_12590;
wire n_12591;
wire n_12595;
wire n_12596;
wire n_12597;
wire n_12598;
wire n_12599;
wire n_1260;
wire n_12600;
wire n_12602;
wire n_12603;
wire n_12604;
wire n_12605;
wire n_12606;
wire n_12607;
wire n_1261;
wire n_12610;
wire n_12611;
wire n_12612;
wire n_12613;
wire n_12614;
wire n_12615;
wire n_12616;
wire n_12617;
wire n_12618;
wire n_12619;
wire n_12620;
wire n_12621;
wire n_12622;
wire n_12623;
wire n_12624;
wire n_12625;
wire n_12626;
wire n_12628;
wire n_12629;
wire n_1263;
wire n_12630;
wire n_12631;
wire n_12632;
wire n_12633;
wire n_12634;
wire n_12635;
wire n_12636;
wire n_12637;
wire n_12638;
wire n_12639;
wire n_1264;
wire n_12640;
wire n_12641;
wire n_12642;
wire n_12643;
wire n_12644;
wire n_12645;
wire n_12646;
wire n_12647;
wire n_12648;
wire n_12649;
wire n_1265;
wire n_12650;
wire n_12651;
wire n_12652;
wire n_12653;
wire n_12654;
wire n_12655;
wire n_12656;
wire n_12658;
wire n_12659;
wire n_1266;
wire n_12660;
wire n_12661;
wire n_12662;
wire n_12663;
wire n_12664;
wire n_12665;
wire n_12666;
wire n_12667;
wire n_12668;
wire n_12669;
wire n_12670;
wire n_12671;
wire n_12672;
wire n_12673;
wire n_12674;
wire n_12675;
wire n_12676;
wire n_12677;
wire n_12678;
wire n_12679;
wire n_12680;
wire n_12681;
wire n_12682;
wire n_12683;
wire n_12684;
wire n_12685;
wire n_12686;
wire n_12688;
wire n_12689;
wire n_1269;
wire n_12692;
wire n_12693;
wire n_12695;
wire n_12696;
wire n_12697;
wire n_12699;
wire n_1270;
wire n_12700;
wire n_12701;
wire n_12702;
wire n_12703;
wire n_12704;
wire n_12705;
wire n_12706;
wire n_12707;
wire n_12709;
wire n_12710;
wire n_12711;
wire n_12712;
wire n_12713;
wire n_12714;
wire n_12715;
wire n_12716;
wire n_12717;
wire n_1272;
wire n_12720;
wire n_12721;
wire n_12722;
wire n_12723;
wire n_12724;
wire n_12725;
wire n_12726;
wire n_12727;
wire n_12728;
wire n_12729;
wire n_1273;
wire n_12731;
wire n_12732;
wire n_12733;
wire n_12734;
wire n_12735;
wire n_12736;
wire n_12737;
wire n_12738;
wire n_1274;
wire n_12741;
wire n_12742;
wire n_12743;
wire n_12744;
wire n_12745;
wire n_12746;
wire n_12747;
wire n_12748;
wire n_12749;
wire n_1275;
wire n_12750;
wire n_12751;
wire n_12752;
wire n_12753;
wire n_12754;
wire n_12756;
wire n_12757;
wire n_12758;
wire n_12759;
wire n_1276;
wire n_12760;
wire n_12761;
wire n_12762;
wire n_12763;
wire n_12764;
wire n_12765;
wire n_12766;
wire n_12767;
wire n_12768;
wire n_12769;
wire n_1277;
wire n_12770;
wire n_12771;
wire n_12772;
wire n_12773;
wire n_12774;
wire n_12775;
wire n_12776;
wire n_12778;
wire n_12779;
wire n_12780;
wire n_12781;
wire n_12783;
wire n_12784;
wire n_12785;
wire n_12786;
wire n_12787;
wire n_12788;
wire n_12789;
wire n_1279;
wire n_12790;
wire n_12791;
wire n_12792;
wire n_12795;
wire n_12797;
wire n_12799;
wire n_1280;
wire n_12801;
wire n_12805;
wire n_12806;
wire n_12809;
wire n_1281;
wire n_12810;
wire n_12811;
wire n_12812;
wire n_12813;
wire n_12814;
wire n_12815;
wire n_12816;
wire n_12817;
wire n_12818;
wire n_12819;
wire n_1282;
wire n_12821;
wire n_12822;
wire n_12823;
wire n_12824;
wire n_12825;
wire n_12826;
wire n_12827;
wire n_12828;
wire n_12829;
wire n_1283;
wire n_12830;
wire n_12831;
wire n_12832;
wire n_12833;
wire n_12834;
wire n_12835;
wire n_12836;
wire n_12837;
wire n_12839;
wire n_12840;
wire n_12841;
wire n_12842;
wire n_12843;
wire n_12845;
wire n_12846;
wire n_12847;
wire n_12848;
wire n_12849;
wire n_1285;
wire n_12850;
wire n_12851;
wire n_12852;
wire n_12853;
wire n_12855;
wire n_12858;
wire n_12859;
wire n_1286;
wire n_12862;
wire n_12863;
wire n_12864;
wire n_12865;
wire n_12866;
wire n_12867;
wire n_12868;
wire n_12869;
wire n_1287;
wire n_12870;
wire n_12871;
wire n_12872;
wire n_12873;
wire n_12874;
wire n_12875;
wire n_12876;
wire n_12877;
wire n_12878;
wire n_12879;
wire n_1288;
wire n_12880;
wire n_12881;
wire n_12882;
wire n_12883;
wire n_12884;
wire n_12885;
wire n_12886;
wire n_12887;
wire n_12888;
wire n_12889;
wire n_1289;
wire n_12890;
wire n_12891;
wire n_12892;
wire n_12893;
wire n_12894;
wire n_12895;
wire n_12896;
wire n_12897;
wire n_12898;
wire n_12899;
wire n_1290;
wire n_12900;
wire n_12901;
wire n_12902;
wire n_12903;
wire n_12904;
wire n_12905;
wire n_12906;
wire n_12907;
wire n_12908;
wire n_1291;
wire n_12911;
wire n_12912;
wire n_12913;
wire n_12914;
wire n_12915;
wire n_12916;
wire n_12917;
wire n_12918;
wire n_12919;
wire n_12920;
wire n_12921;
wire n_12922;
wire n_12923;
wire n_12924;
wire n_12927;
wire n_12928;
wire n_12929;
wire n_1293;
wire n_12930;
wire n_12931;
wire n_12932;
wire n_12933;
wire n_12934;
wire n_12935;
wire n_12936;
wire n_12937;
wire n_12938;
wire n_12939;
wire n_1294;
wire n_12940;
wire n_12941;
wire n_12942;
wire n_12943;
wire n_12946;
wire n_12947;
wire n_12948;
wire n_12949;
wire n_12950;
wire n_12951;
wire n_12952;
wire n_12954;
wire n_12956;
wire n_12957;
wire n_12958;
wire n_12959;
wire n_12960;
wire n_12961;
wire n_12962;
wire n_12963;
wire n_12964;
wire n_12966;
wire n_12968;
wire n_12970;
wire n_12972;
wire n_12974;
wire n_12976;
wire n_12978;
wire n_12980;
wire n_12981;
wire n_12982;
wire n_12983;
wire n_12984;
wire n_12985;
wire n_12986;
wire n_12988;
wire n_1299;
wire n_12992;
wire n_12994;
wire TIMEBOOST_net_776;
wire n_12998;
wire TIMEBOOST_net_11408;
wire TIMEBOOST_net_22081;
wire TIMEBOOST_net_775;
wire TIMEBOOST_net_7413;
wire n_13012;
wire n_13018;
wire n_13020;
wire n_13022;
wire n_13026;
wire n_13027;
wire n_13028;
wire n_13034;
wire n_1304;
wire n_13041;
wire n_13042;
wire n_13043;
wire n_13044;
wire n_13045;
wire n_13046;
wire n_13047;
wire n_13048;
wire n_13049;
wire n_13050;
wire n_13051;
wire n_13052;
wire n_13053;
wire n_13054;
wire n_13055;
wire n_13056;
wire n_13057;
wire n_13058;
wire n_13059;
wire n_1306;
wire n_13060;
wire n_13061;
wire n_13063;
wire n_13064;
wire n_13065;
wire n_13066;
wire n_13067;
wire n_13068;
wire n_13073;
wire n_13074;
wire n_13075;
wire n_13076;
wire n_13077;
wire n_13078;
wire n_13079;
wire n_13080;
wire n_13081;
wire n_13082;
wire n_13083;
wire n_13084;
wire n_13085;
wire n_13086;
wire n_13087;
wire n_13088;
wire n_13089;
wire n_13090;
wire n_13091;
wire n_13093;
wire n_13094;
wire n_13095;
wire n_13097;
wire n_13098;
wire TIMEBOOST_net_21236;
wire n_13102;
wire g65775_db;
wire TIMEBOOST_net_17422;
wire TIMEBOOST_net_22155;
wire TIMEBOOST_net_11415;
wire TIMEBOOST_net_21641;
wire n_13116;
wire n_13117;
wire n_13118;
wire n_13120;
wire n_13122;
wire n_13123;
wire n_13124;
wire n_13125;
wire n_13127;
wire n_13128;
wire n_13129;
wire n_13130;
wire n_13131;
wire n_13132;
wire n_13133;
wire n_13134;
wire n_13135;
wire n_13136;
wire n_13137;
wire n_13138;
wire n_13139;
wire n_13140;
wire n_13141;
wire n_13142;
wire n_13143;
wire n_13144;
wire n_13145;
wire n_13146;
wire n_1315;
wire TIMEBOOST_net_23135;
wire n_1316;
wire TIMEBOOST_net_23133;
wire TIMEBOOST_net_22557;
wire TIMEBOOST_net_16248;
wire TIMEBOOST_net_22643;
wire n_13166;
wire n_13167;
wire n_13168;
wire TIMEBOOST_net_22534;
wire n_1317;
wire TIMEBOOST_net_22516;
wire n_2185;
wire g65698_db;
wire TIMEBOOST_net_17585;
wire n_13179;
wire n_1318;
wire n_13180;
wire TIMEBOOST_net_22548;
wire TIMEBOOST_net_14050;
wire n_13184;
wire TIMEBOOST_net_22622;
wire g65679_db;
wire TIMEBOOST_net_23409;
wire TIMEBOOST_net_11209;
wire TIMEBOOST_net_11208;
wire TIMEBOOST_net_16352;
wire TIMEBOOST_net_16347;
wire TIMEBOOST_net_11207;
wire TIMEBOOST_net_11206;
wire TIMEBOOST_net_16493;
wire TIMEBOOST_net_21173;
wire TIMEBOOST_net_11203;
wire TIMEBOOST_net_21316;
wire TIMEBOOST_net_17421;
wire TIMEBOOST_net_16492;
wire TIMEBOOST_net_11202;
wire TIMEBOOST_net_11511;
wire TIMEBOOST_net_16491;
wire TIMEBOOST_net_22151;
wire TIMEBOOST_net_16764;
wire TIMEBOOST_net_11510;
wire TIMEBOOST_net_11509;
wire n_1322;
wire n_13221;
wire TIMEBOOST_net_14052;
wire TIMEBOOST_net_21116;
wire TIMEBOOST_net_11189;
wire TIMEBOOST_net_11289;
wire n_13228;
wire n_1323;
wire TIMEBOOST_net_8003;
wire n_13249;
wire n_1325;
wire TIMEBOOST_net_21532;
wire TIMEBOOST_net_21734;
wire n_1326;
wire TIMEBOOST_net_22084;
wire TIMEBOOST_net_15364;
wire n_1327;
wire TIMEBOOST_net_21799;
wire n_13273;
wire TIMEBOOST_net_16846;
wire n_13286;
wire n_13287;
wire n_1329;
wire n_13290;
wire n_13291;
wire n_13292;
wire n_13295;
wire n_1330;
wire n_13302;
wire n_13303;
wire n_13304;
wire n_13305;
wire n_13306;
wire n_13308;
wire n_13309;
wire n_1331;
wire n_13310;
wire n_13311;
wire n_13313;
wire n_13314;
wire n_13315;
wire n_13317;
wire n_13318;
wire n_13319;
wire n_1332;
wire n_13320;
wire n_13321;
wire n_13323;
wire TIMEBOOST_net_11204;
wire n_13327;
wire n_13328;
wire n_13329;
wire n_1333;
wire n_13332;
wire n_13333;
wire n_13334;
wire n_13335;
wire n_13337;
wire n_13338;
wire n_13339;
wire n_1334;
wire n_13340;
wire n_13341;
wire n_13342;
wire TIMEBOOST_net_12373;
wire TIMEBOOST_net_14451;
wire n_13346;
wire n_13348;
wire n_13349;
wire n_1335;
wire n_13350;
wire n_13353;
wire n_13354;
wire n_13355;
wire TIMEBOOST_net_22358;
wire n_13357;
wire n_13358;
wire n_13359;
wire TIMEBOOST_net_7488;
wire n_13361;
wire TIMEBOOST_net_13685;
wire n_13363;
wire n_13365;
wire n_13366;
wire n_13367;
wire n_13368;
wire n_13369;
wire n_1337;
wire n_13370;
wire n_13371;
wire n_13372;
wire n_13373;
wire n_13374;
wire n_13375;
wire n_13376;
wire n_13377;
wire n_13378;
wire n_13379;
wire n_1338;
wire n_13380;
wire n_13381;
wire n_13383;
wire n_13384;
wire n_13386;
wire n_13387;
wire n_13388;
wire n_13389;
wire n_13390;
wire n_13391;
wire n_13392;
wire n_13393;
wire n_13394;
wire n_13395;
wire n_13398;
wire n_13399;
wire n_1340;
wire n_13400;
wire n_13401;
wire n_13402;
wire n_13403;
wire n_13404;
wire n_13405;
wire n_13406;
wire n_13407;
wire n_13408;
wire n_13409;
wire n_1341;
wire n_13410;
wire n_13411;
wire n_13412;
wire n_13414;
wire n_13415;
wire n_13416;
wire n_13417;
wire n_13418;
wire n_13419;
wire n_1342;
wire n_13420;
wire n_13421;
wire n_13422;
wire n_13423;
wire n_13424;
wire n_13425;
wire n_13426;
wire n_13427;
wire n_13428;
wire n_13429;
wire n_1343;
wire n_13430;
wire n_13431;
wire n_13432;
wire n_13434;
wire n_1344;
wire n_13441;
wire TIMEBOOST_net_17260;
wire n_13444;
wire n_13447;
wire n_13448;
wire n_1345;
wire n_13450;
wire TIMEBOOST_net_22412;
wire n_1346;
wire TIMEBOOST_net_21567;
wire n_13468;
wire n_13469;
wire n_1347;
wire n_13470;
wire n_13474;
wire n_13475;
wire n_13479;
wire n_13481;
wire n_13482;
wire n_13483;
wire n_13484;
wire n_13485;
wire n_13486;
wire n_13487;
wire n_13488;
wire TIMEBOOST_net_21417;
wire n_1349;
wire n_13490;
wire n_13491;
wire n_13493;
wire n_13494;
wire n_13495;
wire n_13496;
wire n_13497;
wire n_13499;
wire n_135;
wire n_1350;
wire n_13500;
wire n_13502;
wire n_13503;
wire n_13504;
wire n_13505;
wire n_13506;
wire n_13508;
wire n_13509;
wire n_1351;
wire n_13511;
wire n_13512;
wire n_13513;
wire n_13514;
wire n_13515;
wire n_13516;
wire n_13517;
wire n_13518;
wire n_13519;
wire n_1352;
wire n_13520;
wire n_13521;
wire n_13522;
wire n_13523;
wire n_13524;
wire n_13525;
wire n_13526;
wire n_13527;
wire n_13528;
wire n_13529;
wire n_1353;
wire n_13530;
wire n_13531;
wire n_13532;
wire n_13533;
wire n_13534;
wire n_13535;
wire n_13536;
wire n_13537;
wire n_13538;
wire n_13539;
wire n_1354;
wire n_13540;
wire n_13541;
wire n_13543;
wire n_13544;
wire n_13546;
wire n_13547;
wire n_13548;
wire n_1355;
wire n_13550;
wire n_13552;
wire n_13553;
wire n_13554;
wire n_13555;
wire n_13556;
wire n_13557;
wire n_13558;
wire n_13559;
wire n_1356;
wire n_13560;
wire n_13561;
wire n_13562;
wire n_13563;
wire n_13564;
wire n_13565;
wire n_13566;
wire TIMEBOOST_net_6912;
wire n_13568;
wire n_13569;
wire n_1357;
wire TIMEBOOST_net_16516;
wire n_13571;
wire n_13573;
wire n_13574;
wire n_13575;
wire n_13576;
wire n_13577;
wire n_13578;
wire n_13579;
wire n_1358;
wire n_13581;
wire n_13582;
wire n_13585;
wire n_13587;
wire n_1359;
wire n_13591;
wire n_13592;
wire n_13595;
wire n_13597;
wire n_13599;
wire n_13601;
wire n_13603;
wire n_13605;
wire n_13607;
wire n_13608;
wire n_13609;
wire n_1361;
wire n_13611;
wire n_13613;
wire n_13614;
wire n_13616;
wire n_13617;
wire n_13618;
wire n_13619;
wire n_1362;
wire n_13620;
wire n_13621;
wire n_13622;
wire n_13623;
wire n_13624;
wire n_13625;
wire n_13627;
wire n_13628;
wire n_13629;
wire n_1363;
wire n_13631;
wire n_13632;
wire n_13634;
wire n_13635;
wire n_13636;
wire n_13638;
wire n_13640;
wire n_13641;
wire n_13642;
wire n_13643;
wire n_13645;
wire n_13646;
wire n_13647;
wire n_13648;
wire n_1365;
wire n_13650;
wire n_13651;
wire TIMEBOOST_net_11217;
wire n_13653;
wire n_13654;
wire n_13657;
wire n_13658;
wire n_13659;
wire n_1366;
wire n_13661;
wire n_13662;
wire n_13663;
wire n_13664;
wire n_13666;
wire n_13667;
wire n_13668;
wire n_13670;
wire n_13671;
wire n_13672;
wire n_13673;
wire n_13674;
wire n_13678;
wire n_13679;
wire n_13680;
wire n_13681;
wire n_13682;
wire n_13685;
wire n_13686;
wire n_13687;
wire n_13688;
wire n_13689;
wire n_1369;
wire n_13691;
wire n_13692;
wire n_13693;
wire n_13694;
wire n_13695;
wire n_13696;
wire n_13697;
wire n_13698;
wire n_13701;
wire n_13703;
wire n_13704;
wire n_13705;
wire n_13709;
wire n_1371;
wire n_13710;
wire n_13711;
wire n_13712;
wire n_13715;
wire n_13716;
wire n_13717;
wire n_13719;
wire n_1372;
wire n_13720;
wire n_13721;
wire n_13722;
wire n_13724;
wire n_13725;
wire n_13727;
wire n_13728;
wire n_13729;
wire n_1373;
wire n_13731;
wire n_13732;
wire n_13734;
wire n_13735;
wire n_13736;
wire n_13738;
wire n_1374;
wire n_13740;
wire n_13741;
wire n_13743;
wire n_13744;
wire n_13745;
wire TIMEBOOST_net_10284;
wire n_13748;
wire n_13749;
wire n_13750;
wire n_13752;
wire n_13753;
wire n_13754;
wire n_13755;
wire n_13756;
wire n_13757;
wire n_13758;
wire n_13759;
wire n_13760;
wire n_13761;
wire TIMEBOOST_net_14272;
wire n_13763;
wire n_13764;
wire n_13765;
wire n_13766;
wire n_13767;
wire n_13768;
wire n_1377;
wire n_13770;
wire n_13771;
wire n_13772;
wire TIMEBOOST_net_22352;
wire n_13774;
wire n_13775;
wire n_13776;
wire TIMEBOOST_net_16726;
wire TIMEBOOST_net_6913;
wire n_1378;
wire n_13780;
wire n_13781;
wire n_13783;
wire n_13784;
wire n_13785;
wire n_13787;
wire n_13789;
wire n_1379;
wire n_13790;
wire n_13792;
wire n_13793;
wire n_13794;
wire n_13798;
wire n_13806;
wire n_13807;
wire n_13809;
wire n_1381;
wire n_13810;
wire n_13812;
wire n_13813;
wire n_13814;
wire n_13815;
wire n_13816;
wire n_13817;
wire n_13819;
wire n_1382;
wire n_13820;
wire n_13821;
wire n_13822;
wire n_13823;
wire n_13824;
wire n_13825;
wire n_13826;
wire n_13827;
wire n_13828;
wire n_13829;
wire n_1383;
wire n_13830;
wire n_13831;
wire n_1384;
wire n_13842;
wire n_13843;
wire n_13844;
wire TIMEBOOST_net_13894;
wire n_13846;
wire n_13847;
wire TIMEBOOST_net_12982;
wire n_13849;
wire n_1385;
wire TIMEBOOST_net_13232;
wire TIMEBOOST_net_23458;
wire TIMEBOOST_net_7241;
wire n_13854;
wire n_13856;
wire n_13857;
wire TIMEBOOST_net_13240;
wire n_13859;
wire n_13862;
wire TIMEBOOST_net_15434;
wire TIMEBOOST_net_21752;
wire TIMEBOOST_net_21702;
wire n_13868;
wire TIMEBOOST_net_14591;
wire n_1387;
wire TIMEBOOST_net_12898;
wire n_13873;
wire TIMEBOOST_net_21627;
wire TIMEBOOST_net_21742;
wire TIMEBOOST_net_11630;
wire n_1388;
wire TIMEBOOST_net_22075;
wire TIMEBOOST_net_12861;
wire TIMEBOOST_net_16926;
wire TIMEBOOST_net_16925;
wire TIMEBOOST_net_16924;
wire TIMEBOOST_net_21798;
wire TIMEBOOST_net_20442;
wire TIMEBOOST_net_21597;
wire n_1389;
wire n_13891;
wire TIMEBOOST_net_13389;
wire n_139;
wire n_1390;
wire n_13901;
wire n_13903;
wire TIMEBOOST_net_22011;
wire TIMEBOOST_net_21737;
wire n_13907;
wire n_13908;
wire n_1391;
wire n_13910;
wire n_13911;
wire n_13917;
wire n_13918;
wire n_13919;
wire n_1392;
wire n_13920;
wire n_13921;
wire n_13922;
wire n_13923;
wire TIMEBOOST_net_20252;
wire TIMEBOOST_net_23509;
wire n_1393;
wire n_13930;
wire TIMEBOOST_net_22001;
wire TIMEBOOST_net_14651;
wire TIMEBOOST_net_22069;
wire n_13937;
wire n_13938;
wire TIMEBOOST_net_16856;
wire n_1394;
wire TIMEBOOST_net_7219;
wire TIMEBOOST_net_13723;
wire TIMEBOOST_net_12904;
wire TIMEBOOST_net_20251;
wire TIMEBOOST_net_16855;
wire TIMEBOOST_net_17400;
wire TIMEBOOST_net_13230;
wire n_1395;
wire TIMEBOOST_net_21632;
wire TIMEBOOST_net_12903;
wire TIMEBOOST_net_16854;
wire TIMEBOOST_net_16820;
wire TIMEBOOST_net_16853;
wire TIMEBOOST_net_13238;
wire n_1396;
wire TIMEBOOST_net_13239;
wire TIMEBOOST_net_14463;
wire TIMEBOOST_net_16851;
wire TIMEBOOST_net_13236;
wire TIMEBOOST_net_16850;
wire TIMEBOOST_net_14604;
wire n_1397;
wire TIMEBOOST_net_12902;
wire n_13971;
wire n_13972;
wire TIMEBOOST_net_16849;
wire TIMEBOOST_net_23466;
wire TIMEBOOST_net_21601;
wire n_1398;
wire n_13980;
wire TIMEBOOST_net_17531;
wire n_13982;
wire TIMEBOOST_net_13185;
wire TIMEBOOST_net_16873;
wire TIMEBOOST_net_12374;
wire n_13987;
wire n_1399;
wire n_13990;
wire n_13991;
wire n_13993;
wire n_13995;
wire TIMEBOOST_net_13162;
wire n_13997;
wire n_13999;
wire n_14;
wire n_1400;
wire n_14000;
wire TIMEBOOST_net_21900;
wire TIMEBOOST_net_22060;
wire TIMEBOOST_net_16848;
wire n_1401;
wire n_14011;
wire TIMEBOOST_net_16847;
wire TIMEBOOST_net_14654;
wire g52461_da;
wire n_1402;
wire TIMEBOOST_net_7105;
wire TIMEBOOST_net_13161;
wire n_14022;
wire TIMEBOOST_net_21555;
wire TIMEBOOST_net_16842;
wire TIMEBOOST_net_15052;
wire TIMEBOOST_net_23531;
wire n_1403;
wire TIMEBOOST_net_16713;
wire TIMEBOOST_net_15876;
wire TIMEBOOST_net_21322;
wire TIMEBOOST_net_16058;
wire TIMEBOOST_net_20214;
wire TIMEBOOST_net_15524;
wire n_1404;
wire TIMEBOOST_net_10668;
wire TIMEBOOST_net_21373;
wire TIMEBOOST_net_21004;
wire TIMEBOOST_net_16673;
wire TIMEBOOST_net_13194;
wire TIMEBOOST_net_14649;
wire TIMEBOOST_net_16900;
wire n_1405;
wire g64980_db;
wire n_14054;
wire n_14055;
wire TIMEBOOST_net_13174;
wire n_1406;
wire g64314_db;
wire TIMEBOOST_net_13171;
wire TIMEBOOST_net_16684;
wire n_9013;
wire TIMEBOOST_net_23457;
wire n_1407;
wire n_14070;
wire n_14073;
wire n_14074;
wire n_14075;
wire n_14076;
wire n_14077;
wire n_14078;
wire n_14079;
wire n_1408;
wire n_14080;
wire n_14081;
wire n_14082;
wire n_14083;
wire n_14084;
wire n_14085;
wire n_14086;
wire n_14087;
wire n_14088;
wire n_1409;
wire n_14093;
wire n_14094;
wire TIMEBOOST_net_17538;
wire TIMEBOOST_net_21665;
wire n_14099;
wire n_1410;
wire n_14104;
wire TIMEBOOST_net_14655;
wire TIMEBOOST_net_20250;
wire n_1411;
wire n_14111;
wire TIMEBOOST_net_22165;
wire TIMEBOOST_net_16885;
wire TIMEBOOST_net_16884;
wire TIMEBOOST_net_7214;
wire TIMEBOOST_net_7213;
wire TIMEBOOST_net_7212;
wire n_1412;
wire TIMEBOOST_net_16881;
wire TIMEBOOST_net_7211;
wire TIMEBOOST_net_22326;
wire TIMEBOOST_net_13233;
wire TIMEBOOST_net_22479;
wire TIMEBOOST_net_7209;
wire TIMEBOOST_net_7208;
wire n_1413;
wire TIMEBOOST_net_7207;
wire TIMEBOOST_net_22716;
wire TIMEBOOST_net_16875;
wire g64324_db;
wire n_1414;
wire TIMEBOOST_net_22314;
wire n_14142;
wire n_14144;
wire n_1415;
wire TIMEBOOST_net_22267;
wire g52458_da;
wire g52473_da;
wire TIMEBOOST_net_17377;
wire TIMEBOOST_net_16868;
wire n_1416;
wire TIMEBOOST_net_16867;
wire n_14163;
wire TIMEBOOST_net_16906;
wire TIMEBOOST_net_7109;
wire TIMEBOOST_net_7108;
wire TIMEBOOST_net_16905;
wire TIMEBOOST_net_7107;
wire n_1417;
wire TIMEBOOST_net_16904;
wire TIMEBOOST_net_7106;
wire TIMEBOOST_net_15362;
wire TIMEBOOST_net_7104;
wire TIMEBOOST_net_15435;
wire TIMEBOOST_net_7103;
wire TIMEBOOST_net_22249;
wire TIMEBOOST_net_7102;
wire TIMEBOOST_net_7101;
wire n_1418;
wire TIMEBOOST_net_12742;
wire TIMEBOOST_net_15353;
wire TIMEBOOST_net_7098;
wire TIMEBOOST_net_14453;
wire n_1419;
wire TIMEBOOST_net_16717;
wire n_14197;
wire TIMEBOOST_net_21332;
wire TIMEBOOST_net_9763;
wire TIMEBOOST_net_16903;
wire TIMEBOOST_net_7092;
wire TIMEBOOST_net_16902;
wire n_1421;
wire TIMEBOOST_net_16901;
wire TIMEBOOST_net_12876;
wire TIMEBOOST_net_16055;
wire TIMEBOOST_net_14328;
wire n_1422;
wire TIMEBOOST_net_12788;
wire n_14226;
wire TIMEBOOST_net_16899;
wire TIMEBOOST_net_12910;
wire n_1423;
wire TIMEBOOST_net_16898;
wire TIMEBOOST_net_21902;
wire TIMEBOOST_net_16897;
wire n_1424;
wire TIMEBOOST_net_21862;
wire TIMEBOOST_net_12905;
wire TIMEBOOST_net_20266;
wire TIMEBOOST_net_22018;
wire TIMEBOOST_net_17125;
wire n_1425;
wire n_14250;
wire n_14251;
wire n_14252;
wire n_14253;
wire n_14254;
wire n_14255;
wire n_14256;
wire n_14257;
wire n_14258;
wire n_1426;
wire n_14260;
wire n_14261;
wire n_14264;
wire n_14268;
wire n_14269;
wire n_14270;
wire n_14271;
wire n_14272;
wire n_14273;
wire n_14274;
wire n_14275;
wire n_14277;
wire n_1428;
wire n_14283;
wire n_14284;
wire n_14285;
wire n_14286;
wire n_1429;
wire n_14290;
wire n_14291;
wire n_14292;
wire n_14293;
wire n_14295;
wire n_14296;
wire n_14298;
wire n_143;
wire n_14300;
wire n_14301;
wire n_14302;
wire n_14303;
wire n_14304;
wire n_14305;
wire n_14306;
wire n_14307;
wire n_14308;
wire n_14309;
wire n_1431;
wire n_14310;
wire n_14311;
wire n_14312;
wire n_14313;
wire n_14314;
wire n_14315;
wire n_14316;
wire n_14317;
wire n_14318;
wire n_14319;
wire n_1432;
wire n_14320;
wire n_14321;
wire n_14322;
wire n_14323;
wire n_14324;
wire n_14325;
wire n_14326;
wire n_14327;
wire n_14328;
wire n_14329;
wire n_1433;
wire n_14330;
wire n_14331;
wire n_14332;
wire n_14333;
wire n_14334;
wire n_14335;
wire n_14336;
wire n_14337;
wire n_14338;
wire n_14339;
wire n_1434;
wire n_14340;
wire n_14341;
wire n_14342;
wire n_14343;
wire n_14344;
wire n_14345;
wire n_14346;
wire n_14347;
wire n_14348;
wire n_14349;
wire n_1435;
wire n_14350;
wire n_14351;
wire n_14352;
wire n_14353;
wire n_14354;
wire n_14355;
wire n_14356;
wire n_14357;
wire n_14358;
wire n_14359;
wire n_1436;
wire n_14360;
wire n_14361;
wire n_14362;
wire n_14363;
wire n_14364;
wire n_14365;
wire n_14366;
wire n_14367;
wire n_14368;
wire n_14369;
wire n_1437;
wire n_14370;
wire n_14371;
wire n_14372;
wire n_14373;
wire n_14374;
wire n_14375;
wire n_14376;
wire n_14377;
wire n_14378;
wire n_14379;
wire n_1438;
wire n_14380;
wire n_14381;
wire n_14382;
wire n_14383;
wire n_14384;
wire n_14385;
wire n_14386;
wire n_14387;
wire n_14388;
wire n_14389;
wire n_1439;
wire n_14390;
wire n_14391;
wire n_14392;
wire n_14393;
wire n_14394;
wire n_14396;
wire n_14397;
wire TIMEBOOST_net_10300;
wire n_1440;
wire n_14401;
wire n_14402;
wire n_14403;
wire n_14407;
wire n_14408;
wire n_1441;
wire n_14410;
wire n_14413;
wire n_14414;
wire n_14415;
wire n_14416;
wire n_14419;
wire n_1442;
wire n_14420;
wire n_14421;
wire n_14422;
wire n_14426;
wire n_14427;
wire n_14428;
wire n_14429;
wire n_1443;
wire n_14430;
wire n_14431;
wire n_14432;
wire n_14433;
wire n_14434;
wire n_14435;
wire n_14436;
wire n_14437;
wire n_14438;
wire n_14439;
wire n_1444;
wire n_14440;
wire n_14441;
wire n_14442;
wire n_14443;
wire n_14444;
wire n_14445;
wire n_14446;
wire n_14447;
wire n_14448;
wire n_14449;
wire n_1445;
wire n_14451;
wire n_14454;
wire n_14456;
wire n_14457;
wire n_14458;
wire n_14459;
wire n_1446;
wire n_14460;
wire n_14461;
wire n_14462;
wire n_14467;
wire n_14468;
wire n_14469;
wire n_1447;
wire n_14471;
wire n_14472;
wire n_14473;
wire n_14474;
wire n_14475;
wire n_14476;
wire n_14477;
wire n_14478;
wire n_14479;
wire n_1448;
wire n_14480;
wire n_14481;
wire n_14482;
wire n_14483;
wire n_14484;
wire n_14485;
wire n_14486;
wire n_14487;
wire n_14489;
wire n_1449;
wire n_14490;
wire n_14491;
wire n_14493;
wire n_14494;
wire n_14495;
wire n_14497;
wire n_14498;
wire n_14499;
wire n_1450;
wire n_14500;
wire n_14504;
wire n_14505;
wire n_14507;
wire n_14508;
wire n_14510;
wire n_14511;
wire n_14512;
wire n_14513;
wire n_14514;
wire n_14515;
wire n_14517;
wire n_14518;
wire TIMEBOOST_net_16383;
wire n_1452;
wire n_14521;
wire n_14526;
wire TIMEBOOST_net_10055;
wire n_14528;
wire n_14529;
wire n_1453;
wire n_14530;
wire n_14531;
wire n_14532;
wire n_14534;
wire n_14535;
wire n_14536;
wire n_14539;
wire n_1454;
wire n_14541;
wire n_14543;
wire n_14544;
wire n_14545;
wire n_14547;
wire n_14548;
wire n_14549;
wire n_14550;
wire n_14551;
wire n_14554;
wire n_14556;
wire n_14557;
wire n_14558;
wire n_14559;
wire n_14560;
wire n_14563;
wire n_14564;
wire n_14565;
wire n_14566;
wire n_14567;
wire n_14569;
wire n_14570;
wire n_14571;
wire n_14572;
wire TIMEBOOST_net_14245;
wire n_14577;
wire n_14578;
wire n_14579;
wire n_14580;
wire n_14582;
wire n_14583;
wire n_14585;
wire n_14586;
wire n_14588;
wire n_14589;
wire n_1459;
wire n_14590;
wire n_14591;
wire n_14592;
wire n_14593;
wire n_14594;
wire n_14595;
wire n_14596;
wire n_14597;
wire n_14598;
wire n_14599;
wire n_1460;
wire n_14601;
wire n_14602;
wire n_14603;
wire n_14604;
wire n_14605;
wire n_14607;
wire n_14608;
wire n_14609;
wire n_1461;
wire n_14610;
wire n_14611;
wire n_14612;
wire n_14613;
wire n_14614;
wire n_14615;
wire n_14616;
wire n_14617;
wire n_14618;
wire n_14619;
wire n_14620;
wire n_14621;
wire n_14622;
wire n_14623;
wire n_14624;
wire n_14625;
wire n_14626;
wire n_14627;
wire n_14628;
wire n_14629;
wire n_1463;
wire n_14630;
wire n_14631;
wire n_14632;
wire n_14633;
wire n_14634;
wire n_14635;
wire n_14636;
wire n_14637;
wire n_14638;
wire n_14639;
wire n_14640;
wire n_14641;
wire n_14642;
wire n_14643;
wire n_14644;
wire n_14645;
wire n_14646;
wire n_14648;
wire n_14649;
wire n_1465;
wire n_14650;
wire n_14651;
wire n_14652;
wire n_14653;
wire n_14654;
wire n_14655;
wire n_14656;
wire n_14657;
wire n_14658;
wire n_14659;
wire n_14661;
wire n_14662;
wire n_14663;
wire n_14664;
wire n_14665;
wire n_14666;
wire n_14667;
wire n_14668;
wire n_14669;
wire n_1467;
wire n_14670;
wire n_14671;
wire TIMEBOOST_net_11485;
wire n_14674;
wire TIMEBOOST_net_11483;
wire n_14678;
wire TIMEBOOST_net_16840;
wire n_1468;
wire n_14681;
wire n_14682;
wire n_14683;
wire n_14685;
wire n_14686;
wire n_14687;
wire n_14688;
wire n_14689;
wire n_1469;
wire n_14690;
wire n_14691;
wire TIMEBOOST_net_21333;
wire n_14694;
wire n_14695;
wire n_14696;
wire n_14697;
wire n_14698;
wire n_14699;
wire n_1470;
wire n_14700;
wire n_14701;
wire n_14702;
wire n_14703;
wire n_14705;
wire n_14706;
wire n_14708;
wire n_14709;
wire n_1471;
wire n_14710;
wire n_14711;
wire n_14713;
wire n_14715;
wire n_14717;
wire n_14719;
wire n_1472;
wire n_14721;
wire n_14722;
wire n_14723;
wire n_14724;
wire n_14725;
wire n_14726;
wire n_14727;
wire n_14728;
wire n_14730;
wire n_14731;
wire n_14733;
wire n_14734;
wire n_14738;
wire n_1474;
wire n_14740;
wire n_14741;
wire TIMEBOOST_net_16860;
wire TIMEBOOST_net_16859;
wire n_14746;
wire n_14747;
wire TIMEBOOST_net_16858;
wire n_1475;
wire n_14750;
wire n_14751;
wire n_14753;
wire TIMEBOOST_net_11632;
wire n_14755;
wire n_14756;
wire n_14757;
wire n_14759;
wire n_1476;
wire n_14760;
wire n_14761;
wire n_14762;
wire n_14763;
wire n_14764;
wire n_14765;
wire n_14766;
wire n_14767;
wire n_14768;
wire n_14769;
wire n_1477;
wire n_14770;
wire n_14772;
wire n_14773;
wire n_14775;
wire n_14776;
wire n_14777;
wire n_14778;
wire n_1478;
wire n_14780;
wire n_14781;
wire n_14783;
wire n_14784;
wire n_14786;
wire n_14789;
wire n_1479;
wire n_14790;
wire n_14791;
wire n_14792;
wire n_14793;
wire n_14794;
wire n_14796;
wire n_14797;
wire n_14798;
wire n_14799;
wire n_148;
wire n_1480;
wire n_14800;
wire n_14802;
wire n_14803;
wire n_14804;
wire n_14805;
wire n_14806;
wire n_14807;
wire n_14808;
wire n_1481;
wire n_14810;
wire n_14811;
wire n_14812;
wire n_14813;
wire n_14814;
wire n_14815;
wire n_14816;
wire n_14817;
wire n_14818;
wire n_14819;
wire n_1482;
wire n_14821;
wire n_14822;
wire n_14824;
wire n_14825;
wire n_14826;
wire n_14828;
wire n_14829;
wire n_1483;
wire n_14830;
wire n_14832;
wire n_14833;
wire n_14834;
wire n_14836;
wire n_14837;
wire n_14838;
wire n_14839;
wire n_1484;
wire n_14840;
wire n_14841;
wire n_14842;
wire n_14844;
wire n_14845;
wire n_14846;
wire n_14847;
wire n_14848;
wire n_14849;
wire n_1485;
wire n_14850;
wire n_14851;
wire n_14852;
wire n_14853;
wire n_14854;
wire n_14855;
wire n_14856;
wire n_14858;
wire n_14859;
wire n_1486;
wire n_14860;
wire n_14861;
wire n_14862;
wire n_14863;
wire n_14864;
wire n_14865;
wire n_14866;
wire n_14867;
wire n_14869;
wire n_14871;
wire n_14873;
wire n_14875;
wire n_14877;
wire n_14879;
wire n_1488;
wire n_14880;
wire n_14881;
wire n_14883;
wire n_14884;
wire n_14885;
wire n_14887;
wire n_14888;
wire n_14889;
wire n_14890;
wire n_14891;
wire n_14892;
wire n_14893;
wire n_14894;
wire n_14895;
wire n_14896;
wire n_14897;
wire n_14898;
wire n_14899;
wire n_14900;
wire n_14901;
wire n_14902;
wire n_14903;
wire n_14904;
wire n_14905;
wire n_14906;
wire n_14907;
wire n_14908;
wire n_14909;
wire n_14910;
wire n_14911;
wire n_14912;
wire n_14913;
wire n_14914;
wire n_14915;
wire n_14916;
wire n_14917;
wire n_14918;
wire n_14919;
wire n_14920;
wire n_14921;
wire n_14922;
wire n_14923;
wire n_14924;
wire n_14925;
wire n_14926;
wire n_14927;
wire n_14928;
wire n_14929;
wire n_1493;
wire n_14930;
wire n_14931;
wire n_14932;
wire n_14933;
wire n_14934;
wire n_14939;
wire n_1495;
wire n_14956;
wire n_14957;
wire n_14960;
wire n_14961;
wire n_14963;
wire n_14965;
wire n_14967;
wire n_1497;
wire n_14971;
wire n_14981;
wire n_1499;
wire n_15;
wire n_150;
wire n_15001;
wire n_1501;
wire n_15014;
wire n_1502;
wire n_1503;
wire TIMEBOOST_net_13446;
wire n_1504;
wire n_1505;
wire n_15054;
wire n_15055;
wire n_15065;
wire n_1507;
wire n_1508;
wire n_1509;
wire n_1510;
wire n_15117;
wire n_1512;
wire n_15125;
wire n_15128;
wire n_1513;
wire n_1514;
wire n_15142;
wire n_1515;
wire n_15187;
wire n_15188;
wire n_1519;
wire n_15196;
wire n_15197;
wire n_152;
wire n_15204;
wire n_15210;
wire n_15217;
wire n_1522;
wire n_1523;
wire n_15231;
wire n_1524;
wire n_15249;
wire n_15260;
wire n_15261;
wire n_15262;
wire n_15275;
wire n_15276;
wire n_15291;
wire n_15292;
wire n_15295;
wire n_15301;
wire n_15302;
wire n_15313;
wire n_15314;
wire n_15317;
wire n_1532;
wire n_15324;
wire n_15325;
wire n_1533;
wire n_15330;
wire n_15331;
wire n_15347;
wire n_1535;
wire n_1536;
wire n_15365;
wire n_1537;
wire n_15370;
wire n_15371;
wire n_15372;
wire n_15373;
wire n_15376;
wire n_15377;
wire TIMEBOOST_net_16753;
wire n_15385;
wire n_15388;
wire n_15389;
wire n_1539;
wire n_15390;
wire n_15397;
wire n_1540;
wire n_15401;
wire n_15402;
wire n_15403;
wire n_15405;
wire n_15406;
wire n_15407;
wire n_1541;
wire n_15414;
wire n_15417;
wire n_1542;
wire TIMEBOOST_net_22701;
wire n_15434;
wire n_15435;
wire n_15436;
wire n_15438;
wire n_15439;
wire n_15440;
wire n_15441;
wire n_15442;
wire n_15444;
wire n_15445;
wire n_15446;
wire n_1545;
wire n_15453;
wire n_15456;
wire n_15458;
wire n_1546;
wire n_15467;
wire n_1547;
wire n_15474;
wire n_1548;
wire n_1549;
wire n_1551;
wire n_15512;
wire TIMEBOOST_net_11348;
wire n_15514;
wire n_15515;
wire n_15516;
wire n_15517;
wire n_15518;
wire n_15527;
wire n_15528;
wire n_15529;
wire n_1553;
wire n_15534;
wire n_15538;
wire n_15539;
wire n_1554;
wire n_15540;
wire n_15549;
wire n_1555;
wire n_15551;
wire n_15552;
wire n_15553;
wire n_15558;
wire n_15560;
wire n_15562;
wire n_15565;
wire n_15566;
wire n_15567;
wire n_15568;
wire n_15569;
wire n_1557;
wire n_15581;
wire n_15584;
wire n_15585;
wire n_15586;
wire n_15587;
wire n_15589;
wire n_1559;
wire n_15590;
wire n_15591;
wire n_15592;
wire n_15593;
wire n_15594;
wire n_15598;
wire n_156;
wire n_15607;
wire n_1561;
wire n_15611;
wire n_15614;
wire n_1562;
wire n_1563;
wire n_15638;
wire n_1564;
wire n_15645;
wire n_1565;
wire n_1566;
wire n_1567;
wire n_1568;
wire n_15680;
wire n_15689;
wire n_1569;
wire n_15694;
wire n_15695;
wire g64948_db;
wire n_15698;
wire n_15699;
wire n_1571;
wire TIMEBOOST_net_13879;
wire n_15729;
wire n_1573;
wire TIMEBOOST_net_14632;
wire n_15732;
wire n_15733;
wire n_15735;
wire n_15736;
wire n_15738;
wire n_15739;
wire n_1574;
wire n_15741;
wire n_15744;
wire n_15746;
wire n_15748;
wire TIMEBOOST_net_20577;
wire n_15754;
wire n_15755;
wire n_15756;
wire n_15757;
wire n_15758;
wire n_15759;
wire TIMEBOOST_net_23253;
wire n_15760;
wire n_15762;
wire n_15769;
wire TIMEBOOST_net_12496;
wire n_15788;
wire n_15798;
wire n_15802;
wire n_15805;
wire n_15808;
wire n_1581;
wire n_15813;
wire n_1582;
wire n_15823;
wire n_15824;
wire n_1583;
wire TIMEBOOST_net_20179;
wire n_1585;
wire n_15854;
wire n_15856;
wire n_15859;
wire n_1586;
wire n_1588;
wire n_1589;
wire n_1590;
wire n_15908;
wire TIMEBOOST_net_342;
wire TIMEBOOST_net_20975;
wire n_15910;
wire n_15914;
wire n_15915;
wire n_15917;
wire n_15918;
wire n_15919;
wire TIMEBOOST_net_20404;
wire n_15920;
wire TIMEBOOST_net_13366;
wire n_15922;
wire n_15923;
wire n_15924;
wire n_15927;
wire n_15929;
wire n_1593;
wire n_15931;
wire n_15932;
wire n_15935;
wire TIMEBOOST_net_16809;
wire n_15937;
wire n_15939;
wire n_1594;
wire n_15940;
wire n_15941;
wire n_15942;
wire n_1595;
wire n_15958;
wire n_15959;
wire n_15960;
wire n_15969;
wire n_15979;
wire n_1598;
wire n_15980;
wire n_15981;
wire n_15982;
wire n_15985;
wire n_15988;
wire n_1599;
wire n_15994;
wire n_15996;
wire n_15998;
wire n_15999;
wire n_160;
wire n_1600;
wire n_16000;
wire n_16001;
wire n_16002;
wire n_16003;
wire n_16015;
wire n_16016;
wire n_1602;
wire n_16021;
wire n_16022;
wire n_16027;
wire n_1603;
wire n_16030;
wire n_16033;
wire n_16034;
wire n_16036;
wire n_16046;
wire n_16047;
wire n_16048;
wire n_16049;
wire n_1605;
wire n_16052;
wire TIMEBOOST_net_20658;
wire n_16066;
wire TIMEBOOST_net_15706;
wire n_1607;
wire n_16070;
wire n_16071;
wire n_16075;
wire n_16076;
wire n_1608;
wire n_16089;
wire n_1609;
wire n_1610;
wire n_16101;
wire n_16102;
wire n_16103;
wire n_16105;
wire TIMEBOOST_net_20405;
wire n_1612;
wire n_1613;
wire n_16131;
wire n_1614;
wire n_1615;
wire n_16150;
wire n_16151;
wire n_16152;
wire n_16153;
wire n_16154;
wire n_16156;
wire n_16157;
wire TIMEBOOST_net_11296;
wire n_16159;
wire n_1616;
wire n_16160;
wire n_16161;
wire n_16162;
wire n_16163;
wire n_16164;
wire n_16165;
wire TIMEBOOST_net_12449;
wire n_16167;
wire n_16168;
wire n_16169;
wire n_16170;
wire n_16173;
wire n_16175;
wire TIMEBOOST_net_10438;
wire n_16183;
wire n_1619;
wire n_16205;
wire n_16206;
wire n_16207;
wire n_16208;
wire n_16209;
wire n_1621;
wire n_16210;
wire n_16211;
wire n_16212;
wire n_16213;
wire n_16220;
wire n_16221;
wire n_16222;
wire n_16223;
wire n_16224;
wire n_16225;
wire n_16226;
wire n_16227;
wire n_16228;
wire n_16229;
wire n_1623;
wire n_16230;
wire n_16231;
wire n_16233;
wire n_16234;
wire n_16235;
wire n_16236;
wire n_16237;
wire n_16238;
wire n_16239;
wire n_1624;
wire n_16240;
wire n_16241;
wire n_16242;
wire n_16243;
wire n_16244;
wire n_16247;
wire n_16248;
wire n_16249;
wire n_1625;
wire n_16250;
wire n_16251;
wire n_16252;
wire n_16253;
wire n_16254;
wire n_16255;
wire n_16256;
wire n_16257;
wire n_16258;
wire n_16259;
wire n_1626;
wire n_16260;
wire n_16261;
wire n_16262;
wire n_16264;
wire n_16265;
wire n_16268;
wire n_16271;
wire n_16273;
wire n_16275;
wire n_1628;
wire n_16280;
wire n_16284;
wire n_16285;
wire n_16286;
wire n_16287;
wire n_16288;
wire n_16289;
wire n_1629;
wire n_16290;
wire n_16291;
wire n_16293;
wire n_16299;
wire n_1630;
wire n_16300;
wire n_16301;
wire n_16304;
wire n_16305;
wire n_16306;
wire n_16307;
wire n_16309;
wire n_1631;
wire n_16310;
wire n_16311;
wire n_16313;
wire n_16317;
wire n_1632;
wire n_16322;
wire n_16325;
wire n_16326;
wire n_1633;
wire n_16330;
wire n_16331;
wire n_16332;
wire n_16334;
wire TIMEBOOST_net_13041;
wire n_1634;
wire n_1635;
wire n_16350;
wire n_16351;
wire n_16352;
wire n_16354;
wire n_16358;
wire n_16364;
wire n_16368;
wire n_16388;
wire n_16389;
wire n_1639;
wire n_16390;
wire n_16391;
wire n_16392;
wire n_16393;
wire n_16394;
wire n_16395;
wire n_16396;
wire n_16397;
wire n_16398;
wire n_16399;
wire n_1640;
wire n_16400;
wire n_16401;
wire n_16402;
wire n_16403;
wire n_16404;
wire n_16406;
wire n_16408;
wire n_16409;
wire n_1641;
wire n_16410;
wire n_16411;
wire n_16412;
wire n_16413;
wire n_1642;
wire n_16424;
wire n_16425;
wire n_16427;
wire n_16428;
wire n_16429;
wire n_1643;
wire TIMEBOOST_net_16519;
wire n_16433;
wire n_16434;
wire n_16435;
wire n_16436;
wire n_16437;
wire n_16438;
wire n_16439;
wire n_16441;
wire n_16442;
wire n_16444;
wire n_16445;
wire n_1645;
wire n_16451;
wire n_16452;
wire n_16455;
wire n_16456;
wire TIMEBOOST_net_21855;
wire TIMEBOOST_net_13396;
wire n_16459;
wire TIMEBOOST_net_23395;
wire n_16460;
wire n_16462;
wire n_1647;
wire n_16474;
wire n_16475;
wire n_1648;
wire n_16485;
wire n_16486;
wire n_16487;
wire n_1649;
wire n_16490;
wire n_16491;
wire n_16492;
wire n_16493;
wire n_16494;
wire n_16495;
wire n_16496;
wire n_16497;
wire n_16499;
wire n_16501;
wire n_16503;
wire n_16504;
wire n_16507;
wire n_16511;
wire n_16512;
wire n_16513;
wire n_16516;
wire n_1652;
wire n_16520;
wire n_16521;
wire n_16523;
wire n_16524;
wire n_16533;
wire n_16534;
wire n_16535;
wire n_16536;
wire n_16537;
wire n_16538;
wire n_16539;
wire n_1654;
wire n_16540;
wire n_16541;
wire n_16542;
wire n_16543;
wire n_16544;
wire n_16547;
wire n_1655;
wire n_16550;
wire n_16552;
wire n_16553;
wire n_16554;
wire n_1656;
wire n_16560;
wire n_16564;
wire n_16566;
wire n_1657;
wire n_16572;
wire n_16573;
wire n_16576;
wire n_16577;
wire n_16578;
wire n_16579;
wire n_1658;
wire n_16581;
wire n_16582;
wire n_16583;
wire n_16584;
wire n_16585;
wire n_16586;
wire n_16587;
wire n_16588;
wire n_16589;
wire n_1659;
wire n_16591;
wire n_16592;
wire n_16594;
wire n_16595;
wire n_16596;
wire n_16597;
wire n_16599;
wire n_1660;
wire n_16600;
wire n_16601;
wire n_16602;
wire n_16603;
wire n_16605;
wire TIMEBOOST_net_12906;
wire TIMEBOOST_net_14265;
wire TIMEBOOST_net_12907;
wire n_16610;
wire n_16611;
wire n_16614;
wire n_16615;
wire n_16616;
wire n_16617;
wire n_1662;
wire n_16622;
wire n_16623;
wire n_16624;
wire n_16625;
wire TIMEBOOST_net_22322;
wire TIMEBOOST_net_23335;
wire TIMEBOOST_net_21520;
wire n_16635;
wire n_16637;
wire n_16657;
wire n_1666;
wire n_1667;
wire n_1668;
wire n_16685;
wire n_1669;
wire n_16690;
wire n_16695;
wire n_16696;
wire n_16698;
wire n_1673;
wire n_16738;
wire n_1674;
wire n_16748;
wire n_1675;
wire n_16763;
wire n_1677;
wire n_16779;
wire n_1678;
wire n_1679;
wire n_16791;
wire n_16798;
wire n_168;
wire n_1680;
wire n_1681;
wire n_16810;
wire n_16816;
wire n_16818;
wire n_1683;
wire n_16834;
wire n_16835;
wire n_16836;
wire n_16837;
wire n_16838;
wire n_16839;
wire n_1684;
wire n_16840;
wire n_16841;
wire n_16842;
wire n_16843;
wire n_16844;
wire n_16845;
wire n_16848;
wire n_16849;
wire n_1685;
wire n_16850;
wire n_16851;
wire n_16852;
wire n_16853;
wire n_16854;
wire n_16855;
wire n_1686;
wire n_16860;
wire n_16864;
wire n_16867;
wire n_16871;
wire n_16876;
wire n_1688;
wire n_16888;
wire n_1689;
wire n_16891;
wire n_169;
wire n_1690;
wire n_16904;
wire n_16906;
wire n_16910;
wire n_16911;
wire n_16914;
wire n_16916;
wire n_1692;
wire n_1693;
wire n_16936;
wire n_1694;
wire n_16940;
wire n_16942;
wire n_16945;
wire n_16949;
wire n_1695;
wire n_16952;
wire n_1696;
wire n_16963;
wire n_16964;
wire n_16966;
wire n_16967;
wire n_1697;
wire n_16970;
wire n_16974;
wire n_16976;
wire n_16977;
wire n_1698;
wire n_16980;
wire n_16981;
wire n_16984;
wire n_16985;
wire n_16986;
wire n_16987;
wire n_1699;
wire n_16992;
wire n_17;
wire n_1701;
wire n_17016;
wire n_17017;
wire g52465_da;
wire TIMEBOOST_net_16872;
wire TIMEBOOST_net_23467;
wire TIMEBOOST_net_22416;
wire n_17021;
wire n_17027;
wire n_17028;
wire n_17029;
wire n_17030;
wire n_17031;
wire n_17032;
wire n_17034;
wire n_17035;
wire n_17036;
wire n_17039;
wire n_1704;
wire n_17040;
wire n_17041;
wire n_17042;
wire n_17043;
wire n_17044;
wire n_17045;
wire n_17046;
wire n_17048;
wire n_17049;
wire n_17050;
wire n_17051;
wire n_1707;
wire n_1709;
wire n_1714;
wire n_1715;
wire n_1716;
wire TIMEBOOST_net_20929;
wire n_1719;
wire n_1721;
wire n_1724;
wire n_1737;
wire n_1739;
wire n_1740;
wire n_1742;
wire n_1743;
wire n_1746;
wire n_1748;
wire n_1750;
wire n_1752;
wire n_1754;
wire n_1755;
wire n_1758;
wire n_1759;
wire n_177;
wire n_1774;
wire n_1777;
wire n_1779;
wire n_1780;
wire n_1781;
wire n_1782;
wire n_1784;
wire n_1785;
wire n_1786;
wire n_1787;
wire n_1788;
wire n_1789;
wire n_1790;
wire n_1793;
wire n_1794;
wire n_1795;
wire n_1798;
wire n_1799;
wire n_18;
wire n_1800;
wire n_1802;
wire n_1803;
wire n_1804;
wire n_1805;
wire n_1806;
wire n_1808;
wire n_1809;
wire n_181;
wire n_1810;
wire n_1812;
wire n_1813;
wire n_1814;
wire n_1815;
wire n_1816;
wire n_1817;
wire n_1819;
wire n_1820;
wire n_1821;
wire n_1822;
wire n_1823;
wire n_1824;
wire n_1825;
wire n_1826;
wire n_1827;
wire n_1828;
wire n_1829;
wire n_1832;
wire n_1834;
wire n_1838;
wire TIMEBOOST_net_13107;
wire n_1845;
wire TIMEBOOST_net_16365;
wire n_1847;
wire n_1848;
wire TIMEBOOST_net_20583;
wire TIMEBOOST_net_17505;
wire n_1852;
wire n_1854;
wire n_1855;
wire n_1858;
wire n_1859;
wire n_1860;
wire n_1862;
wire n_1864;
wire n_1865;
wire n_1867;
wire n_1870;
wire n_1871;
wire n_1872;
wire n_1873;
wire n_1876;
wire n_1879;
wire n_188;
wire n_1880;
wire n_1881;
wire TIMEBOOST_net_13397;
wire n_1886;
wire n_1889;
wire n_1893;
wire n_1895;
wire n_1896;
wire TIMEBOOST_net_23556;
wire n_1901;
wire n_1903;
wire n_1904;
wire n_1905;
wire n_1906;
wire n_1907;
wire n_1909;
wire n_191;
wire n_1912;
wire TIMEBOOST_net_20508;
wire n_1915;
wire n_1916;
wire n_1919;
wire n_1920;
wire n_1921;
wire n_1924;
wire n_193;
wire TIMEBOOST_net_13088;
wire TIMEBOOST_net_23123;
wire n_1934;
wire n_1935;
wire n_1936;
wire n_1937;
wire n_1938;
wire TIMEBOOST_net_10825;
wire n_1942;
wire n_1943;
wire n_1944;
wire TIMEBOOST_net_22861;
wire n_1946;
wire n_1948;
wire n_1949;
wire n_1950;
wire n_1952;
wire n_1953;
wire n_1955;
wire n_1956;
wire n_1959;
wire n_1960;
wire n_1961;
wire n_1963;
wire n_1964;
wire n_1965;
wire n_1966;
wire n_1967;
wire n_1968;
wire n_1969;
wire n_1970;
wire n_1971;
wire n_1972;
wire n_1973;
wire n_1974;
wire n_1975;
wire n_1976;
wire TIMEBOOST_net_22951;
wire n_1979;
wire n_1981;
wire n_1985;
wire n_1986;
wire n_1987;
wire n_1989;
wire n_1990;
wire n_1992;
wire n_1993;
wire n_1994;
wire n_1995;
wire TIMEBOOST_net_23124;
wire n_1998;
wire n_1999;
wire n_2;
wire n_200;
wire n_2000;
wire n_2001;
wire n_2002;
wire TIMEBOOST_net_15375;
wire n_2007;
wire n_2008;
wire n_2009;
wire n_2010;
wire n_2011;
wire n_2012;
wire n_2013;
wire n_2014;
wire TIMEBOOST_net_15873;
wire n_2016;
wire n_2017;
wire n_2018;
wire n_2019;
wire n_202;
wire n_2022;
wire n_2023;
wire n_2024;
wire n_2027;
wire n_2028;
wire n_2029;
wire n_2031;
wire n_2034;
wire n_2035;
wire n_2036;
wire n_2037;
wire TIMEBOOST_net_8767;
wire n_204;
wire n_2040;
wire n_2041;
wire n_2042;
wire n_2043;
wire n_2044;
wire n_2046;
wire n_2047;
wire n_2049;
wire n_205;
wire n_2051;
wire n_2052;
wire n_2053;
wire n_2054;
wire n_2055;
wire n_2056;
wire n_2057;
wire n_2059;
wire n_206;
wire TIMEBOOST_net_22776;
wire n_2061;
wire n_2065;
wire n_2066;
wire n_2067;
wire n_2068;
wire n_2069;
wire n_207;
wire n_2070;
wire n_2071;
wire n_2072;
wire n_2074;
wire n_2075;
wire n_2076;
wire n_2077;
wire n_2078;
wire n_2079;
wire n_208;
wire n_2080;
wire n_2082;
wire n_2083;
wire n_2084;
wire n_2086;
wire n_2087;
wire n_2088;
wire n_2092;
wire n_2094;
wire n_21;
wire n_2100;
wire n_2101;
wire n_2102;
wire n_2103;
wire n_2104;
wire n_2105;
wire n_2106;
wire n_2108;
wire n_211;
wire n_2110;
wire n_2111;
wire n_2113;
wire n_2114;
wire n_2115;
wire n_2116;
wire n_2117;
wire n_2119;
wire n_2120;
wire n_2121;
wire n_2122;
wire n_2125;
wire n_2126;
wire n_2127;
wire n_2129;
wire n_213;
wire n_2131;
wire n_2132;
wire n_2134;
wire n_2135;
wire n_2136;
wire n_2137;
wire n_2138;
wire n_2140;
wire n_2146;
wire n_2147;
wire TIMEBOOST_net_21613;
wire n_2151;
wire n_2152;
wire n_2153;
wire n_2154;
wire n_2155;
wire TIMEBOOST_net_23480;
wire n_2158;
wire n_2159;
wire n_2161;
wire n_2162;
wire n_2163;
wire n_2165;
wire TIMEBOOST_net_20162;
wire n_2170;
wire n_2171;
wire n_2172;
wire TIMEBOOST_net_23479;
wire n_2174;
wire n_2175;
wire n_2176;
wire n_2177;
wire n_2178;
wire n_2179;
wire n_2180;
wire TIMEBOOST_net_16877;
wire n_2184;
wire TIMEBOOST_net_22512;
wire n_2186;
wire n_2187;
wire n_2189;
wire n_2191;
wire n_2192;
wire n_2193;
wire n_2194;
wire n_2195;
wire n_2197;
wire n_2198;
wire n_2199;
wire n_22;
wire n_2200;
wire n_2201;
wire n_2202;
wire n_2203;
wire n_2205;
wire n_2206;
wire n_2207;
wire n_2209;
wire n_221;
wire n_2210;
wire n_2211;
wire n_2212;
wire n_2213;
wire n_2214;
wire n_2215;
wire n_2218;
wire n_2219;
wire n_2223;
wire n_2224;
wire n_2225;
wire n_2226;
wire n_2227;
wire n_2228;
wire n_2229;
wire n_2230;
wire n_2231;
wire n_2232;
wire n_2233;
wire n_2234;
wire n_2235;
wire n_2236;
wire n_2237;
wire n_2238;
wire n_2243;
wire n_2244;
wire n_2245;
wire n_2246;
wire n_2247;
wire n_2248;
wire n_2249;
wire n_2250;
wire n_2251;
wire n_2252;
wire n_2253;
wire n_2254;
wire n_2255;
wire n_2256;
wire n_2257;
wire n_2258;
wire n_2259;
wire n_2260;
wire n_2261;
wire n_2262;
wire n_2263;
wire n_2264;
wire n_2266;
wire TIMEBOOST_net_14663;
wire n_2269;
wire n_227;
wire n_2271;
wire n_2272;
wire n_2273;
wire n_2274;
wire n_2275;
wire n_2276;
wire n_2280;
wire n_2281;
wire n_2284;
wire n_2285;
wire n_2286;
wire n_2287;
wire n_2289;
wire n_2291;
wire n_2292;
wire n_2293;
wire n_2295;
wire n_2297;
wire TIMEBOOST_net_7531;
wire n_2299;
wire n_23;
wire n_230;
wire n_2300;
wire n_2301;
wire n_2302;
wire n_2303;
wire n_2304;
wire n_2305;
wire n_2306;
wire n_2308;
wire n_231;
wire n_2311;
wire n_2313;
wire n_2314;
wire n_2315;
wire n_2316;
wire n_2319;
wire n_232;
wire n_2326;
wire n_2327;
wire n_2328;
wire n_2329;
wire n_233;
wire n_2331;
wire n_2337;
wire n_2339;
wire n_234;
wire n_2341;
wire n_2343;
wire n_2344;
wire n_2345;
wire n_2347;
wire n_2349;
wire n_235;
wire n_2350;
wire n_2351;
wire n_2352;
wire n_2353;
wire n_2354;
wire n_2356;
wire n_2358;
wire n_2359;
wire n_236;
wire n_2361;
wire n_2362;
wire n_2363;
wire n_2364;
wire n_2366;
wire n_2367;
wire n_2369;
wire n_2370;
wire n_2371;
wire n_2372;
wire n_2373;
wire n_2374;
wire n_2376;
wire n_2377;
wire TIMEBOOST_net_20665;
wire n_2380;
wire n_2386;
wire n_2387;
wire TIMEBOOST_net_21297;
wire n_2390;
wire n_2392;
wire n_2395;
wire n_2396;
wire n_2397;
wire n_2398;
wire n_2399;
wire n_24;
wire n_2400;
wire n_2401;
wire n_2402;
wire n_2405;
wire n_2406;
wire n_2407;
wire n_2409;
wire n_2410;
wire n_2411;
wire n_2412;
wire n_2414;
wire n_2415;
wire n_2416;
wire n_2418;
wire n_2419;
wire n_242;
wire n_2420;
wire n_2421;
wire n_2422;
wire n_2423;
wire n_2424;
wire n_2425;
wire n_2426;
wire n_2427;
wire n_2428;
wire n_2429;
wire n_243;
wire n_2430;
wire n_2431;
wire n_2432;
wire n_2433;
wire n_2434;
wire n_2435;
wire n_2436;
wire n_2437;
wire n_2438;
wire TIMEBOOST_net_158;
wire n_2440;
wire n_2441;
wire n_2442;
wire n_2443;
wire n_2445;
wire n_2446;
wire n_2447;
wire n_2449;
wire n_245;
wire n_2451;
wire n_2453;
wire n_2456;
wire n_2457;
wire n_2458;
wire n_2459;
wire n_2460;
wire n_2461;
wire n_2462;
wire n_2463;
wire n_2464;
wire n_2468;
wire n_2469;
wire n_247;
wire n_2471;
wire n_2473;
wire n_2474;
wire n_2475;
wire n_2476;
wire n_2477;
wire n_2478;
wire n_2479;
wire n_2482;
wire n_2483;
wire n_2485;
wire n_2486;
wire n_2487;
wire n_2488;
wire n_249;
wire n_2490;
wire n_2491;
wire n_2492;
wire n_2493;
wire n_2494;
wire n_2496;
wire n_2497;
wire n_2498;
wire n_2499;
wire n_2500;
wire n_2501;
wire n_2502;
wire n_2503;
wire n_2504;
wire n_2505;
wire n_2507;
wire n_2508;
wire n_2509;
wire n_251;
wire n_2510;
wire n_2512;
wire n_2513;
wire n_2514;
wire n_2515;
wire n_2516;
wire n_2517;
wire n_2518;
wire n_2519;
wire n_2520;
wire n_2521;
wire n_2522;
wire n_2524;
wire n_2526;
wire n_2527;
wire n_2528;
wire n_2530;
wire n_2531;
wire n_2533;
wire n_2534;
wire n_2536;
wire n_2537;
wire n_2539;
wire n_2540;
wire n_2541;
wire n_2542;
wire n_2543;
wire n_2544;
wire n_2545;
wire n_2546;
wire n_2547;
wire n_255;
wire n_2552;
wire n_2553;
wire n_2555;
wire n_2556;
wire n_2557;
wire n_2558;
wire n_2559;
wire n_2560;
wire n_2562;
wire n_2564;
wire n_2566;
wire n_2567;
wire n_2568;
wire n_2569;
wire n_257;
wire n_2570;
wire n_2571;
wire n_2572;
wire n_2573;
wire n_2574;
wire n_2575;
wire n_2576;
wire n_2577;
wire n_2579;
wire n_2580;
wire n_2581;
wire n_2582;
wire n_2583;
wire n_2584;
wire n_2585;
wire n_2586;
wire n_2587;
wire n_2588;
wire n_2590;
wire n_2592;
wire n_2593;
wire n_2594;
wire n_2595;
wire n_2596;
wire n_2597;
wire n_2598;
wire n_2599;
wire n_26;
wire n_2600;
wire n_2601;
wire n_2602;
wire n_2603;
wire n_2604;
wire n_2605;
wire n_2606;
wire n_2608;
wire n_2609;
wire n_261;
wire n_2610;
wire n_2611;
wire n_2612;
wire n_2613;
wire n_2614;
wire TIMEBOOST_net_12483;
wire n_2616;
wire n_2619;
wire n_2620;
wire n_2621;
wire n_2622;
wire n_2623;
wire n_2624;
wire n_2625;
wire TIMEBOOST_net_23314;
wire n_2629;
wire n_263;
wire n_2630;
wire n_2631;
wire n_2632;
wire n_2633;
wire n_2634;
wire n_2635;
wire n_2636;
wire n_2637;
wire n_2638;
wire n_2639;
wire n_2640;
wire n_2641;
wire n_2643;
wire n_2644;
wire n_2645;
wire n_2646;
wire n_2648;
wire n_2649;
wire n_2651;
wire n_2652;
wire n_2653;
wire n_2654;
wire n_2655;
wire n_2656;
wire n_2657;
wire n_2658;
wire n_2659;
wire n_2660;
wire n_2661;
wire n_2662;
wire n_2663;
wire n_2664;
wire n_2665;
wire n_2666;
wire n_2667;
wire n_2668;
wire n_2669;
wire n_2670;
wire n_2671;
wire n_2672;
wire n_2673;
wire n_2674;
wire n_2675;
wire n_2676;
wire n_2677;
wire n_2678;
wire n_2679;
wire n_268;
wire n_2680;
wire n_2681;
wire n_2682;
wire n_2683;
wire n_2684;
wire n_2685;
wire n_2687;
wire n_2691;
wire n_2692;
wire n_2693;
wire n_2694;
wire n_2695;
wire n_2696;
wire n_2697;
wire n_2698;
wire n_2699;
wire n_27;
wire n_2700;
wire n_2701;
wire n_2702;
wire n_2705;
wire n_2706;
wire n_2707;
wire n_2708;
wire n_2709;
wire n_271;
wire n_2710;
wire n_2711;
wire n_2712;
wire n_2713;
wire n_2714;
wire n_2715;
wire n_2716;
wire n_2717;
wire n_2718;
wire n_2719;
wire n_272;
wire n_2720;
wire n_2721;
wire n_2722;
wire n_2723;
wire n_2725;
wire n_2726;
wire n_2727;
wire n_2728;
wire n_2729;
wire n_2730;
wire n_2731;
wire n_2732;
wire n_2734;
wire n_2735;
wire n_2738;
wire n_2739;
wire n_2740;
wire n_2742;
wire n_2744;
wire n_2745;
wire n_2746;
wire n_2747;
wire n_2748;
wire n_2750;
wire n_2751;
wire n_2752;
wire n_2753;
wire n_2754;
wire n_2755;
wire n_2756;
wire n_2757;
wire n_276;
wire n_2761;
wire n_2762;
wire n_2763;
wire n_2764;
wire n_2765;
wire n_2767;
wire n_2768;
wire n_2769;
wire n_277;
wire n_2770;
wire n_2774;
wire n_2775;
wire n_2776;
wire n_2777;
wire n_2778;
wire n_2779;
wire n_278;
wire n_2780;
wire n_2781;
wire n_2782;
wire n_2783;
wire n_2784;
wire n_2785;
wire n_2786;
wire n_2787;
wire n_2788;
wire n_2789;
wire n_279;
wire n_2790;
wire n_2792;
wire n_2793;
wire n_2794;
wire n_2795;
wire n_2797;
wire n_2799;
wire n_28;
wire n_2801;
wire TIMEBOOST_net_14795;
wire n_2803;
wire n_2804;
wire TIMEBOOST_net_15881;
wire n_2806;
wire n_2807;
wire n_2809;
wire n_2812;
wire n_2813;
wire n_2814;
wire n_2815;
wire n_2818;
wire n_2819;
wire n_282;
wire n_2820;
wire n_2821;
wire n_2822;
wire n_2823;
wire n_2824;
wire n_2825;
wire n_2826;
wire n_2828;
wire n_2829;
wire n_2830;
wire n_2831;
wire n_2833;
wire n_2834;
wire n_2835;
wire n_2836;
wire n_2838;
wire n_2839;
wire n_2840;
wire n_2841;
wire n_2842;
wire n_2843;
wire n_2844;
wire n_2846;
wire n_2847;
wire n_2848;
wire n_2849;
wire n_285;
wire n_2851;
wire n_2852;
wire n_2853;
wire n_2854;
wire n_2855;
wire n_2856;
wire n_2857;
wire n_2858;
wire n_2859;
wire n_2860;
wire n_2864;
wire n_2865;
wire n_2866;
wire n_2867;
wire n_2868;
wire n_2869;
wire n_287;
wire n_2870;
wire n_2871;
wire n_2872;
wire n_2873;
wire n_2874;
wire n_2876;
wire n_2877;
wire n_2878;
wire n_288;
wire n_2883;
wire n_2887;
wire n_2888;
wire n_2897;
wire n_2898;
wire n_290;
wire n_2900;
wire n_2902;
wire n_2904;
wire n_2905;
wire n_2906;
wire n_2907;
wire n_2909;
wire n_2910;
wire n_2913;
wire n_2914;
wire n_2915;
wire n_2916;
wire n_2917;
wire n_2918;
wire n_2919;
wire n_292;
wire n_2920;
wire n_2921;
wire n_2922;
wire n_2924;
wire n_2925;
wire n_2926;
wire n_2927;
wire n_2929;
wire n_2930;
wire n_2931;
wire n_2932;
wire n_2933;
wire n_2934;
wire n_2935;
wire n_2937;
wire n_2938;
wire n_2939;
wire n_294;
wire n_2940;
wire n_2941;
wire n_2942;
wire n_2943;
wire n_2946;
wire n_2947;
wire n_2948;
wire n_2949;
wire n_2950;
wire n_2951;
wire n_2952;
wire n_2953;
wire n_2954;
wire n_2955;
wire n_2956;
wire n_2957;
wire n_2958;
wire n_2959;
wire n_2960;
wire n_2961;
wire n_2962;
wire n_2963;
wire n_2964;
wire n_2965;
wire n_2966;
wire n_2967;
wire n_2968;
wire n_2969;
wire n_297;
wire n_2970;
wire n_2971;
wire n_2972;
wire n_2973;
wire n_2979;
wire n_298;
wire n_2980;
wire n_2981;
wire n_2982;
wire n_2983;
wire n_2984;
wire n_2986;
wire n_2987;
wire n_2988;
wire n_2989;
wire n_2990;
wire n_2991;
wire n_2992;
wire n_2993;
wire n_2995;
wire n_2996;
wire n_2997;
wire n_2998;
wire n_2999;
wire n_300;
wire n_3000;
wire n_3001;
wire n_3004;
wire n_3005;
wire n_3006;
wire n_3007;
wire n_3008;
wire n_3013;
wire n_3014;
wire n_3015;
wire n_3016;
wire TIMEBOOST_net_14848;
wire n_3018;
wire n_3019;
wire n_302;
wire n_3020;
wire n_3021;
wire n_3022;
wire n_3023;
wire n_3024;
wire n_3025;
wire n_3026;
wire n_3027;
wire n_3028;
wire n_303;
wire n_3030;
wire n_3031;
wire n_3032;
wire n_3033;
wire n_3034;
wire n_3036;
wire n_3037;
wire n_3039;
wire n_304;
wire n_3040;
wire n_3041;
wire n_3042;
wire n_3043;
wire n_3044;
wire n_3045;
wire n_3046;
wire n_3047;
wire n_3048;
wire n_3049;
wire n_3050;
wire n_3051;
wire n_3052;
wire n_3053;
wire n_3054;
wire n_3055;
wire n_3057;
wire n_3058;
wire n_3059;
wire n_306;
wire n_3060;
wire n_3061;
wire n_3062;
wire n_3064;
wire n_3066;
wire n_3068;
wire n_307;
wire n_3070;
wire n_3071;
wire n_3072;
wire n_3073;
wire n_3074;
wire n_3076;
wire n_3077;
wire n_3078;
wire n_3079;
wire n_3080;
wire n_3081;
wire n_3083;
wire n_3084;
wire n_3087;
wire n_3089;
wire n_3090;
wire n_3107;
wire n_3108;
wire n_3109;
wire n_3110;
wire n_3111;
wire n_3112;
wire n_3114;
wire n_3115;
wire n_3116;
wire n_3117;
wire n_3118;
wire n_3119;
wire n_3120;
wire n_3123;
wire n_3125;
wire n_3126;
wire TIMEBOOST_net_22278;
wire n_313;
wire n_3130;
wire n_3131;
wire n_3132;
wire n_3133;
wire n_3134;
wire n_3135;
wire n_3136;
wire n_3137;
wire n_3138;
wire n_3139;
wire n_3140;
wire n_3141;
wire n_3142;
wire n_3147;
wire n_3148;
wire n_3151;
wire n_3152;
wire n_3153;
wire n_3154;
wire n_3156;
wire n_3157;
wire n_3158;
wire n_3159;
wire n_3160;
wire n_3162;
wire n_3163;
wire n_3164;
wire n_3166;
wire n_3167;
wire n_3168;
wire n_3169;
wire n_317;
wire n_3170;
wire n_3171;
wire n_3172;
wire n_3173;
wire n_3174;
wire n_3175;
wire n_3178;
wire n_3179;
wire n_3184;
wire n_3185;
wire n_3189;
wire n_319;
wire n_3190;
wire n_3191;
wire n_3192;
wire n_3193;
wire n_3194;
wire n_3195;
wire n_3196;
wire n_3197;
wire n_3198;
wire n_3199;
wire n_320;
wire n_3200;
wire n_3201;
wire n_3202;
wire n_3203;
wire n_3204;
wire n_3206;
wire n_3209;
wire n_321;
wire n_3210;
wire n_3211;
wire TIMEBOOST_net_23500;
wire TIMEBOOST_net_21215;
wire n_3216;
wire n_3217;
wire n_3219;
wire n_3220;
wire n_3221;
wire n_3222;
wire n_3223;
wire n_3224;
wire n_3226;
wire n_3227;
wire n_3228;
wire n_3229;
wire n_323;
wire n_3231;
wire n_3232;
wire n_3233;
wire n_3235;
wire n_3236;
wire n_3237;
wire n_3238;
wire n_324;
wire n_3241;
wire n_3245;
wire n_3246;
wire n_3247;
wire n_3248;
wire n_325;
wire n_3250;
wire n_3251;
wire n_3252;
wire n_3254;
wire n_3255;
wire n_3256;
wire n_3257;
wire n_3258;
wire n_3259;
wire n_326;
wire n_3260;
wire n_3261;
wire n_3262;
wire n_3265;
wire n_3266;
wire n_3267;
wire n_3268;
wire TIMEBOOST_net_9498;
wire n_3271;
wire n_3273;
wire n_3274;
wire n_3275;
wire n_3276;
wire n_3277;
wire n_3278;
wire n_3279;
wire n_3280;
wire n_3281;
wire n_3282;
wire TIMEBOOST_net_22437;
wire TIMEBOOST_net_21827;
wire TIMEBOOST_net_9606;
wire n_3289;
wire n_329;
wire n_3290;
wire n_3292;
wire n_3293;
wire n_3294;
wire n_3295;
wire n_3296;
wire n_3297;
wire n_3298;
wire n_3301;
wire n_3302;
wire n_3304;
wire n_3305;
wire n_3306;
wire n_331;
wire n_3310;
wire n_3313;
wire n_3314;
wire n_3315;
wire n_3316;
wire n_3317;
wire n_3318;
wire n_3319;
wire n_3320;
wire n_3321;
wire n_3323;
wire n_3324;
wire n_3325;
wire n_3326;
wire n_3327;
wire n_3329;
wire n_333;
wire n_3330;
wire n_3331;
wire n_3332;
wire n_3333;
wire n_3334;
wire n_3335;
wire n_3337;
wire n_3338;
wire n_3339;
wire n_3341;
wire n_3342;
wire n_3344;
wire n_3345;
wire n_3346;
wire n_3347;
wire TIMEBOOST_net_11009;
wire TIMEBOOST_net_11008;
wire n_335;
wire n_3350;
wire n_3351;
wire n_3352;
wire n_3353;
wire n_3354;
wire n_3355;
wire TIMEBOOST_net_16747;
wire n_3357;
wire n_3358;
wire n_3359;
wire n_336;
wire TIMEBOOST_net_17536;
wire n_3361;
wire n_3363;
wire n_3364;
wire n_3365;
wire n_3366;
wire n_3367;
wire n_3368;
wire n_337;
wire n_3370;
wire n_3371;
wire n_3372;
wire n_3373;
wire n_3374;
wire n_3375;
wire n_3376;
wire n_3377;
wire n_3378;
wire n_3379;
wire n_3380;
wire n_3381;
wire n_3384;
wire n_3385;
wire n_3386;
wire n_3387;
wire n_3388;
wire n_3389;
wire n_3390;
wire n_3391;
wire n_3392;
wire n_3393;
wire n_3395;
wire n_3399;
wire n_34;
wire n_340;
wire n_3402;
wire n_3403;
wire n_3404;
wire n_3406;
wire n_3407;
wire n_3408;
wire n_3409;
wire n_341;
wire n_3410;
wire n_3413;
wire n_3415;
wire n_3416;
wire n_3417;
wire n_3419;
wire n_342;
wire n_3420;
wire n_3421;
wire n_3422;
wire n_3423;
wire n_3424;
wire n_3425;
wire n_3428;
wire n_3429;
wire n_343;
wire n_3432;
wire n_3436;
wire n_3437;
wire n_3438;
wire n_3440;
wire n_3443;
wire n_3444;
wire n_3445;
wire n_3446;
wire n_3447;
wire n_3448;
wire n_3449;
wire n_345;
wire n_3450;
wire n_3453;
wire n_3454;
wire n_3455;
wire TIMEBOOST_net_17256;
wire TIMEBOOST_net_16741;
wire n_3462;
wire n_3463;
wire n_3464;
wire n_3465;
wire n_3466;
wire n_3467;
wire n_3468;
wire TIMEBOOST_net_10731;
wire n_3471;
wire n_3472;
wire n_3474;
wire n_3475;
wire n_3476;
wire n_3477;
wire n_3478;
wire n_3479;
wire n_3480;
wire n_3481;
wire TIMEBOOST_net_16695;
wire n_3484;
wire n_3485;
wire n_3486;
wire n_3487;
wire n_3488;
wire n_3489;
wire n_349;
wire n_3490;
wire n_3491;
wire n_3492;
wire n_3493;
wire TIMEBOOST_net_16744;
wire TIMEBOOST_net_16740;
wire n_3496;
wire n_3497;
wire n_3498;
wire n_3499;
wire n_350;
wire n_3501;
wire n_3502;
wire n_3503;
wire n_3504;
wire n_3505;
wire TIMEBOOST_net_20571;
wire TIMEBOOST_net_20580;
wire n_351;
wire n_3510;
wire TIMEBOOST_net_23269;
wire TIMEBOOST_net_13960;
wire TIMEBOOST_net_20576;
wire TIMEBOOST_net_14866;
wire TIMEBOOST_net_21145;
wire TIMEBOOST_net_20954;
wire n_3523;
wire n_3524;
wire TIMEBOOST_net_23252;
wire TIMEBOOST_net_20562;
wire TIMEBOOST_net_20948;
wire TIMEBOOST_net_20945;
wire TIMEBOOST_net_21144;
wire TIMEBOOST_net_20963;
wire TIMEBOOST_net_21139;
wire TIMEBOOST_net_20966;
wire n_354;
wire TIMEBOOST_net_14512;
wire TIMEBOOST_net_21140;
wire TIMEBOOST_net_20962;
wire TIMEBOOST_net_20968;
wire TIMEBOOST_net_22925;
wire TIMEBOOST_net_13957;
wire TIMEBOOST_net_20560;
wire TIMEBOOST_net_20964;
wire TIMEBOOST_net_21121;
wire TIMEBOOST_net_22996;
wire TIMEBOOST_net_21120;
wire TIMEBOOST_net_16723;
wire TIMEBOOST_net_23364;
wire TIMEBOOST_net_8654;
wire TIMEBOOST_net_20848;
wire TIMEBOOST_net_22703;
wire TIMEBOOST_net_20578;
wire n_3568;
wire TIMEBOOST_net_20559;
wire n_357;
wire TIMEBOOST_net_20366;
wire TIMEBOOST_net_20378;
wire TIMEBOOST_net_20581;
wire TIMEBOOST_net_23071;
wire TIMEBOOST_net_20585;
wire TIMEBOOST_net_23365;
wire n_358;
wire TIMEBOOST_net_20959;
wire TIMEBOOST_net_20814;
wire TIMEBOOST_net_21041;
wire TIMEBOOST_net_20952;
wire TIMEBOOST_net_22688;
wire TIMEBOOST_net_22099;
wire TIMEBOOST_net_20950;
wire TIMEBOOST_net_17118;
wire n_3591;
wire n_3592;
wire n_3593;
wire TIMEBOOST_net_20561;
wire TIMEBOOST_net_17547;
wire n_3598;
wire TIMEBOOST_net_20476;
wire n_36;
wire n_360;
wire TIMEBOOST_net_20350;
wire TIMEBOOST_net_23236;
wire TIMEBOOST_net_20410;
wire n_3608;
wire TIMEBOOST_net_20409;
wire n_3616;
wire TIMEBOOST_net_20574;
wire TIMEBOOST_net_20813;
wire n_362;
wire TIMEBOOST_net_20354;
wire TIMEBOOST_net_20980;
wire TIMEBOOST_net_20603;
wire TIMEBOOST_net_22883;
wire n_3627;
wire TIMEBOOST_net_20351;
wire TIMEBOOST_net_20348;
wire TIMEBOOST_net_20485;
wire n_3636;
wire TIMEBOOST_net_20820;
wire n_364;
wire TIMEBOOST_net_23264;
wire TIMEBOOST_net_23459;
wire TIMEBOOST_net_20740;
wire n_3650;
wire TIMEBOOST_net_20582;
wire TIMEBOOST_net_20586;
wire TIMEBOOST_net_20831;
wire n_3655;
wire TIMEBOOST_net_20587;
wire n_366;
wire TIMEBOOST_net_23475;
wire TIMEBOOST_net_20730;
wire TIMEBOOST_net_20715;
wire n_3665;
wire TIMEBOOST_net_21009;
wire n_3667;
wire TIMEBOOST_net_20818;
wire n_3672;
wire TIMEBOOST_net_23503;
wire TIMEBOOST_net_20430;
wire TIMEBOOST_net_20521;
wire n_3677;
wire n_3678;
wire TIMEBOOST_net_20979;
wire TIMEBOOST_net_20520;
wire TIMEBOOST_net_20602;
wire n_369;
wire n_3691;
wire TIMEBOOST_net_20597;
wire TIMEBOOST_net_20353;
wire TIMEBOOST_net_20352;
wire TIMEBOOST_net_21958;
wire n_3697;
wire n_370;
wire TIMEBOOST_net_20748;
wire TIMEBOOST_net_20510;
wire TIMEBOOST_net_23181;
wire TIMEBOOST_net_20827;
wire TIMEBOOST_net_23485;
wire TIMEBOOST_net_20572;
wire TIMEBOOST_net_21137;
wire TIMEBOOST_net_23530;
wire TIMEBOOST_net_20558;
wire TIMEBOOST_net_20738;
wire n_372;
wire n_3721;
wire TIMEBOOST_net_20751;
wire TIMEBOOST_net_20753;
wire TIMEBOOST_net_21296;
wire n_373;
wire TIMEBOOST_net_20594;
wire TIMEBOOST_net_21850;
wire TIMEBOOST_net_20474;
wire TIMEBOOST_net_20544;
wire n_3738;
wire n_3739;
wire n_374;
wire n_3740;
wire n_3741;
wire TIMEBOOST_net_20734;
wire n_3744;
wire TIMEBOOST_net_20270;
wire TIMEBOOST_net_20846;
wire n_3747;
wire n_3749;
wire n_375;
wire TIMEBOOST_net_21813;
wire n_3752;
wire n_3754;
wire n_3755;
wire TIMEBOOST_net_20573;
wire TIMEBOOST_net_20414;
wire TIMEBOOST_net_20823;
wire n_376;
wire n_3760;
wire n_3761;
wire TIMEBOOST_net_20413;
wire n_3763;
wire n_3764;
wire n_3765;
wire n_3768;
wire n_377;
wire n_3770;
wire n_3774;
wire TIMEBOOST_net_20554;
wire n_3777;
wire TIMEBOOST_net_23219;
wire TIMEBOOST_net_23172;
wire n_378;
wire n_3780;
wire n_3781;
wire n_3783;
wire n_3785;
wire n_3786;
wire TIMEBOOST_net_23180;
wire TIMEBOOST_net_20824;
wire n_3791;
wire n_3792;
wire n_3794;
wire n_3795;
wire n_3796;
wire n_3797;
wire n_3798;
wire n_3799;
wire n_38;
wire n_3800;
wire n_3805;
wire n_3806;
wire n_3807;
wire n_3808;
wire n_3809;
wire n_3810;
wire n_3811;
wire n_3812;
wire TIMEBOOST_net_16669;
wire TIMEBOOST_net_13350;
wire n_3815;
wire TIMEBOOST_net_23132;
wire TIMEBOOST_net_20509;
wire n_382;
wire TIMEBOOST_net_20475;
wire TIMEBOOST_net_23142;
wire TIMEBOOST_net_21203;
wire TIMEBOOST_net_17365;
wire n_3827;
wire n_3830;
wire n_3832;
wire TIMEBOOST_net_23489;
wire n_3838;
wire n_384;
wire n_3840;
wire TIMEBOOST_net_20513;
wire TIMEBOOST_net_20491;
wire n_3843;
wire n_3844;
wire n_3846;
wire TIMEBOOST_net_23158;
wire n_3848;
wire n_385;
wire n_3850;
wire n_3852;
wire n_3853;
wire TIMEBOOST_net_16008;
wire n_3856;
wire n_3857;
wire n_3858;
wire n_386;
wire n_3861;
wire n_3863;
wire TIMEBOOST_net_15942;
wire n_3869;
wire TIMEBOOST_net_20636;
wire n_3872;
wire TIMEBOOST_net_13089;
wire n_3875;
wire n_3876;
wire TIMEBOOST_net_20495;
wire n_3879;
wire n_3880;
wire n_3885;
wire n_3886;
wire n_3887;
wire n_389;
wire n_3890;
wire TIMEBOOST_net_17360;
wire TIMEBOOST_net_17482;
wire TIMEBOOST_net_20638;
wire TIMEBOOST_net_23393;
wire n_3900;
wire TIMEBOOST_net_17483;
wire n_3904;
wire n_3905;
wire n_3906;
wire n_4369;
wire n_391;
wire n_3910;
wire n_3912;
wire n_3917;
wire TIMEBOOST_net_23170;
wire n_3921;
wire n_3922;
wire n_3923;
wire n_3925;
wire TIMEBOOST_net_21210;
wire n_3929;
wire n_393;
wire n_3930;
wire n_3931;
wire TIMEBOOST_net_8580;
wire TIMEBOOST_net_22138;
wire n_3939;
wire TIMEBOOST_net_17434;
wire TIMEBOOST_net_15102;
wire n_3947;
wire n_3948;
wire TIMEBOOST_net_13525;
wire n_395;
wire TIMEBOOST_net_17128;
wire n_3951;
wire n_3954;
wire n_3955;
wire n_3957;
wire n_3958;
wire TIMEBOOST_net_21211;
wire n_396;
wire n_3960;
wire TIMEBOOST_net_20171;
wire n_3963;
wire TIMEBOOST_net_13512;
wire n_3968;
wire n_3969;
wire n_397;
wire n_3970;
wire n_3972;
wire TIMEBOOST_net_21212;
wire TIMEBOOST_net_21214;
wire TIMEBOOST_net_20160;
wire n_3978;
wire TIMEBOOST_net_20174;
wire n_398;
wire TIMEBOOST_net_21038;
wire TIMEBOOST_net_17429;
wire n_3982;
wire TIMEBOOST_net_17431;
wire TIMEBOOST_net_20534;
wire n_3988;
wire n_3991;
wire n_3993;
wire TIMEBOOST_net_20882;
wire n_3995;
wire TIMEBOOST_net_20178;
wire TIMEBOOST_net_14925;
wire n_40;
wire TIMEBOOST_net_13524;
wire n_4001;
wire TIMEBOOST_net_17436;
wire TIMEBOOST_net_20970;
wire n_4005;
wire TIMEBOOST_net_17435;
wire TIMEBOOST_net_17437;
wire n_4009;
wire n_401;
wire n_4010;
wire TIMEBOOST_net_17433;
wire n_4013;
wire n_4014;
wire TIMEBOOST_net_17430;
wire TIMEBOOST_net_17548;
wire n_4024;
wire n_4025;
wire n_4026;
wire TIMEBOOST_net_12478;
wire n_4029;
wire n_4031;
wire n_4032;
wire n_4033;
wire TIMEBOOST_net_20176;
wire TIMEBOOST_net_17124;
wire n_4037;
wire n_4038;
wire TIMEBOOST_net_17131;
wire n_404;
wire TIMEBOOST_net_15552;
wire n_4043;
wire n_4044;
wire n_4045;
wire n_4046;
wire n_4047;
wire TIMEBOOST_net_21060;
wire n_405;
wire n_4051;
wire n_4053;
wire TIMEBOOST_net_17129;
wire TIMEBOOST_net_21213;
wire n_4056;
wire n_4057;
wire TIMEBOOST_net_20175;
wire n_4061;
wire n_4062;
wire TIMEBOOST_net_21216;
wire n_4064;
wire n_4065;
wire n_4067;
wire TIMEBOOST_net_20172;
wire n_4069;
wire n_407;
wire TIMEBOOST_net_23315;
wire n_4072;
wire n_4073;
wire n_4074;
wire n_4075;
wire TIMEBOOST_net_23397;
wire n_4077;
wire n_4078;
wire n_408;
wire n_4080;
wire n_4084;
wire n_4085;
wire n_4086;
wire n_4088;
wire n_409;
wire n_4090;
wire n_4092;
wire n_4093;
wire n_4095;
wire n_4096;
wire n_4097;
wire n_4098;
wire n_4100;
wire n_4101;
wire n_4102;
wire n_4103;
wire n_4104;
wire n_4105;
wire n_4106;
wire n_4107;
wire n_4108;
wire n_4109;
wire n_411;
wire n_4111;
wire n_4112;
wire n_4113;
wire n_4114;
wire n_4115;
wire n_4119;
wire n_412;
wire n_4123;
wire n_4125;
wire n_413;
wire n_4130;
wire n_4131;
wire n_4132;
wire n_4134;
wire n_4135;
wire n_4136;
wire n_4137;
wire n_4138;
wire n_4140;
wire n_4142;
wire n_4143;
wire n_4144;
wire n_4145;
wire n_4146;
wire n_4149;
wire n_4151;
wire n_4152;
wire n_4153;
wire n_4154;
wire n_4155;
wire TIMEBOOST_net_20953;
wire n_4157;
wire n_4158;
wire n_416;
wire n_4160;
wire n_4161;
wire n_4162;
wire n_4165;
wire n_4167;
wire n_4168;
wire n_4169;
wire n_4170;
wire n_4171;
wire n_4172;
wire n_4177;
wire TIMEBOOST_net_11425;
wire n_4188;
wire n_419;
wire TIMEBOOST_net_11013;
wire TIMEBOOST_net_23396;
wire TIMEBOOST_net_16751;
wire TIMEBOOST_net_21118;
wire TIMEBOOST_net_11011;
wire n_4196;
wire n_4197;
wire n_4198;
wire TIMEBOOST_net_20691;
wire n_42;
wire n_420;
wire n_4200;
wire n_4201;
wire n_4202;
wire TIMEBOOST_net_11288;
wire n_4205;
wire n_4206;
wire n_4207;
wire n_4208;
wire n_4209;
wire n_4210;
wire n_4211;
wire n_4212;
wire n_4213;
wire n_4214;
wire n_4216;
wire TIMEBOOST_net_20949;
wire n_4222;
wire TIMEBOOST_net_20856;
wire n_4225;
wire TIMEBOOST_net_23150;
wire TIMEBOOST_net_23383;
wire TIMEBOOST_net_16431;
wire TIMEBOOST_net_20843;
wire TIMEBOOST_net_23359;
wire TIMEBOOST_net_23522;
wire TIMEBOOST_net_20761;
wire TIMEBOOST_net_13959;
wire n_424;
wire TIMEBOOST_net_20967;
wire TIMEBOOST_net_20965;
wire TIMEBOOST_net_23120;
wire n_425;
wire TIMEBOOST_net_13958;
wire TIMEBOOST_net_21138;
wire TIMEBOOST_net_21131;
wire TIMEBOOST_net_21142;
wire n_4261;
wire TIMEBOOST_net_20863;
wire n_4265;
wire TIMEBOOST_net_20955;
wire TIMEBOOST_net_17525;
wire n_4273;
wire TIMEBOOST_net_20930;
wire TIMEBOOST_net_23516;
wire n_4280;
wire TIMEBOOST_net_20739;
wire TIMEBOOST_net_20957;
wire TIMEBOOST_net_23526;
wire TIMEBOOST_net_23520;
wire TIMEBOOST_net_15875;
wire n_430;
wire n_4302;
wire TIMEBOOST_net_20722;
wire TIMEBOOST_net_23501;
wire TIMEBOOST_net_23495;
wire TIMEBOOST_net_20754;
wire TIMEBOOST_net_20596;
wire n_4312;
wire TIMEBOOST_net_23258;
wire TIMEBOOST_net_20765;
wire TIMEBOOST_net_21190;
wire TIMEBOOST_net_20847;
wire n_432;
wire TIMEBOOST_net_21722;
wire TIMEBOOST_net_20666;
wire n_4323;
wire TIMEBOOST_net_17439;
wire n_4327;
wire TIMEBOOST_net_20763;
wire n_433;
wire n_4330;
wire TIMEBOOST_net_20727;
wire TIMEBOOST_net_20604;
wire TIMEBOOST_net_20468;
wire TIMEBOOST_net_20720;
wire TIMEBOOST_net_20663;
wire n_434;
wire TIMEBOOST_net_20477;
wire TIMEBOOST_net_341;
wire n_4343;
wire TIMEBOOST_net_23507;
wire n_4345;
wire TIMEBOOST_net_23476;
wire n_4359;
wire TIMEBOOST_net_21037;
wire n_4349;
wire TIMEBOOST_net_23462;
wire TIMEBOOST_net_20465;
wire TIMEBOOST_net_20762;
wire TIMEBOOST_net_20764;
wire n_4357;
wire n_4358;
wire TIMEBOOST_net_20725;
wire n_436;
wire TIMEBOOST_net_23474;
wire TIMEBOOST_net_16975;
wire TIMEBOOST_net_21675;
wire TIMEBOOST_net_7592;
wire TIMEBOOST_net_21014;
wire TIMEBOOST_net_21135;
wire TIMEBOOST_net_23514;
wire TIMEBOOST_net_22792;
wire n_4382;
wire TIMEBOOST_net_23540;
wire TIMEBOOST_net_20757;
wire TIMEBOOST_net_20718;
wire TIMEBOOST_net_20759;
wire n_439;
wire TIMEBOOST_net_13136;
wire n_4392;
wire TIMEBOOST_net_23499;
wire n_4394;
wire TIMEBOOST_net_20969;
wire n_4396;
wire TIMEBOOST_net_20600;
wire TIMEBOOST_net_23306;
wire n_4399;
wire n_440;
wire TIMEBOOST_net_20598;
wire n_4402;
wire n_4403;
wire TIMEBOOST_net_20756;
wire n_4406;
wire n_4409;
wire n_4410;
wire TIMEBOOST_net_20732;
wire TIMEBOOST_net_20737;
wire TIMEBOOST_net_20736;
wire TIMEBOOST_net_20731;
wire TIMEBOOST_net_20728;
wire n_4417;
wire TIMEBOOST_net_23508;
wire TIMEBOOST_net_21141;
wire TIMEBOOST_net_13249;
wire TIMEBOOST_net_8653;
wire n_4429;
wire TIMEBOOST_net_23477;
wire n_4437;
wire n_4438;
wire TIMEBOOST_net_17438;
wire n_4442;
wire n_4444;
wire TIMEBOOST_net_20601;
wire n_4447;
wire TIMEBOOST_net_20972;
wire n_4450;
wire n_4452;
wire TIMEBOOST_net_20768;
wire n_4454;
wire n_4456;
wire TIMEBOOST_net_20726;
wire TIMEBOOST_net_20332;
wire n_4460;
wire TIMEBOOST_net_20721;
wire TIMEBOOST_net_20263;
wire TIMEBOOST_net_20767;
wire n_4465;
wire n_4466;
wire TIMEBOOST_net_20479;
wire TIMEBOOST_net_20758;
wire n_447;
wire n_4470;
wire n_4472;
wire n_4473;
wire TIMEBOOST_net_20667;
wire n_4476;
wire n_4477;
wire n_4479;
wire n_4480;
wire TIMEBOOST_net_20478;
wire n_4482;
wire TIMEBOOST_net_20755;
wire TIMEBOOST_net_23152;
wire TIMEBOOST_net_23137;
wire n_4488;
wire n_4490;
wire TIMEBOOST_net_23136;
wire n_4493;
wire TIMEBOOST_net_21133;
wire n_4495;
wire TIMEBOOST_net_20766;
wire n_4497;
wire n_4498;
wire TIMEBOOST_net_21028;
wire TIMEBOOST_net_23154;
wire n_4501;
wire n_4504;
wire n_4505;
wire TIMEBOOST_net_23148;
wire n_4508;
wire n_4509;
wire n_4510;
wire n_4511;
wire n_4512;
wire n_4513;
wire n_4514;
wire n_4516;
wire n_4517;
wire n_4519;
wire n_4520;
wire n_4521;
wire n_4522;
wire n_4523;
wire n_4524;
wire n_4527;
wire n_4528;
wire n_4532;
wire n_4533;
wire n_4534;
wire n_4535;
wire n_4536;
wire n_4537;
wire n_454;
wire n_4591;
wire n_4592;
wire n_4594;
wire TIMEBOOST_net_17522;
wire n_4598;
wire n_46;
wire n_4601;
wire n_4603;
wire n_4605;
wire n_4607;
wire TIMEBOOST_net_10722;
wire TIMEBOOST_net_17313;
wire n_4610;
wire n_4611;
wire TIMEBOOST_net_22256;
wire n_4614;
wire n_4616;
wire n_4617;
wire n_4618;
wire n_4619;
wire n_4621;
wire n_4623;
wire n_4625;
wire n_4627;
wire n_4628;
wire n_4629;
wire n_4630;
wire n_4631;
wire n_4632;
wire n_4633;
wire n_4634;
wire n_4635;
wire n_4636;
wire n_4637;
wire n_4638;
wire n_4639;
wire n_4641;
wire n_4642;
wire n_4644;
wire n_4645;
wire TIMEBOOST_net_21130;
wire n_4647;
wire n_4649;
wire n_4652;
wire n_4654;
wire n_4655;
wire TIMEBOOST_net_21134;
wire n_4658;
wire n_4659;
wire n_4660;
wire n_4661;
wire n_4662;
wire n_4663;
wire n_4664;
wire n_4666;
wire n_4667;
wire n_4668;
wire n_4669;
wire n_4671;
wire n_4672;
wire n_4674;
wire n_4675;
wire n_4677;
wire n_4679;
wire n_4680;
wire n_4681;
wire n_4683;
wire n_4685;
wire n_4686;
wire TIMEBOOST_net_11012;
wire n_4688;
wire TIMEBOOST_net_11010;
wire n_4691;
wire n_4692;
wire n_4693;
wire n_4694;
wire n_4695;
wire n_4696;
wire n_4697;
wire TIMEBOOST_net_16748;
wire n_4699;
wire n_47;
wire n_4700;
wire n_4702;
wire n_4703;
wire n_4704;
wire TIMEBOOST_net_23394;
wire TIMEBOOST_net_16746;
wire n_4707;
wire n_4708;
wire n_471;
wire n_4711;
wire n_4712;
wire n_4713;
wire n_4714;
wire n_4715;
wire TIMEBOOST_net_320;
wire n_4717;
wire n_4718;
wire n_4719;
wire n_4720;
wire n_4721;
wire n_4722;
wire n_4723;
wire n_4725;
wire n_4726;
wire n_4727;
wire n_4728;
wire n_4729;
wire n_4730;
wire n_4732;
wire n_4733;
wire n_4734;
wire n_4735;
wire n_4736;
wire n_4737;
wire n_4739;
wire n_4740;
wire n_4741;
wire n_4743;
wire TIMEBOOST_net_22195;
wire n_4746;
wire TIMEBOOST_net_13704;
wire TIMEBOOST_net_16966;
wire TIMEBOOST_net_13601;
wire TIMEBOOST_net_12762;
wire TIMEBOOST_net_20349;
wire TIMEBOOST_net_13225;
wire TIMEBOOST_net_8231;
wire g62021_db;
wire TIMEBOOST_net_23321;
wire g61989_db;
wire TIMEBOOST_net_7473;
wire TIMEBOOST_net_21720;
wire TIMEBOOST_net_13597;
wire TIMEBOOST_net_8236;
wire TIMEBOOST_net_16844;
wire TIMEBOOST_net_13593;
wire n_3269;
wire TIMEBOOST_net_7472;
wire TIMEBOOST_net_13594;
wire TIMEBOOST_net_237;
wire n_4778;
wire TIMEBOOST_net_13595;
wire n_4780;
wire n_4781;
wire n_4782;
wire n_4783;
wire n_4784;
wire n_4785;
wire n_4786;
wire n_4792;
wire n_4793;
wire n_4795;
wire n_4796;
wire n_4797;
wire n_4798;
wire n_4799;
wire n_4800;
wire n_4802;
wire n_4803;
wire n_4806;
wire n_4807;
wire n_4808;
wire n_4809;
wire n_4811;
wire n_4812;
wire n_4813;
wire n_4814;
wire n_4815;
wire n_4816;
wire n_4818;
wire n_4819;
wire n_4820;
wire n_4822;
wire n_4823;
wire n_4824;
wire n_4825;
wire n_4826;
wire n_4828;
wire n_4830;
wire n_4831;
wire n_4832;
wire n_4833;
wire n_4834;
wire n_4835;
wire n_4836;
wire n_4837;
wire n_4838;
wire n_4839;
wire n_4840;
wire n_4841;
wire n_4842;
wire n_4843;
wire n_4844;
wire n_4845;
wire n_4846;
wire n_4847;
wire n_4848;
wire n_4849;
wire n_4851;
wire n_4853;
wire n_4855;
wire n_4856;
wire n_4857;
wire n_4858;
wire n_4859;
wire n_4860;
wire n_4861;
wire n_4862;
wire n_4863;
wire n_4864;
wire n_4866;
wire n_4867;
wire n_4868;
wire n_4869;
wire n_4870;
wire n_4871;
wire n_4872;
wire n_4873;
wire n_4874;
wire n_4875;
wire n_4877;
wire n_4878;
wire n_4879;
wire n_4880;
wire n_4881;
wire n_4883;
wire n_4884;
wire TIMEBOOST_net_17035;
wire n_4886;
wire TIMEBOOST_net_23245;
wire n_4889;
wire n_4890;
wire n_4891;
wire n_4892;
wire TIMEBOOST_net_17545;
wire n_4894;
wire n_4895;
wire n_4896;
wire n_4897;
wire n_4899;
wire n_4900;
wire n_4901;
wire n_4902;
wire n_4903;
wire n_4904;
wire n_4905;
wire n_4906;
wire n_4907;
wire n_4908;
wire n_4909;
wire n_4911;
wire n_4912;
wire n_4913;
wire n_4914;
wire n_4915;
wire n_4917;
wire n_4918;
wire n_4920;
wire n_4922;
wire n_4924;
wire n_4926;
wire n_4928;
wire n_4930;
wire n_4932;
wire n_4934;
wire n_4936;
wire n_4939;
wire n_4941;
wire n_4943;
wire n_4945;
wire n_4947;
wire n_4949;
wire n_4951;
wire n_4953;
wire n_4955;
wire n_4957;
wire n_4959;
wire n_4961;
wire n_4963;
wire n_4965;
wire n_4968;
wire n_497;
wire n_4970;
wire n_4973;
wire n_4975;
wire n_4978;
wire n_4980;
wire n_4982;
wire n_4984;
wire n_4986;
wire n_4988;
wire n_4991;
wire n_4993;
wire n_4996;
wire n_4999;
wire n_50;
wire n_5001;
wire n_5003;
wire n_5006;
wire n_5009;
wire n_5012;
wire n_5014;
wire n_5016;
wire n_5018;
wire n_5021;
wire n_5023;
wire n_5025;
wire n_5027;
wire n_5029;
wire n_5031;
wire n_5033;
wire n_5036;
wire n_5038;
wire n_504;
wire n_5040;
wire n_5042;
wire n_5044;
wire n_5046;
wire n_5048;
wire n_5050;
wire n_5052;
wire n_5054;
wire n_5056;
wire n_5058;
wire n_5060;
wire n_5062;
wire n_5064;
wire n_5066;
wire n_5068;
wire n_5071;
wire n_5074;
wire n_5076;
wire n_5078;
wire n_5080;
wire n_5082;
wire n_5084;
wire n_5086;
wire n_5088;
wire n_5090;
wire n_5092;
wire n_5094;
wire n_5096;
wire n_5098;
wire n_5100;
wire n_5102;
wire n_5104;
wire n_5106;
wire n_5108;
wire n_5110;
wire n_5112;
wire n_5114;
wire n_5116;
wire n_5118;
wire n_512;
wire n_5120;
wire n_5122;
wire n_5124;
wire n_5126;
wire n_5128;
wire n_513;
wire n_5130;
wire n_5132;
wire n_5134;
wire n_5136;
wire n_5138;
wire n_5140;
wire n_5143;
wire n_5146;
wire n_5149;
wire n_5151;
wire n_5153;
wire n_5156;
wire n_5158;
wire n_5161;
wire n_5163;
wire n_5166;
wire n_5168;
wire n_5170;
wire n_5172;
wire n_5174;
wire n_5176;
wire n_5179;
wire n_518;
wire n_5181;
wire n_5183;
wire n_5185;
wire n_5188;
wire n_519;
wire n_5190;
wire n_5192;
wire n_5194;
wire n_5196;
wire n_5198;
wire n_520;
wire n_5200;
wire n_5203;
wire n_5205;
wire n_5207;
wire n_521;
wire n_5210;
wire n_5212;
wire n_5214;
wire n_5216;
wire n_5218;
wire n_522;
wire n_5221;
wire n_5223;
wire n_5225;
wire n_5227;
wire n_5228;
wire n_5229;
wire n_523;
wire n_5230;
wire n_5232;
wire n_5235;
wire n_5237;
wire n_524;
wire n_5240;
wire n_5242;
wire n_5244;
wire n_5246;
wire n_5248;
wire n_525;
wire n_5251;
wire n_5253;
wire n_5255;
wire n_5258;
wire n_526;
wire n_5260;
wire n_5263;
wire n_5265;
wire n_5267;
wire n_5269;
wire n_527;
wire n_5272;
wire n_5275;
wire n_5277;
wire n_5279;
wire n_528;
wire n_5281;
wire n_5283;
wire n_5285;
wire n_5288;
wire n_529;
wire n_5290;
wire n_5293;
wire n_5296;
wire n_5298;
wire n_530;
wire n_5300;
wire n_5303;
wire n_5305;
wire n_5308;
wire n_531;
wire n_5311;
wire n_5313;
wire n_5315;
wire n_5318;
wire n_532;
wire n_5320;
wire n_5323;
wire n_5325;
wire n_5327;
wire n_533;
wire n_5330;
wire n_5332;
wire n_5335;
wire n_5337;
wire n_5339;
wire n_534;
wire n_5342;
wire n_5345;
wire n_5347;
wire n_5349;
wire n_535;
wire n_5351;
wire n_5354;
wire n_5356;
wire n_5358;
wire n_536;
wire n_5361;
wire n_5363;
wire n_5366;
wire n_5368;
wire n_5371;
wire n_5373;
wire n_5376;
wire n_5378;
wire n_538;
wire n_5380;
wire n_5383;
wire n_5386;
wire n_5388;
wire n_539;
wire n_5391;
wire n_5393;
wire n_5396;
wire n_5399;
wire n_540;
wire n_5402;
wire n_5404;
wire n_5406;
wire n_5409;
wire n_541;
wire n_5412;
wire n_5414;
wire n_5416;
wire n_5418;
wire n_5421;
wire n_5424;
wire n_5427;
wire n_5429;
wire n_5431;
wire n_5433;
wire n_5435;
wire n_5438;
wire n_544;
wire n_5441;
wire n_5444;
wire n_5446;
wire n_5448;
wire n_545;
wire n_5450;
wire n_5452;
wire n_5454;
wire n_5456;
wire n_5458;
wire n_546;
wire n_5461;
wire n_5463;
wire n_5465;
wire n_5467;
wire n_547;
wire n_5470;
wire n_5472;
wire n_5474;
wire n_5476;
wire n_5478;
wire n_5481;
wire n_5483;
wire n_5486;
wire n_5489;
wire n_549;
wire n_5491;
wire n_5493;
wire n_5495;
wire n_5497;
wire n_5499;
wire n_550;
wire n_5501;
wire n_5503;
wire n_5505;
wire n_5507;
wire n_5509;
wire n_551;
wire n_5511;
wire n_5513;
wire n_5515;
wire n_5517;
wire n_5519;
wire n_5521;
wire n_5523;
wire n_5526;
wire n_5528;
wire n_5531;
wire n_5534;
wire n_5537;
wire n_5539;
wire n_554;
wire n_5541;
wire n_5543;
wire n_5545;
wire n_5546;
wire n_5547;
wire n_5548;
wire n_5549;
wire n_5552;
wire n_5553;
wire n_5554;
wire n_5555;
wire n_5556;
wire n_5557;
wire n_5558;
wire n_5559;
wire n_5561;
wire n_5563;
wire n_5565;
wire n_5566;
wire n_5567;
wire n_5568;
wire n_5569;
wire n_5570;
wire n_5571;
wire n_5572;
wire n_5573;
wire n_5574;
wire n_5575;
wire n_5576;
wire n_5577;
wire n_5578;
wire n_5579;
wire n_558;
wire n_5580;
wire n_5581;
wire n_5582;
wire n_5583;
wire n_5585;
wire n_5587;
wire n_5588;
wire n_5589;
wire n_559;
wire n_5591;
wire n_5592;
wire n_5593;
wire n_5594;
wire n_5595;
wire n_5597;
wire n_5598;
wire n_560;
wire n_5600;
wire n_5601;
wire n_5603;
wire n_5604;
wire n_5606;
wire n_5607;
wire n_5608;
wire n_5609;
wire n_561;
wire n_5611;
wire n_5612;
wire n_5614;
wire n_5616;
wire n_5617;
wire n_5618;
wire n_5619;
wire n_562;
wire n_5620;
wire n_5622;
wire n_5623;
wire n_5625;
wire n_5626;
wire n_5627;
wire n_5628;
wire n_563;
wire n_5630;
wire n_5631;
wire n_5632;
wire n_5633;
wire n_5634;
wire n_5635;
wire n_5636;
wire n_5637;
wire n_5638;
wire n_5639;
wire n_564;
wire n_5640;
wire n_5641;
wire n_5642;
wire n_5643;
wire n_5644;
wire TIMEBOOST_net_10977;
wire n_5646;
wire n_5648;
wire n_5649;
wire n_565;
wire n_5650;
wire n_5651;
wire n_5652;
wire n_5654;
wire n_5655;
wire n_5656;
wire n_5657;
wire n_5658;
wire n_566;
wire n_5660;
wire n_5662;
wire n_5663;
wire n_5664;
wire n_5666;
wire n_5668;
wire n_5669;
wire n_567;
wire n_5670;
wire n_5672;
wire n_5673;
wire n_5675;
wire n_5676;
wire n_5678;
wire n_5679;
wire n_568;
wire n_5681;
wire n_5682;
wire n_5684;
wire n_5686;
wire n_5687;
wire n_5688;
wire n_5689;
wire n_5691;
wire n_5694;
wire n_5696;
wire n_5699;
wire n_57;
wire n_5701;
wire n_5702;
wire n_5703;
wire n_5704;
wire n_5705;
wire n_5707;
wire n_5708;
wire n_5709;
wire n_5710;
wire n_5712;
wire n_5713;
wire n_5716;
wire n_5717;
wire n_5718;
wire n_5722;
wire n_5723;
wire n_5724;
wire n_5725;
wire n_5728;
wire TIMEBOOST_net_14587;
wire n_573;
wire n_5730;
wire n_5731;
wire n_5732;
wire n_5733;
wire n_5735;
wire n_5736;
wire n_5737;
wire n_5739;
wire n_574;
wire n_5740;
wire n_5741;
wire n_5742;
wire n_5743;
wire n_5744;
wire n_5745;
wire n_5747;
wire n_5748;
wire TIMEBOOST_net_21330;
wire n_5750;
wire n_5751;
wire TIMEBOOST_net_21342;
wire n_5753;
wire n_5754;
wire n_5755;
wire n_5757;
wire n_5758;
wire TIMEBOOST_net_17081;
wire n_5763;
wire n_5766;
wire n_5768;
wire n_5769;
wire n_5770;
wire n_5772;
wire n_5774;
wire n_5776;
wire n_5778;
wire n_5780;
wire n_5782;
wire n_5784;
wire n_5786;
wire n_5788;
wire n_5790;
wire n_5792;
wire n_5794;
wire n_5796;
wire n_5798;
wire n_580;
wire n_5800;
wire n_5802;
wire n_5804;
wire n_5806;
wire n_5808;
wire n_581;
wire n_5810;
wire n_5812;
wire n_5814;
wire n_5816;
wire n_5819;
wire n_582;
wire n_5822;
wire n_5824;
wire n_5827;
wire n_583;
wire n_5830;
wire n_5833;
wire n_5836;
wire n_5838;
wire n_584;
wire n_5840;
wire n_5842;
wire n_5844;
wire n_5846;
wire n_5848;
wire n_585;
wire n_5850;
wire n_5852;
wire n_5854;
wire n_5856;
wire n_5858;
wire n_586;
wire n_5860;
wire n_5862;
wire n_5864;
wire n_5866;
wire n_5868;
wire n_587;
wire n_5870;
wire n_5872;
wire n_5874;
wire n_5876;
wire n_5878;
wire n_588;
wire n_5880;
wire n_5882;
wire n_5884;
wire n_5886;
wire n_5888;
wire n_5890;
wire n_5892;
wire n_5894;
wire n_5896;
wire n_5898;
wire n_5900;
wire n_5902;
wire n_5904;
wire n_5906;
wire n_5908;
wire n_5910;
wire n_5912;
wire n_5914;
wire n_5916;
wire n_5918;
wire n_592;
wire n_5920;
wire n_5922;
wire n_5924;
wire n_5926;
wire n_5928;
wire n_593;
wire n_5930;
wire n_5932;
wire n_5934;
wire n_5936;
wire n_5938;
wire n_594;
wire n_5940;
wire n_5942;
wire n_5944;
wire n_5946;
wire n_5948;
wire n_595;
wire n_5950;
wire n_5952;
wire n_5954;
wire n_5956;
wire n_5958;
wire n_596;
wire n_5960;
wire n_5962;
wire n_5964;
wire n_5966;
wire n_5967;
wire n_5969;
wire n_597;
wire n_5971;
wire n_5973;
wire n_5975;
wire n_5977;
wire n_5979;
wire n_598;
wire n_5981;
wire n_5983;
wire n_5985;
wire n_5987;
wire n_5989;
wire n_599;
wire n_5991;
wire n_5993;
wire n_5995;
wire n_5997;
wire n_5999;
wire n_6;
wire n_600;
wire n_6001;
wire n_6003;
wire n_6005;
wire n_6007;
wire n_6009;
wire n_601;
wire n_6011;
wire n_6013;
wire n_6015;
wire n_6017;
wire n_6019;
wire n_602;
wire n_6021;
wire n_6023;
wire n_6025;
wire n_6027;
wire n_6029;
wire n_603;
wire n_6031;
wire n_6033;
wire n_6035;
wire n_6037;
wire n_6039;
wire n_604;
wire n_6040;
wire n_6041;
wire n_6043;
wire n_6045;
wire n_6047;
wire n_6049;
wire n_605;
wire n_6051;
wire n_6053;
wire n_6054;
wire n_6056;
wire n_6058;
wire n_606;
wire n_6060;
wire n_6061;
wire n_6063;
wire n_6065;
wire n_6067;
wire n_6069;
wire n_607;
wire n_6071;
wire n_6073;
wire n_6075;
wire n_6077;
wire n_6079;
wire n_6081;
wire n_6083;
wire n_6085;
wire n_6087;
wire n_6089;
wire n_609;
wire n_6091;
wire n_6093;
wire n_6095;
wire n_6097;
wire n_6099;
wire n_61;
wire n_610;
wire n_6101;
wire n_6103;
wire n_6105;
wire n_6107;
wire n_6109;
wire n_611;
wire n_6111;
wire n_6112;
wire n_6115;
wire n_6117;
wire n_6119;
wire n_612;
wire n_6121;
wire n_6123;
wire n_6125;
wire n_6127;
wire n_6129;
wire n_613;
wire n_6132;
wire n_6135;
wire n_6136;
wire n_6138;
wire n_614;
wire n_6140;
wire n_6142;
wire n_6144;
wire n_6146;
wire n_6148;
wire n_615;
wire n_6150;
wire n_6152;
wire n_6154;
wire n_6156;
wire n_6158;
wire n_616;
wire n_6160;
wire n_6162;
wire n_6164;
wire n_6166;
wire n_6168;
wire n_617;
wire n_6171;
wire n_6173;
wire n_6175;
wire n_6177;
wire n_6179;
wire n_6181;
wire n_6184;
wire n_6186;
wire n_6189;
wire n_6191;
wire n_6193;
wire n_6195;
wire n_6196;
wire n_6199;
wire n_620;
wire n_6200;
wire n_6201;
wire n_6204;
wire n_6206;
wire n_6208;
wire n_621;
wire n_6211;
wire n_6213;
wire n_6216;
wire n_6218;
wire n_622;
wire n_6221;
wire n_6223;
wire n_6226;
wire n_6228;
wire n_623;
wire n_6230;
wire n_6231;
wire n_6232;
wire n_6234;
wire n_6235;
wire n_6238;
wire n_624;
wire n_6240;
wire n_6243;
wire n_6246;
wire n_6249;
wire n_625;
wire n_6252;
wire n_6254;
wire n_6257;
wire n_6259;
wire n_626;
wire n_6261;
wire n_6264;
wire n_6266;
wire n_6268;
wire n_627;
wire n_6271;
wire n_6273;
wire n_6276;
wire n_6278;
wire n_6281;
wire n_6284;
wire n_6286;
wire n_6287;
wire n_6289;
wire n_629;
wire n_6292;
wire n_6295;
wire n_6297;
wire n_6298;
wire n_6301;
wire n_6303;
wire n_6305;
wire n_6308;
wire n_6311;
wire n_6313;
wire n_6315;
wire n_6318;
wire n_6319;
wire n_6321;
wire n_6323;
wire n_6325;
wire n_6327;
wire n_6329;
wire n_6331;
wire n_6333;
wire n_6334;
wire n_6335;
wire n_6337;
wire n_6338;
wire n_6340;
wire n_6342;
wire n_6344;
wire n_6345;
wire n_6347;
wire n_6348;
wire n_6350;
wire n_6353;
wire n_6355;
wire n_6356;
wire n_6358;
wire n_6361;
wire n_6364;
wire n_6366;
wire n_6369;
wire n_6371;
wire n_6372;
wire n_6373;
wire n_6374;
wire n_6376;
wire n_6379;
wire n_6382;
wire n_6384;
wire n_6386;
wire n_6388;
wire n_639;
wire n_6390;
wire n_6391;
wire n_6393;
wire n_6395;
wire n_6398;
wire n_640;
wire n_6400;
wire n_6402;
wire n_6405;
wire n_6407;
wire n_641;
wire n_6410;
wire n_6413;
wire n_6415;
wire n_6417;
wire n_642;
wire n_6420;
wire n_6423;
wire n_6425;
wire n_6427;
wire n_643;
wire n_6430;
wire n_6431;
wire n_6433;
wire n_6435;
wire n_6436;
wire n_6438;
wire n_6440;
wire n_6443;
wire n_6446;
wire n_6448;
wire n_645;
wire n_6451;
wire n_6453;
wire n_6456;
wire n_6458;
wire n_646;
wire n_6461;
wire n_6463;
wire n_6465;
wire n_6468;
wire n_6470;
wire n_6473;
wire n_6475;
wire n_6477;
wire n_648;
wire n_6480;
wire n_6483;
wire n_6485;
wire n_6488;
wire n_649;
wire n_6490;
wire n_6493;
wire n_6495;
wire n_6498;
wire n_65;
wire n_650;
wire n_6501;
wire n_6504;
wire n_6506;
wire n_6509;
wire n_6512;
wire n_6514;
wire n_6516;
wire n_6518;
wire n_652;
wire n_6521;
wire n_6523;
wire n_6526;
wire n_6528;
wire n_653;
wire n_6530;
wire n_6532;
wire n_6534;
wire n_6536;
wire n_6538;
wire n_6541;
wire n_6543;
wire n_6546;
wire n_6548;
wire n_655;
wire n_6550;
wire n_6553;
wire n_6554;
wire n_6556;
wire n_6558;
wire n_656;
wire n_6561;
wire n_6563;
wire n_6566;
wire n_6567;
wire n_6569;
wire n_657;
wire n_6572;
wire n_6575;
wire n_6578;
wire n_658;
wire n_6580;
wire n_6582;
wire n_6585;
wire n_6587;
wire n_6589;
wire n_659;
wire n_6592;
wire n_6594;
wire n_6596;
wire n_6598;
wire n_660;
wire n_6601;
wire n_6603;
wire n_6605;
wire n_6607;
wire n_661;
wire n_6610;
wire n_6613;
wire n_6615;
wire n_6617;
wire n_662;
wire n_6620;
wire n_6621;
wire n_6623;
wire n_6624;
wire n_6626;
wire n_6629;
wire n_663;
wire n_6631;
wire n_6634;
wire n_6636;
wire n_6639;
wire n_664;
wire n_6641;
wire n_6644;
wire n_6645;
wire n_6647;
wire n_6649;
wire n_665;
wire n_6651;
wire n_6654;
wire n_6657;
wire n_6659;
wire n_666;
wire n_6662;
wire n_6665;
wire n_6668;
wire n_667;
wire n_6670;
wire n_6672;
wire n_6674;
wire n_6676;
wire n_6678;
wire n_668;
wire n_6680;
wire n_6682;
wire n_6684;
wire n_6686;
wire n_6689;
wire n_669;
wire n_6691;
wire n_6693;
wire n_6695;
wire n_6697;
wire n_6699;
wire n_67;
wire n_670;
wire n_6701;
wire n_6703;
wire n_6705;
wire n_6707;
wire n_6709;
wire n_671;
wire n_6712;
wire n_6714;
wire n_6716;
wire n_6718;
wire n_672;
wire n_6720;
wire n_6722;
wire n_6724;
wire n_6726;
wire n_6729;
wire n_673;
wire n_6731;
wire n_6733;
wire n_6735;
wire n_6738;
wire n_674;
wire n_6741;
wire n_6743;
wire n_6745;
wire n_6747;
wire n_6749;
wire n_675;
wire n_6752;
wire n_6754;
wire n_6757;
wire n_6759;
wire n_676;
wire n_6761;
wire n_6763;
wire n_6766;
wire n_6768;
wire n_677;
wire n_6770;
wire n_6772;
wire n_6774;
wire n_6776;
wire n_6778;
wire n_678;
wire n_6781;
wire n_6783;
wire n_6785;
wire n_6788;
wire n_6789;
wire n_6791;
wire n_6793;
wire n_6795;
wire n_6797;
wire n_6799;
wire n_6801;
wire n_6804;
wire n_6806;
wire n_6809;
wire n_681;
wire n_6812;
wire n_6814;
wire n_6816;
wire n_6819;
wire n_6821;
wire n_6824;
wire n_6826;
wire n_6828;
wire n_6830;
wire n_6833;
wire n_6835;
wire n_6837;
wire n_6840;
wire n_6842;
wire n_6845;
wire n_6847;
wire n_6849;
wire n_6851;
wire n_6853;
wire n_6855;
wire n_6857;
wire n_6859;
wire n_6861;
wire n_6863;
wire n_6865;
wire n_6867;
wire n_6868;
wire n_6869;
wire n_6871;
wire n_6872;
wire n_6875;
wire n_6876;
wire n_6878;
wire n_6880;
wire n_6883;
wire n_6885;
wire n_6886;
wire n_6887;
wire n_6889;
wire n_689;
wire n_6892;
wire n_6895;
wire n_6897;
wire n_6898;
wire n_6900;
wire n_6902;
wire n_6903;
wire n_6905;
wire n_6908;
wire n_691;
wire n_6910;
wire n_6911;
wire n_6913;
wire n_6915;
wire n_6917;
wire n_6919;
wire n_692;
wire n_6920;
wire n_6922;
wire n_6924;
wire n_6926;
wire n_6929;
wire n_6932;
wire n_6934;
wire n_6935;
wire n_6937;
wire n_6940;
wire n_6941;
wire n_6942;
wire n_6943;
wire n_6944;
wire n_6946;
wire n_6948;
wire n_695;
wire n_6951;
wire n_6953;
wire n_6956;
wire n_6958;
wire n_696;
wire n_6961;
wire n_6963;
wire n_6965;
wire n_6967;
wire n_6969;
wire n_6971;
wire n_6973;
wire n_6975;
wire n_6977;
wire n_6978;
wire n_6980;
wire n_6982;
wire n_6983;
wire n_6984;
wire n_6985;
wire n_6986;
wire n_6987;
wire n_6989;
wire n_6991;
wire n_6992;
wire n_6993;
wire n_6994;
wire n_6995;
wire n_6996;
wire n_6997;
wire n_6998;
wire n_6999;
wire n_700;
wire n_7000;
wire n_7001;
wire n_7002;
wire n_7003;
wire n_7004;
wire n_7005;
wire n_7006;
wire n_7007;
wire n_7008;
wire n_7009;
wire n_7010;
wire n_7011;
wire n_7012;
wire n_7013;
wire n_7014;
wire n_7015;
wire n_7016;
wire n_7018;
wire n_7019;
wire n_7027;
wire n_7028;
wire n_7029;
wire n_703;
wire n_7030;
wire n_7031;
wire n_7032;
wire n_7033;
wire n_7038;
wire n_7039;
wire n_7040;
wire n_7043;
wire n_7044;
wire n_7045;
wire n_7046;
wire n_7047;
wire n_7048;
wire n_7049;
wire n_705;
wire n_7050;
wire n_7051;
wire n_7052;
wire n_7053;
wire n_7054;
wire n_7055;
wire n_7056;
wire n_7057;
wire n_7058;
wire n_7059;
wire n_7060;
wire n_7061;
wire n_7062;
wire n_7063;
wire n_7064;
wire n_7065;
wire n_7066;
wire n_7067;
wire n_7068;
wire n_7069;
wire n_707;
wire n_7070;
wire n_7071;
wire n_7072;
wire n_7073;
wire n_7074;
wire n_7075;
wire TIMEBOOST_net_11210;
wire n_7078;
wire n_7079;
wire n_708;
wire n_7080;
wire n_7081;
wire n_7082;
wire n_7083;
wire n_7084;
wire TIMEBOOST_net_20386;
wire TIMEBOOST_net_16514;
wire TIMEBOOST_net_17104;
wire TIMEBOOST_net_17455;
wire n_709;
wire n_7091;
wire n_7092;
wire n_7093;
wire n_7094;
wire n_7095;
wire n_7096;
wire n_7102;
wire n_7108;
wire n_711;
wire n_7110;
wire n_7112;
wire n_7114;
wire n_7115;
wire n_7117;
wire n_7119;
wire n_7121;
wire n_7122;
wire n_7123;
wire n_7125;
wire n_7126;
wire n_7128;
wire n_713;
wire n_7130;
wire n_7132;
wire n_7134;
wire n_7135;
wire n_7136;
wire n_7137;
wire n_7139;
wire n_7141;
wire n_7143;
wire n_7145;
wire n_7147;
wire n_7149;
wire n_715;
wire n_7151;
wire n_7153;
wire n_7155;
wire n_7157;
wire n_7159;
wire n_716;
wire n_7161;
wire n_7163;
wire n_7165;
wire n_7168;
wire n_7171;
wire n_7174;
wire n_7177;
wire n_7180;
wire n_7182;
wire n_7185;
wire n_7187;
wire n_7189;
wire n_7191;
wire n_7193;
wire n_7195;
wire n_7197;
wire n_72;
wire n_7200;
wire n_7203;
wire n_7205;
wire n_7207;
wire n_7209;
wire n_721;
wire n_7210;
wire n_7211;
wire n_7212;
wire n_7213;
wire n_7214;
wire n_7216;
wire n_7218;
wire n_722;
wire n_7220;
wire TIMEBOOST_net_17551;
wire TIMEBOOST_net_20161;
wire n_7226;
wire n_7227;
wire n_7228;
wire n_7229;
wire n_7231;
wire n_7232;
wire n_7233;
wire n_7234;
wire n_7235;
wire n_7236;
wire n_7237;
wire n_7238;
wire n_7239;
wire n_7240;
wire n_7241;
wire n_7242;
wire n_7243;
wire n_7244;
wire n_7245;
wire n_7246;
wire n_7247;
wire n_7248;
wire n_7249;
wire n_725;
wire n_7250;
wire n_7251;
wire n_7252;
wire n_7253;
wire n_7254;
wire n_7255;
wire n_7256;
wire n_7257;
wire n_7258;
wire n_7259;
wire n_7260;
wire n_7261;
wire n_7262;
wire n_7263;
wire n_7264;
wire n_7265;
wire n_7266;
wire n_7267;
wire n_7268;
wire n_7269;
wire n_727;
wire n_7270;
wire n_7271;
wire n_7272;
wire n_7273;
wire n_7274;
wire n_7275;
wire n_7276;
wire n_7277;
wire n_7278;
wire n_7279;
wire n_7280;
wire n_7281;
wire n_7282;
wire n_7283;
wire n_7284;
wire n_7285;
wire n_7286;
wire n_7287;
wire n_7288;
wire n_7289;
wire n_729;
wire n_7290;
wire n_7291;
wire n_7293;
wire n_7294;
wire n_7295;
wire n_7296;
wire n_7297;
wire n_7298;
wire n_730;
wire n_7300;
wire n_7307;
wire n_7308;
wire n_7309;
wire n_731;
wire n_7310;
wire n_7311;
wire n_7312;
wire n_7313;
wire n_7315;
wire n_7316;
wire n_7317;
wire TIMEBOOST_net_20983;
wire n_7320;
wire n_7321;
wire n_7322;
wire n_7324;
wire n_7325;
wire TIMEBOOST_net_767;
wire n_7329;
wire n_733;
wire n_7330;
wire n_7333;
wire TIMEBOOST_net_22438;
wire TIMEBOOST_net_14340;
wire n_7338;
wire n_7339;
wire n_734;
wire n_7341;
wire TIMEBOOST_net_11329;
wire n_7350;
wire n_736;
wire n_7362;
wire n_7364;
wire n_7366;
wire n_7368;
wire n_7369;
wire n_737;
wire n_7371;
wire n_7373;
wire n_7374;
wire n_7375;
wire n_7377;
wire n_7379;
wire n_738;
wire n_7381;
wire n_7383;
wire n_7385;
wire n_7386;
wire n_7387;
wire n_7388;
wire n_739;
wire n_7390;
wire n_7392;
wire n_7393;
wire n_7396;
wire n_7397;
wire n_7398;
wire n_7399;
wire n_74;
wire n_740;
wire n_7400;
wire n_7401;
wire n_7404;
wire n_7405;
wire n_7406;
wire n_7407;
wire n_7408;
wire n_7409;
wire n_741;
wire n_7410;
wire n_7411;
wire n_7412;
wire n_7413;
wire n_7414;
wire n_7415;
wire n_7416;
wire n_7417;
wire n_7418;
wire n_7419;
wire n_742;
wire n_7420;
wire n_7421;
wire n_7422;
wire n_7423;
wire n_7424;
wire n_7425;
wire n_7426;
wire n_7427;
wire n_7428;
wire n_7429;
wire n_743;
wire n_7430;
wire n_7431;
wire n_7432;
wire n_7433;
wire n_7434;
wire n_7435;
wire n_7436;
wire n_7437;
wire n_7438;
wire n_7439;
wire n_744;
wire n_7440;
wire n_7442;
wire n_7443;
wire n_7444;
wire n_7445;
wire n_7446;
wire n_7447;
wire n_7448;
wire n_7449;
wire n_745;
wire n_7450;
wire n_7451;
wire n_7452;
wire n_7453;
wire n_7454;
wire n_7455;
wire n_7456;
wire n_7457;
wire n_7458;
wire n_7459;
wire n_746;
wire n_7460;
wire n_7461;
wire n_7462;
wire n_7463;
wire n_7464;
wire n_7465;
wire n_7466;
wire n_7467;
wire n_7468;
wire n_7469;
wire n_747;
wire n_7470;
wire n_7472;
wire n_7473;
wire n_7474;
wire n_7475;
wire n_7476;
wire n_7477;
wire n_7478;
wire n_7479;
wire n_748;
wire n_7480;
wire n_7481;
wire n_7482;
wire n_7483;
wire n_7484;
wire n_7485;
wire n_7486;
wire n_7487;
wire n_7488;
wire n_7489;
wire n_7490;
wire n_7491;
wire n_7492;
wire n_7493;
wire n_7494;
wire n_7495;
wire n_7496;
wire n_7497;
wire n_7498;
wire n_7499;
wire n_75;
wire n_7500;
wire n_7504;
wire n_7505;
wire n_7508;
wire n_7509;
wire n_7510;
wire n_7511;
wire n_7512;
wire n_7513;
wire n_7514;
wire n_7515;
wire n_7516;
wire n_7517;
wire n_7518;
wire n_7519;
wire n_7521;
wire n_7522;
wire n_7523;
wire n_7524;
wire n_7525;
wire n_7527;
wire n_7528;
wire n_7529;
wire n_7530;
wire n_7531;
wire n_7532;
wire n_7534;
wire n_7535;
wire n_7538;
wire n_7539;
wire n_7540;
wire n_7541;
wire n_7542;
wire n_7543;
wire n_7544;
wire n_7547;
wire n_7548;
wire n_7550;
wire n_7551;
wire n_7552;
wire n_7557;
wire n_7558;
wire n_7559;
wire n_7560;
wire n_7561;
wire n_7562;
wire n_7564;
wire n_7565;
wire n_7567;
wire n_7568;
wire n_7569;
wire n_7571;
wire n_7574;
wire n_7575;
wire n_7576;
wire n_7577;
wire n_7578;
wire n_7579;
wire n_7580;
wire n_7581;
wire n_7582;
wire n_7583;
wire n_7584;
wire n_7585;
wire n_7586;
wire n_7587;
wire n_7588;
wire n_7589;
wire n_7590;
wire n_7591;
wire n_7592;
wire n_7593;
wire n_7594;
wire n_7595;
wire n_7596;
wire n_7597;
wire n_7598;
wire n_7599;
wire n_76;
wire n_7600;
wire n_7601;
wire n_7602;
wire n_7603;
wire n_7604;
wire n_7605;
wire n_7606;
wire n_7607;
wire n_7608;
wire n_7609;
wire n_7610;
wire n_7611;
wire n_7612;
wire n_7613;
wire n_7614;
wire n_7615;
wire n_7616;
wire n_7617;
wire n_7618;
wire n_7619;
wire n_7620;
wire n_7621;
wire n_7622;
wire n_7624;
wire n_7625;
wire n_7626;
wire n_7627;
wire n_7628;
wire n_7629;
wire n_763;
wire n_7630;
wire n_7631;
wire n_7632;
wire n_7633;
wire n_7634;
wire n_7635;
wire n_7636;
wire n_7637;
wire n_7638;
wire n_7639;
wire n_7640;
wire n_7642;
wire n_7643;
wire n_7645;
wire n_7646;
wire n_7647;
wire n_7648;
wire n_7649;
wire n_7650;
wire n_7651;
wire n_7652;
wire n_7653;
wire n_7654;
wire n_7655;
wire n_7656;
wire n_7657;
wire n_7658;
wire n_7661;
wire n_7663;
wire n_7664;
wire n_7665;
wire n_7666;
wire n_7667;
wire n_7669;
wire n_7671;
wire n_7672;
wire n_7673;
wire n_7677;
wire n_7679;
wire n_7681;
wire n_7683;
wire n_7684;
wire n_7685;
wire n_7687;
wire n_7689;
wire n_7692;
wire n_7694;
wire n_7695;
wire n_7697;
wire n_7698;
wire n_7699;
wire n_7701;
wire n_7702;
wire n_7704;
wire n_7705;
wire n_7706;
wire n_7707;
wire n_7708;
wire n_7709;
wire n_7712;
wire n_7714;
wire n_7715;
wire n_7716;
wire n_7717;
wire n_7718;
wire n_7719;
wire n_7720;
wire n_7721;
wire n_7722;
wire n_7723;
wire n_7724;
wire n_7725;
wire n_7726;
wire TIMEBOOST_net_21359;
wire n_7731;
wire n_7733;
wire n_7734;
wire n_7735;
wire n_7737;
wire n_7738;
wire n_7739;
wire n_7740;
wire n_7742;
wire n_7743;
wire n_7744;
wire n_7745;
wire n_7746;
wire n_7747;
wire n_7749;
wire n_7750;
wire n_7751;
wire n_7752;
wire n_7753;
wire n_7754;
wire n_7755;
wire n_7756;
wire n_7757;
wire n_7759;
wire n_7760;
wire n_7761;
wire n_7762;
wire n_7764;
wire n_7766;
wire n_7767;
wire n_7768;
wire n_7769;
wire n_7771;
wire n_7773;
wire n_7774;
wire n_7776;
wire n_7777;
wire n_7779;
wire n_7780;
wire n_7781;
wire n_7782;
wire n_7783;
wire n_7785;
wire n_7786;
wire n_7787;
wire n_7788;
wire n_7789;
wire n_779;
wire n_7790;
wire n_7791;
wire n_7792;
wire n_7793;
wire n_7794;
wire n_7795;
wire n_7796;
wire n_7797;
wire n_7798;
wire n_7799;
wire n_7800;
wire n_7801;
wire n_7802;
wire n_7803;
wire n_7804;
wire n_7805;
wire n_7806;
wire n_7807;
wire n_7808;
wire n_7809;
wire n_7810;
wire n_7811;
wire n_7812;
wire n_7813;
wire n_7814;
wire n_7815;
wire n_7816;
wire n_7817;
wire n_7818;
wire n_7819;
wire n_7820;
wire n_7821;
wire n_7822;
wire n_7823;
wire n_7824;
wire n_7826;
wire n_7828;
wire n_783;
wire n_7830;
wire n_7833;
wire n_7835;
wire n_7836;
wire n_7838;
wire n_784;
wire n_7840;
wire n_7842;
wire n_7844;
wire n_7845;
wire n_7847;
wire n_7849;
wire n_785;
wire n_7851;
wire n_7853;
wire n_7855;
wire n_7857;
wire n_7859;
wire n_7861;
wire n_7863;
wire n_7865;
wire n_7867;
wire n_7869;
wire n_7871;
wire n_7873;
wire n_7875;
wire n_7877;
wire n_7879;
wire n_7881;
wire n_7883;
wire n_7885;
wire n_7887;
wire n_7889;
wire n_7891;
wire n_7893;
wire n_7895;
wire n_7897;
wire n_7899;
wire n_790;
wire n_7901;
wire n_7903;
wire n_7905;
wire n_7907;
wire n_7909;
wire n_791;
wire n_7911;
wire n_7913;
wire n_7915;
wire n_7917;
wire n_7919;
wire n_7921;
wire n_7923;
wire n_7925;
wire n_7927;
wire n_7929;
wire n_7931;
wire n_7933;
wire n_7935;
wire n_7937;
wire n_7939;
wire n_7941;
wire n_7943;
wire n_7945;
wire n_7947;
wire n_7949;
wire n_7951;
wire n_7953;
wire n_7955;
wire n_7957;
wire n_7959;
wire n_7961;
wire n_7963;
wire n_7965;
wire n_7967;
wire n_7969;
wire n_7971;
wire n_7973;
wire n_7975;
wire n_7977;
wire n_7979;
wire n_798;
wire n_7981;
wire n_7983;
wire n_7985;
wire n_7987;
wire n_7989;
wire n_7991;
wire n_7993;
wire n_7995;
wire n_7997;
wire n_7999;
wire n_8001;
wire n_8003;
wire n_8005;
wire n_8007;
wire n_8009;
wire n_8012;
wire n_8014;
wire n_8017;
wire n_8019;
wire n_802;
wire n_8021;
wire n_8024;
wire n_8027;
wire n_8030;
wire n_8032;
wire n_8034;
wire n_8036;
wire n_8039;
wire n_8041;
wire n_8044;
wire n_8047;
wire n_8049;
wire n_8052;
wire n_8054;
wire n_8056;
wire n_8059;
wire n_8060;
wire n_8062;
wire n_8064;
wire n_8066;
wire n_8068;
wire n_8069;
wire n_8071;
wire n_8073;
wire n_8076;
wire n_8079;
wire TIMEBOOST_net_20169;
wire n_8082;
wire n_8084;
wire n_8087;
wire n_8089;
wire n_8092;
wire n_8094;
wire n_8097;
wire n_8100;
wire n_8102;
wire n_8105;
wire n_8107;
wire n_8109;
wire n_8111;
wire n_8114;
wire n_8116;
wire n_8118;
wire n_8119;
wire n_812;
wire n_8121;
wire n_8123;
wire n_8125;
wire n_8128;
wire n_813;
wire n_8130;
wire n_8132;
wire n_8135;
wire n_8137;
wire n_8139;
wire n_8140;
wire n_8142;
wire n_8144;
wire n_8147;
wire n_815;
wire n_8150;
wire n_8152;
wire n_8154;
wire n_8157;
wire n_8159;
wire n_816;
wire n_8161;
wire n_8163;
wire n_8166;
wire n_8168;
wire n_817;
wire n_8171;
wire n_8173;
wire n_8175;
wire n_8176;
wire n_8178;
wire n_8180;
wire n_8182;
wire n_8184;
wire n_8186;
wire n_8189;
wire n_819;
wire n_8191;
wire n_8193;
wire n_8196;
wire n_8198;
wire n_8200;
wire n_8203;
wire n_8205;
wire n_8208;
wire n_8210;
wire n_8213;
wire n_8215;
wire n_8218;
wire n_8220;
wire n_8223;
wire n_8226;
wire n_8229;
wire n_8231;
wire n_8232;
wire n_8234;
wire n_8236;
wire n_8239;
wire n_824;
wire n_8241;
wire n_8244;
wire n_8246;
wire n_8248;
wire n_8251;
wire n_8253;
wire n_8255;
wire n_8258;
wire n_826;
wire n_8260;
wire n_8262;
wire n_8264;
wire n_8267;
wire n_8269;
wire n_8271;
wire n_8272;
wire n_8274;
wire n_8277;
wire n_8279;
wire n_8281;
wire n_8283;
wire n_8285;
wire n_8288;
wire n_829;
wire n_8291;
wire n_8293;
wire n_8295;
wire n_8297;
wire n_8299;
wire n_83;
wire n_8302;
wire n_8304;
wire n_8307;
wire n_8309;
wire n_8311;
wire n_8313;
wire n_8316;
wire n_8319;
wire n_832;
wire n_8321;
wire n_8323;
wire n_8325;
wire n_8327;
wire n_8329;
wire n_833;
wire n_8331;
wire n_8333;
wire n_8335;
wire n_8337;
wire n_8339;
wire n_8341;
wire n_8344;
wire n_8346;
wire n_8349;
wire n_8351;
wire n_8353;
wire n_8355;
wire n_8358;
wire n_836;
wire n_8360;
wire n_8362;
wire n_8364;
wire n_8366;
wire n_8368;
wire n_837;
wire n_8371;
wire n_8373;
wire n_8376;
wire n_8379;
wire n_838;
wire n_8382;
wire n_8384;
wire n_8387;
wire n_8389;
wire n_839;
wire n_8391;
wire n_8393;
wire n_8395;
wire n_8397;
wire n_84;
wire n_840;
wire n_8400;
wire n_8402;
wire n_8404;
wire n_8406;
wire n_8407;
wire n_8409;
wire n_841;
wire n_8411;
wire n_8413;
wire n_8415;
wire n_8417;
wire n_8419;
wire n_842;
wire n_8421;
wire n_8423;
wire n_8426;
wire n_8428;
wire n_843;
wire n_8430;
wire n_8431;
wire n_8432;
wire n_8433;
wire n_8434;
wire n_8436;
wire n_8437;
wire n_8438;
wire n_8439;
wire n_844;
wire n_8440;
wire n_8441;
wire n_8442;
wire n_8444;
wire n_8445;
wire n_8446;
wire n_8447;
wire n_8448;
wire n_8449;
wire n_845;
wire n_8450;
wire n_8451;
wire n_8452;
wire n_8453;
wire n_8454;
wire n_8455;
wire n_8456;
wire n_8457;
wire n_8458;
wire n_8459;
wire n_8460;
wire n_8461;
wire n_8462;
wire n_8463;
wire n_8464;
wire n_8465;
wire n_8466;
wire n_8467;
wire n_8468;
wire n_8469;
wire n_847;
wire n_8470;
wire n_8472;
wire n_8474;
wire n_8476;
wire n_8477;
wire n_8478;
wire n_8480;
wire n_8481;
wire n_8482;
wire n_8483;
wire n_8484;
wire n_8485;
wire n_8486;
wire n_8487;
wire n_8488;
wire n_8489;
wire n_849;
wire n_8492;
wire n_8493;
wire n_8494;
wire n_8495;
wire n_8496;
wire n_8498;
wire n_85;
wire n_850;
wire TIMEBOOST_net_11487;
wire n_8501;
wire n_8502;
wire n_8503;
wire n_8504;
wire n_8505;
wire n_8506;
wire n_8508;
wire n_8509;
wire n_851;
wire n_8510;
wire n_8511;
wire n_8512;
wire n_8513;
wire n_8514;
wire n_8515;
wire n_8516;
wire n_8517;
wire n_8518;
wire n_8519;
wire n_852;
wire n_8520;
wire n_8521;
wire n_8522;
wire n_8523;
wire n_8524;
wire n_8525;
wire n_8526;
wire n_8527;
wire n_8528;
wire n_8529;
wire n_853;
wire n_8530;
wire n_8531;
wire TIMEBOOST_net_13587;
wire n_8535;
wire n_8538;
wire TIMEBOOST_net_14808;
wire n_8540;
wire n_8541;
wire n_8542;
wire n_8547;
wire n_8548;
wire n_8549;
wire n_855;
wire n_8550;
wire n_8551;
wire n_8552;
wire n_8553;
wire n_8554;
wire n_8555;
wire n_8556;
wire n_8557;
wire n_8558;
wire n_8559;
wire n_8560;
wire n_8561;
wire n_8562;
wire n_8563;
wire n_8564;
wire n_8565;
wire n_8566;
wire n_8567;
wire n_8568;
wire n_8569;
wire n_8571;
wire n_8572;
wire n_8573;
wire n_8574;
wire n_8575;
wire n_8576;
wire n_8579;
wire n_858;
wire n_8582;
wire n_8583;
wire n_8585;
wire n_8588;
wire n_8589;
wire n_8590;
wire n_8591;
wire n_8595;
wire n_8596;
wire n_8597;
wire n_8598;
wire n_8601;
wire n_8602;
wire n_8603;
wire n_8604;
wire n_8605;
wire n_8606;
wire n_8607;
wire n_8609;
wire n_861;
wire n_8611;
wire n_8613;
wire n_8615;
wire n_8616;
wire n_8617;
wire n_8618;
wire n_8619;
wire n_8620;
wire n_8621;
wire n_8622;
wire n_8623;
wire n_8624;
wire n_8625;
wire n_8626;
wire n_8627;
wire n_8628;
wire n_8629;
wire n_863;
wire n_8630;
wire n_8631;
wire n_8632;
wire n_8633;
wire n_8634;
wire n_8635;
wire n_8636;
wire n_8637;
wire n_8638;
wire n_864;
wire n_8640;
wire n_8641;
wire n_8642;
wire n_8643;
wire n_8644;
wire n_8645;
wire n_8646;
wire n_8647;
wire n_8648;
wire n_8649;
wire n_865;
wire n_8650;
wire n_8651;
wire n_8652;
wire TIMEBOOST_net_23358;
wire n_8655;
wire n_8656;
wire n_8657;
wire n_8658;
wire n_8659;
wire n_866;
wire n_8660;
wire n_8661;
wire n_8662;
wire n_8664;
wire n_8665;
wire n_8668;
wire n_8669;
wire n_867;
wire n_8672;
wire n_8673;
wire n_8674;
wire n_8675;
wire n_8676;
wire n_8677;
wire n_868;
wire n_8680;
wire n_8682;
wire n_8686;
wire n_8687;
wire n_8688;
wire n_869;
wire n_8692;
wire n_8693;
wire n_8694;
wire n_8695;
wire n_8697;
wire n_8699;
wire n_870;
wire n_8701;
wire n_8703;
wire n_8705;
wire n_8707;
wire n_8708;
wire n_8709;
wire n_871;
wire n_8711;
wire n_8712;
wire n_8713;
wire n_8714;
wire n_8716;
wire n_8717;
wire n_872;
wire n_8721;
wire n_8723;
wire n_8724;
wire n_8725;
wire n_8726;
wire n_8727;
wire n_8728;
wire n_8730;
wire n_8731;
wire n_8732;
wire n_8733;
wire n_8734;
wire n_874;
wire TIMEBOOST_net_10377;
wire TIMEBOOST_net_10314;
wire TIMEBOOST_net_10378;
wire n_8745;
wire n_8747;
wire n_8749;
wire n_875;
wire n_8750;
wire n_8751;
wire n_8752;
wire TIMEBOOST_net_16378;
wire n_8757;
wire n_8759;
wire n_876;
wire n_8760;
wire n_8765;
wire n_877;
wire n_878;
wire n_8780;
wire n_8782;
wire n_8784;
wire n_879;
wire n_8790;
wire n_8792;
wire n_8794;
wire TIMEBOOST_net_10056;
wire n_8796;
wire n_880;
wire n_8800;
wire n_8801;
wire n_881;
wire n_8818;
wire n_8819;
wire n_882;
wire n_8820;
wire n_883;
wire n_8831;
wire n_8832;
wire TIMEBOOST_net_16783;
wire TIMEBOOST_net_16784;
wire TIMEBOOST_net_16785;
wire TIMEBOOST_net_16786;
wire TIMEBOOST_net_23494;
wire n_884;
wire TIMEBOOST_net_23528;
wire n_8842;
wire n_8843;
wire n_8846;
wire n_8847;
wire n_8848;
wire n_8849;
wire n_885;
wire n_8850;
wire n_8851;
wire n_8852;
wire n_8853;
wire n_8854;
wire n_8855;
wire n_8857;
wire n_8859;
wire n_886;
wire n_8860;
wire n_8861;
wire n_8863;
wire n_8864;
wire n_8866;
wire n_8867;
wire n_887;
wire n_8871;
wire n_8872;
wire n_8874;
wire n_8875;
wire n_8876;
wire n_8877;
wire n_8879;
wire n_888;
wire n_8880;
wire n_8884;
wire n_8887;
wire n_8888;
wire n_8889;
wire n_889;
wire n_8890;
wire n_8892;
wire n_8896;
wire n_8897;
wire n_8898;
wire n_8899;
wire n_890;
wire n_8900;
wire n_8902;
wire n_8904;
wire n_8906;
wire n_8908;
wire n_891;
wire n_8910;
wire n_8912;
wire n_8914;
wire n_8916;
wire n_8917;
wire n_8919;
wire n_892;
wire n_8920;
wire n_8921;
wire n_8924;
wire n_8926;
wire n_8927;
wire n_8928;
wire n_893;
wire n_8932;
wire n_8934;
wire n_8935;
wire n_8939;
wire n_894;
wire n_8940;
wire n_8941;
wire n_8943;
wire n_8944;
wire n_8945;
wire n_8946;
wire n_8947;
wire n_8949;
wire n_895;
wire n_8950;
wire TIMEBOOST_net_14149;
wire TIMEBOOST_net_10293;
wire n_8953;
wire n_8954;
wire n_8955;
wire n_8957;
wire n_8959;
wire n_896;
wire n_8960;
wire n_8961;
wire n_8962;
wire n_8963;
wire n_8964;
wire n_8965;
wire n_8966;
wire n_8967;
wire n_8968;
wire n_8969;
wire n_897;
wire n_8970;
wire n_8971;
wire n_8973;
wire n_8975;
wire n_8977;
wire n_8979;
wire n_898;
wire n_8981;
wire n_8983;
wire n_8986;
wire n_8989;
wire n_899;
wire TIMEBOOST_net_21051;
wire TIMEBOOST_net_17481;
wire n_8993;
wire TIMEBOOST_net_17432;
wire TIMEBOOST_net_12949;
wire n_8996;
wire n_8997;
wire TIMEBOOST_net_21967;
wire n_9;
wire n_900;
wire TIMEBOOST_net_12513;
wire n_9001;
wire n_9002;
wire n_9003;
wire n_9004;
wire TIMEBOOST_net_23483;
wire n_9007;
wire n_9008;
wire n_9009;
wire n_901;
wire n_9011;
wire n_9012;
wire TIMEBOOST_net_14414;
wire TIMEBOOST_net_23478;
wire n_9017;
wire TIMEBOOST_net_13694;
wire TIMEBOOST_net_21439;
wire n_902;
wire n_9020;
wire n_9021;
wire n_9022;
wire n_9024;
wire n_9025;
wire n_9026;
wire n_9028;
wire TIMEBOOST_net_23468;
wire n_903;
wire TIMEBOOST_net_23416;
wire n_9034;
wire n_9035;
wire TIMEBOOST_net_17094;
wire TIMEBOOST_net_17244;
wire n_904;
wire TIMEBOOST_net_13098;
wire n_9041;
wire n_9045;
wire n_9046;
wire TIMEBOOST_net_12576;
wire TIMEBOOST_net_13130;
wire n_9049;
wire n_905;
wire n_9050;
wire TIMEBOOST_net_12414;
wire n_9053;
wire n_9054;
wire TIMEBOOST_net_13113;
wire n_9057;
wire n_9059;
wire n_906;
wire n_9060;
wire n_9061;
wire TIMEBOOST_net_13117;
wire n_9064;
wire TIMEBOOST_net_12426;
wire n_9068;
wire n_9069;
wire n_907;
wire TIMEBOOST_net_12447;
wire n_9071;
wire n_9072;
wire n_9073;
wire TIMEBOOST_net_20139;
wire TIMEBOOST_net_23349;
wire n_9076;
wire n_9077;
wire TIMEBOOST_net_12451;
wire TIMEBOOST_net_17480;
wire n_908;
wire TIMEBOOST_net_23443;
wire n_9081;
wire n_9082;
wire TIMEBOOST_net_12420;
wire n_9085;
wire n_9086;
wire TIMEBOOST_net_12444;
wire TIMEBOOST_net_13118;
wire n_9089;
wire n_909;
wire n_9090;
wire TIMEBOOST_net_12422;
wire n_9093;
wire n_9094;
wire n_9095;
wire TIMEBOOST_net_13111;
wire n_9097;
wire n_9098;
wire TIMEBOOST_net_21449;
wire n_910;
wire TIMEBOOST_net_21825;
wire n_9102;
wire TIMEBOOST_net_12448;
wire TIMEBOOST_net_13097;
wire n_9105;
wire n_9106;
wire TIMEBOOST_net_21472;
wire TIMEBOOST_net_15039;
wire TIMEBOOST_net_21822;
wire n_911;
wire n_9110;
wire TIMEBOOST_net_12746;
wire n_9112;
wire n_9114;
wire n_9115;
wire n_9116;
wire n_9118;
wire TIMEBOOST_net_12547;
wire n_912;
wire n_9120;
wire TIMEBOOST_net_12549;
wire n_9122;
wire n_9123;
wire n_9124;
wire n_9125;
wire n_9126;
wire TIMEBOOST_net_12544;
wire TIMEBOOST_net_13112;
wire n_9129;
wire n_913;
wire n_9130;
wire TIMEBOOST_net_12541;
wire n_9134;
wire TIMEBOOST_net_17130;
wire TIMEBOOST_net_17242;
wire TIMEBOOST_net_21084;
wire TIMEBOOST_net_21976;
wire n_914;
wire n_9140;
wire TIMEBOOST_net_14276;
wire n_9143;
wire n_9144;
wire n_9145;
wire n_9146;
wire n_915;
wire n_9152;
wire n_9153;
wire n_9154;
wire n_9155;
wire n_916;
wire n_9160;
wire n_9163;
wire n_9168;
wire n_917;
wire n_9170;
wire n_9171;
wire n_9172;
wire n_9173;
wire n_9174;
wire n_9175;
wire n_9176;
wire n_9177;
wire n_9178;
wire n_9179;
wire n_918;
wire n_9180;
wire n_9181;
wire n_9182;
wire n_9183;
wire n_9184;
wire n_9185;
wire n_9187;
wire n_9188;
wire n_9189;
wire n_919;
wire n_9191;
wire n_9192;
wire n_9194;
wire n_9197;
wire n_9198;
wire n_9199;
wire n_920;
wire n_9200;
wire n_9201;
wire n_9202;
wire n_9203;
wire n_9204;
wire n_9205;
wire n_9206;
wire n_9207;
wire n_9208;
wire n_9209;
wire n_921;
wire n_9210;
wire n_9214;
wire n_9215;
wire n_9216;
wire n_9218;
wire n_9219;
wire n_922;
wire n_9220;
wire n_9221;
wire TIMEBOOST_net_13749;
wire n_9223;
wire n_9224;
wire TIMEBOOST_net_13750;
wire n_9226;
wire n_9227;
wire n_9228;
wire n_9229;
wire n_923;
wire n_9230;
wire n_9231;
wire n_9232;
wire n_9233;
wire n_9234;
wire n_9235;
wire n_9236;
wire n_9237;
wire n_9238;
wire n_9239;
wire n_924;
wire n_9241;
wire n_925;
wire n_9256;
wire n_926;
wire n_9260;
wire n_9261;
wire n_9262;
wire n_9265;
wire n_9269;
wire n_927;
wire n_9270;
wire n_9271;
wire n_9272;
wire n_9274;
wire n_9276;
wire n_9277;
wire n_928;
wire n_9280;
wire n_9283;
wire n_9284;
wire n_9285;
wire n_9286;
wire n_9287;
wire n_929;
wire n_9290;
wire n_9293;
wire n_9294;
wire n_9295;
wire n_9296;
wire n_9297;
wire n_9298;
wire n_9299;
wire n_930;
wire n_9301;
wire n_9303;
wire n_9305;
wire n_9306;
wire n_9307;
wire n_9309;
wire n_931;
wire n_9311;
wire n_9312;
wire n_9315;
wire n_9319;
wire n_9320;
wire n_9321;
wire n_9322;
wire n_9325;
wire n_9328;
wire n_9329;
wire n_9330;
wire n_9331;
wire n_9332;
wire n_9334;
wire n_9335;
wire n_9336;
wire n_9338;
wire n_9340;
wire n_9341;
wire n_9342;
wire n_9343;
wire n_9348;
wire n_9350;
wire n_9353;
wire n_9355;
wire n_9358;
wire n_9361;
wire n_9363;
wire n_9366;
wire n_9368;
wire n_937;
wire n_9371;
wire n_9372;
wire n_9374;
wire n_9377;
wire n_9379;
wire n_938;
wire n_9381;
wire n_9383;
wire n_9385;
wire n_9387;
wire n_9389;
wire n_939;
wire n_9391;
wire n_9393;
wire n_9396;
wire n_9398;
wire n_940;
wire n_9400;
wire n_9402;
wire TIMEBOOST_net_23554;
wire n_9405;
wire TIMEBOOST_net_22274;
wire n_9407;
wire n_9408;
wire n_941;
wire n_9411;
wire n_9412;
wire n_9413;
wire n_9414;
wire n_9418;
wire n_9419;
wire n_9423;
wire TIMEBOOST_net_21170;
wire n_9426;
wire n_9427;
wire n_9428;
wire n_943;
wire n_9430;
wire n_9431;
wire n_9432;
wire n_9433;
wire TIMEBOOST_net_21996;
wire n_9435;
wire n_9436;
wire n_9437;
wire n_9439;
wire n_944;
wire n_9440;
wire n_9441;
wire n_9443;
wire n_9444;
wire n_9448;
wire TIMEBOOST_net_20180;
wire n_945;
wire n_9450;
wire n_9452;
wire n_9454;
wire n_9455;
wire n_9456;
wire TIMEBOOST_net_7320;
wire TIMEBOOST_net_21992;
wire n_9459;
wire n_946;
wire n_9460;
wire TIMEBOOST_net_23403;
wire n_9462;
wire n_9463;
wire TIMEBOOST_net_13297;
wire n_9466;
wire n_9467;
wire TIMEBOOST_net_23399;
wire n_9469;
wire n_947;
wire n_9472;
wire n_9473;
wire n_9474;
wire n_9475;
wire n_9477;
wire n_9478;
wire n_948;
wire n_9480;
wire n_9481;
wire TIMEBOOST_net_12951;
wire TIMEBOOST_net_21983;
wire n_9484;
wire n_9485;
wire n_9486;
wire n_9487;
wire n_9488;
wire n_9490;
wire n_9491;
wire n_9493;
wire n_9494;
wire n_9498;
wire n_9499;
wire n_95;
wire n_950;
wire n_9500;
wire n_9501;
wire n_9502;
wire TIMEBOOST_net_21063;
wire TIMEBOOST_net_13875;
wire n_9506;
wire g65856_db;
wire TIMEBOOST_net_21995;
wire n_9509;
wire n_951;
wire n_9510;
wire TIMEBOOST_net_14058;
wire TIMEBOOST_net_13891;
wire n_9513;
wire TIMEBOOST_net_13889;
wire TIMEBOOST_net_13890;
wire n_9516;
wire n_9517;
wire n_9518;
wire n_9519;
wire n_952;
wire TIMEBOOST_net_23392;
wire n_9524;
wire n_9525;
wire TIMEBOOST_net_13874;
wire n_9528;
wire n_9529;
wire TIMEBOOST_net_17361;
wire n_9531;
wire TIMEBOOST_net_10819;
wire n_9534;
wire TIMEBOOST_net_23234;
wire TIMEBOOST_net_23470;
wire n_9539;
wire n_9542;
wire TIMEBOOST_net_13115;
wire n_9544;
wire TIMEBOOST_net_20523;
wire n_9546;
wire n_9547;
wire n_9548;
wire n_9550;
wire TIMEBOOST_net_21860;
wire n_9554;
wire n_9556;
wire n_9557;
wire TIMEBOOST_net_16048;
wire n_956;
wire n_9561;
wire TIMEBOOST_net_13095;
wire n_9563;
wire TIMEBOOST_net_23198;
wire n_9565;
wire n_9569;
wire n_957;
wire TIMEBOOST_net_14612;
wire n_9572;
wire n_9573;
wire n_9575;
wire n_9576;
wire TIMEBOOST_net_14559;
wire TIMEBOOST_net_12543;
wire TIMEBOOST_net_17446;
wire n_9582;
wire n_9583;
wire n_9584;
wire n_9585;
wire n_9586;
wire n_9588;
wire n_9589;
wire n_959;
wire n_9590;
wire n_9591;
wire n_9593;
wire TIMEBOOST_net_21157;
wire TIMEBOOST_net_21587;
wire n_9598;
wire n_960;
wire n_9604;
wire TIMEBOOST_net_15678;
wire TIMEBOOST_net_13120;
wire TIMEBOOST_net_13387;
wire n_961;
wire TIMEBOOST_net_13385;
wire n_9612;
wire n_9613;
wire n_9615;
wire n_9617;
wire n_9619;
wire TIMEBOOST_net_22157;
wire n_9623;
wire TIMEBOOST_net_12427;
wire TIMEBOOST_net_13431;
wire n_9626;
wire TIMEBOOST_net_21146;
wire TIMEBOOST_net_13119;
wire n_963;
wire n_9631;
wire TIMEBOOST_net_13121;
wire TIMEBOOST_net_22673;
wire n_9637;
wire n_964;
wire n_9642;
wire TIMEBOOST_net_13381;
wire n_9647;
wire n_9648;
wire n_9649;
wire n_965;
wire n_9651;
wire n_9653;
wire n_9655;
wire TIMEBOOST_net_13114;
wire n_9658;
wire n_9659;
wire TIMEBOOST_net_20526;
wire TIMEBOOST_net_7039;
wire n_9663;
wire n_9667;
wire n_9670;
wire n_9671;
wire TIMEBOOST_net_12443;
wire n_9674;
wire n_3676;
wire TIMEBOOST_net_23496;
wire n_9680;
wire n_9682;
wire n_9683;
wire n_9684;
wire n_9685;
wire n_9686;
wire n_9687;
wire TIMEBOOST_net_13116;
wire n_969;
wire n_9690;
wire n_9692;
wire n_9693;
wire n_9694;
wire n_9696;
wire n_9697;
wire n_9700;
wire n_9701;
wire n_9702;
wire n_9705;
wire n_9706;
wire n_9707;
wire n_9708;
wire n_9709;
wire n_971;
wire n_9710;
wire n_9711;
wire n_9712;
wire n_9713;
wire n_9714;
wire n_9716;
wire n_9717;
wire n_9718;
wire n_9719;
wire TIMEBOOST_net_21149;
wire n_9725;
wire n_9726;
wire TIMEBOOST_net_12417;
wire TIMEBOOST_net_20879;
wire n_9729;
wire n_973;
wire n_9732;
wire n_9733;
wire n_9737;
wire n_4232;
wire n_9741;
wire TIMEBOOST_net_23488;
wire n_9744;
wire n_9745;
wire TIMEBOOST_net_21163;
wire n_9747;
wire n_9748;
wire n_9750;
wire n_9751;
wire n_9752;
wire g52400_db;
wire n_9756;
wire TIMEBOOST_net_15555;
wire TIMEBOOST_net_21150;
wire n_976;
wire n_9761;
wire n_9763;
wire TIMEBOOST_net_16359;
wire n_9767;
wire TIMEBOOST_net_12442;
wire n_977;
wire n_9770;
wire TIMEBOOST_net_14887;
wire TIMEBOOST_net_21402;
wire n_9776;
wire n_9777;
wire n_9779;
wire n_978;
wire n_9781;
wire n_9783;
wire TIMEBOOST_net_21265;
wire n_9786;
wire TIMEBOOST_net_12548;
wire n_9788;
wire n_9789;
wire n_9793;
wire TIMEBOOST_net_13108;
wire n_9796;
wire n_9798;
wire n_980;
wire TIMEBOOST_net_13110;
wire n_9802;
wire n_9804;
wire TIMEBOOST_net_12470;
wire n_9807;
wire TIMEBOOST_net_13423;
wire TIMEBOOST_net_14747;
wire TIMEBOOST_net_12469;
wire TIMEBOOST_net_21403;
wire n_9814;
wire n_9816;
wire n_9818;
wire n_982;
wire n_9820;
wire n_9823;
wire TIMEBOOST_net_21484;
wire n_9825;
wire n_9826;
wire TIMEBOOST_net_21184;
wire n_9828;
wire n_983;
wire n_9830;
wire n_9831;
wire n_9832;
wire TIMEBOOST_net_13093;
wire n_9834;
wire TIMEBOOST_net_13094;
wire n_9836;
wire n_9837;
wire TIMEBOOST_net_13091;
wire n_9839;
wire TIMEBOOST_net_17354;
wire n_9841;
wire n_9842;
wire n_9843;
wire n_9844;
wire n_9846;
wire n_9847;
wire TIMEBOOST_net_23547;
wire n_9849;
wire n_9850;
wire n_9851;
wire TIMEBOOST_net_21268;
wire n_9853;
wire n_9854;
wire n_9855;
wire n_9856;
wire n_9857;
wire n_9858;
wire n_9859;
wire n_9860;
wire n_9861;
wire n_9862;
wire TIMEBOOST_net_23481;
wire n_9864;
wire n_9865;
wire n_9867;
wire n_9868;
wire n_9869;
wire n_987;
wire n_9872;
wire n_9874;
wire TIMEBOOST_net_14917;
wire n_9876;
wire TIMEBOOST_net_13109;
wire n_9878;
wire n_9879;
wire n_988;
wire n_9880;
wire n_9881;
wire n_9882;
wire n_9883;
wire n_9884;
wire TIMEBOOST_net_10600;
wire n_9886;
wire n_9887;
wire n_9888;
wire n_9889;
wire n_9890;
wire n_9891;
wire n_9894;
wire n_9895;
wire TIMEBOOST_net_23190;
wire n_9897;
wire n_9898;
wire n_9899;
wire n_990;
wire n_9901;
wire n_9902;
wire TIMEBOOST_net_13429;
wire n_9904;
wire n_9906;
wire n_9908;
wire n_9910;
wire n_9912;
wire n_9914;
wire n_9916;
wire n_9918;
wire n_992;
wire n_9920;
wire n_9922;
wire n_9924;
wire n_9926;
wire n_9928;
wire n_993;
wire n_9931;
wire n_9932;
wire n_994;
wire n_9941;
wire n_9942;
wire n_9947;
wire n_9950;
wire n_9953;
wire n_9956;
wire n_996;
wire n_9962;
wire n_9968;
wire n_9971;
wire n_9975;
wire n_9976;
wire n_9979;
wire n_998;
wire n_9982;
wire n_9988;
wire n_999;
wire n_9991;
wire n_9992;
wire n_9993;
wire n_9997;
wire out_bckp_irdy_out;
wire out_bckp_perr_en_out;
wire output_backup_devsel_out_reg_Q;
wire output_backup_par_en_out_reg_Q;
wire output_backup_par_out_reg_Q;
wire output_backup_perr_out_reg_Q;
wire output_backup_serr_en_out_reg_Q;
wire output_backup_stop_out_reg_Q;
wire output_backup_tar_ad_en_out_reg_Q;
wire output_backup_trdy_out_reg_Q;
wire parchk_pci_ad_out_in;
wire parchk_pci_ad_out_in_1168;
wire parchk_pci_ad_out_in_1169;
wire parchk_pci_ad_out_in_1170;
wire parchk_pci_ad_out_in_1171;
wire parchk_pci_ad_out_in_1172;
wire parchk_pci_ad_out_in_1173;
wire parchk_pci_ad_out_in_1174;
wire parchk_pci_ad_out_in_1175;
wire parchk_pci_ad_out_in_1176;
wire parchk_pci_ad_out_in_1177;
wire parchk_pci_ad_out_in_1178;
wire parchk_pci_ad_out_in_1179;
wire parchk_pci_ad_out_in_1180;
wire parchk_pci_ad_out_in_1181;
wire parchk_pci_ad_out_in_1182;
wire parchk_pci_ad_out_in_1183;
wire parchk_pci_ad_out_in_1184;
wire parchk_pci_ad_out_in_1185;
wire parchk_pci_ad_out_in_1186;
wire parchk_pci_ad_out_in_1187;
wire parchk_pci_ad_out_in_1188;
wire parchk_pci_ad_out_in_1189;
wire parchk_pci_ad_out_in_1190;
wire parchk_pci_ad_out_in_1191;
wire parchk_pci_ad_out_in_1192;
wire parchk_pci_ad_out_in_1193;
wire parchk_pci_ad_out_in_1194;
wire parchk_pci_ad_out_in_1195;
wire parchk_pci_ad_out_in_1196;
wire parchk_pci_ad_out_in_1197;
wire parchk_pci_ad_out_in_1198;
wire parchk_pci_ad_reg_in;
wire parchk_pci_ad_reg_in_1205;
wire parchk_pci_ad_reg_in_1206;
wire parchk_pci_ad_reg_in_1207;
wire parchk_pci_ad_reg_in_1208;
wire parchk_pci_ad_reg_in_1209;
wire parchk_pci_ad_reg_in_1210;
wire parchk_pci_ad_reg_in_1211;
wire parchk_pci_ad_reg_in_1212;
wire parchk_pci_ad_reg_in_1213;
wire parchk_pci_ad_reg_in_1214;
wire parchk_pci_ad_reg_in_1215;
wire parchk_pci_ad_reg_in_1216;
wire parchk_pci_ad_reg_in_1217;
wire parchk_pci_ad_reg_in_1218;
wire parchk_pci_ad_reg_in_1219;
wire parchk_pci_ad_reg_in_1220;
wire parchk_pci_ad_reg_in_1221;
wire parchk_pci_ad_reg_in_1222;
wire parchk_pci_ad_reg_in_1223;
wire parchk_pci_ad_reg_in_1224;
wire parchk_pci_ad_reg_in_1225;
wire parchk_pci_ad_reg_in_1226;
wire parchk_pci_ad_reg_in_1227;
wire parchk_pci_ad_reg_in_1228;
wire parchk_pci_ad_reg_in_1229;
wire parchk_pci_ad_reg_in_1230;
wire parchk_pci_ad_reg_in_1231;
wire parchk_pci_ad_reg_in_1232;
wire parchk_pci_ad_reg_in_1233;
wire parchk_pci_ad_reg_in_1235;
wire parchk_pci_cbe_en_in;
wire parchk_pci_cbe_out_in;
wire parchk_pci_cbe_out_in_1202;
wire parchk_pci_cbe_out_in_1203;
wire parchk_pci_cbe_out_in_1204;
wire parchk_pci_cbe_reg_in;
wire parchk_pci_cbe_reg_in_1236;
wire parchk_pci_cbe_reg_in_1237;
wire parchk_pci_cbe_reg_in_1238;
wire parchk_pci_frame_en_in;
wire parchk_pci_frame_reg_in;
wire parchk_pci_irdy_en_in;
wire parchk_pci_par_en_in;
wire parchk_pci_perr_out_in;
wire parchk_pci_serr_en_in;
wire parchk_pci_serr_out_in;
wire parchk_pci_trdy_en_in;
wire parchk_pci_trdy_reg_in;
wire parity_checker_check_for_serr_on_second;
wire parity_checker_check_for_serr_on_second_reg_Q;
wire parity_checker_check_perr;
wire parity_checker_check_perr_reg_Q;
wire parity_checker_frame_and_irdy_en_prev;
wire parity_checker_frame_and_irdy_en_prev_prev;
wire parity_checker_frame_dec2;
wire parity_checker_master_perr_report;
wire parity_checker_master_perr_report_reg_Q;
wire parity_checker_pci_perr_en_reg;
wire parity_checker_perr_sampled;
wire pci_inti_conf_int_in;
wire pci_resi_conf_soft_res_in;
wire pci_target_unit_del_sync_addr_in;
wire pci_target_unit_del_sync_addr_in_204;
wire pci_target_unit_del_sync_addr_in_205;
wire pci_target_unit_del_sync_addr_in_206;
wire pci_target_unit_del_sync_addr_in_207;
wire pci_target_unit_del_sync_addr_in_208;
wire pci_target_unit_del_sync_addr_in_209;
wire pci_target_unit_del_sync_addr_in_210;
wire pci_target_unit_del_sync_addr_in_211;
wire pci_target_unit_del_sync_addr_in_212;
wire pci_target_unit_del_sync_addr_in_213;
wire pci_target_unit_del_sync_addr_in_214;
wire pci_target_unit_del_sync_addr_in_215;
wire pci_target_unit_del_sync_addr_in_216;
wire pci_target_unit_del_sync_addr_in_217;
wire pci_target_unit_del_sync_addr_in_218;
wire pci_target_unit_del_sync_addr_in_219;
wire pci_target_unit_del_sync_addr_in_220;
wire pci_target_unit_del_sync_addr_in_221;
wire pci_target_unit_del_sync_addr_in_222;
wire pci_target_unit_del_sync_addr_in_223;
wire pci_target_unit_del_sync_addr_in_224;
wire pci_target_unit_del_sync_addr_in_225;
wire pci_target_unit_del_sync_addr_in_226;
wire pci_target_unit_del_sync_addr_in_227;
wire pci_target_unit_del_sync_addr_in_228;
wire pci_target_unit_del_sync_addr_in_229;
wire pci_target_unit_del_sync_addr_in_230;
wire pci_target_unit_del_sync_addr_in_231;
wire pci_target_unit_del_sync_addr_in_232;
wire pci_target_unit_del_sync_addr_in_233;
wire pci_target_unit_del_sync_addr_in_234;
wire pci_target_unit_del_sync_bc_in;
wire pci_target_unit_del_sync_bc_in_201;
wire pci_target_unit_del_sync_bc_in_202;
wire pci_target_unit_del_sync_bc_in_203;
wire pci_target_unit_del_sync_be_out_reg_0__Q;
wire pci_target_unit_del_sync_be_out_reg_1__Q;
wire pci_target_unit_del_sync_be_out_reg_2__Q;
wire pci_target_unit_del_sync_be_out_reg_3__Q;
wire pci_target_unit_del_sync_comp_cycle_count_0_;
wire pci_target_unit_del_sync_comp_cycle_count_10_;
wire pci_target_unit_del_sync_comp_cycle_count_11_;
wire pci_target_unit_del_sync_comp_cycle_count_12_;
wire pci_target_unit_del_sync_comp_cycle_count_13_;
wire pci_target_unit_del_sync_comp_cycle_count_14_;
wire pci_target_unit_del_sync_comp_cycle_count_15_;
wire pci_target_unit_del_sync_comp_cycle_count_1_;
wire pci_target_unit_del_sync_comp_cycle_count_2_;
wire pci_target_unit_del_sync_comp_cycle_count_3_;
wire pci_target_unit_del_sync_comp_cycle_count_4_;
wire pci_target_unit_del_sync_comp_cycle_count_5_;
wire pci_target_unit_del_sync_comp_cycle_count_6_;
wire pci_target_unit_del_sync_comp_cycle_count_7_;
wire pci_target_unit_del_sync_comp_cycle_count_8_;
wire pci_target_unit_del_sync_comp_cycle_count_9_;
wire pci_target_unit_del_sync_comp_cycle_count_reg_16__Q;
wire pci_target_unit_del_sync_comp_done_reg_clr;
wire pci_target_unit_del_sync_comp_done_reg_clr_reg_Q;
wire pci_target_unit_del_sync_comp_done_reg_main;
wire pci_target_unit_del_sync_comp_done_reg_main_reg_Q;
wire pci_target_unit_del_sync_comp_flush_out_reg_Q;
wire pci_target_unit_del_sync_comp_in;
wire pci_target_unit_del_sync_comp_rty_exp_clr;
wire pci_target_unit_del_sync_comp_rty_exp_clr_reg_Q;
wire pci_target_unit_del_sync_comp_rty_exp_reg;
wire pci_target_unit_del_sync_req_comp_pending;
wire pci_target_unit_del_sync_req_comp_pending_sample;
wire pci_target_unit_del_sync_req_comp_pending_sample_reg_Q;
wire pci_target_unit_del_sync_req_done_reg;
wire pci_target_unit_del_sync_req_rty_exp_clr;
wire pci_target_unit_del_sync_req_rty_exp_clr_reg_Q;
wire pci_target_unit_del_sync_req_rty_exp_reg;
wire pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__Q;
wire pci_target_unit_del_sync_sync_comp_done;
wire pci_target_unit_del_sync_sync_comp_req_pending;
wire pci_target_unit_del_sync_sync_comp_rty_exp_clr;
wire pci_target_unit_del_sync_sync_req_comp_pending;
wire pci_target_unit_del_sync_sync_req_rty_exp;
wire pci_target_unit_fifos_inGreyCount_0_;
wire pci_target_unit_fifos_inGreyCount_reg_0__Q;
wire pci_target_unit_fifos_inGreyCount_reg_1__Q;
wire pci_target_unit_fifos_outGreyCount_0_;
wire pci_target_unit_fifos_outGreyCount_reg_0__Q;
wire pci_target_unit_fifos_outGreyCount_reg_1__Q;
wire pci_target_unit_fifos_pcir_control_in_192;
wire pci_target_unit_fifos_pcir_data_in;
wire pci_target_unit_fifos_pcir_data_in_158;
wire pci_target_unit_fifos_pcir_data_in_159;
wire pci_target_unit_fifos_pcir_data_in_160;
wire pci_target_unit_fifos_pcir_data_in_161;
wire pci_target_unit_fifos_pcir_data_in_162;
wire pci_target_unit_fifos_pcir_data_in_163;
wire pci_target_unit_fifos_pcir_data_in_164;
wire pci_target_unit_fifos_pcir_data_in_165;
wire pci_target_unit_fifos_pcir_data_in_166;
wire pci_target_unit_fifos_pcir_data_in_167;
wire pci_target_unit_fifos_pcir_data_in_168;
wire pci_target_unit_fifos_pcir_data_in_169;
wire pci_target_unit_fifos_pcir_data_in_170;
wire pci_target_unit_fifos_pcir_data_in_171;
wire pci_target_unit_fifos_pcir_data_in_172;
wire pci_target_unit_fifos_pcir_data_in_173;
wire pci_target_unit_fifos_pcir_data_in_174;
wire pci_target_unit_fifos_pcir_data_in_175;
wire pci_target_unit_fifos_pcir_data_in_176;
wire pci_target_unit_fifos_pcir_data_in_177;
wire pci_target_unit_fifos_pcir_data_in_178;
wire pci_target_unit_fifos_pcir_data_in_179;
wire pci_target_unit_fifos_pcir_data_in_180;
wire pci_target_unit_fifos_pcir_data_in_181;
wire pci_target_unit_fifos_pcir_data_in_182;
wire pci_target_unit_fifos_pcir_data_in_183;
wire pci_target_unit_fifos_pcir_data_in_184;
wire pci_target_unit_fifos_pcir_data_in_185;
wire pci_target_unit_fifos_pcir_data_in_186;
wire pci_target_unit_fifos_pcir_data_in_187;
wire pci_target_unit_fifos_pcir_data_in_188;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_39;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_40;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_100;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_101;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_;
wire pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q;
wire pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q;
wire pci_target_unit_fifos_pcir_flush_in;
wire pci_target_unit_fifos_pcir_wenable_in;
wire pci_target_unit_fifos_pcir_whole_waddr;
wire pci_target_unit_fifos_pcir_whole_waddr_94;
wire pci_target_unit_fifos_pciw_addr_data_in;
wire pci_target_unit_fifos_pciw_addr_data_in_121;
wire pci_target_unit_fifos_pciw_addr_data_in_122;
wire pci_target_unit_fifos_pciw_addr_data_in_123;
wire pci_target_unit_fifos_pciw_addr_data_in_124;
wire pci_target_unit_fifos_pciw_addr_data_in_125;
wire pci_target_unit_fifos_pciw_addr_data_in_126;
wire pci_target_unit_fifos_pciw_addr_data_in_127;
wire pci_target_unit_fifos_pciw_addr_data_in_128;
wire pci_target_unit_fifos_pciw_addr_data_in_129;
wire pci_target_unit_fifos_pciw_addr_data_in_130;
wire pci_target_unit_fifos_pciw_addr_data_in_131;
wire pci_target_unit_fifos_pciw_addr_data_in_132;
wire pci_target_unit_fifos_pciw_addr_data_in_133;
wire pci_target_unit_fifos_pciw_addr_data_in_134;
wire pci_target_unit_fifos_pciw_addr_data_in_135;
wire pci_target_unit_fifos_pciw_addr_data_in_136;
wire pci_target_unit_fifos_pciw_addr_data_in_137;
wire pci_target_unit_fifos_pciw_addr_data_in_138;
wire pci_target_unit_fifos_pciw_addr_data_in_139;
wire pci_target_unit_fifos_pciw_addr_data_in_140;
wire pci_target_unit_fifos_pciw_addr_data_in_141;
wire pci_target_unit_fifos_pciw_addr_data_in_142;
wire pci_target_unit_fifos_pciw_addr_data_in_143;
wire pci_target_unit_fifos_pciw_addr_data_in_144;
wire pci_target_unit_fifos_pciw_addr_data_in_145;
wire pci_target_unit_fifos_pciw_addr_data_in_146;
wire pci_target_unit_fifos_pciw_addr_data_in_147;
wire pci_target_unit_fifos_pciw_addr_data_in_148;
wire pci_target_unit_fifos_pciw_addr_data_in_149;
wire pci_target_unit_fifos_pciw_addr_data_in_150;
wire pci_target_unit_fifos_pciw_addr_data_in_151;
wire pci_target_unit_fifos_pciw_cbe_in;
wire pci_target_unit_fifos_pciw_cbe_in_152;
wire pci_target_unit_fifos_pciw_cbe_in_153;
wire pci_target_unit_fifos_pciw_cbe_in_154;
wire pci_target_unit_fifos_pciw_control_in;
wire pci_target_unit_fifos_pciw_control_in_155;
wire pci_target_unit_fifos_pciw_control_in_156;
wire pci_target_unit_fifos_pciw_control_in_157;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_74;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_75;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q;
wire pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus2;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_94;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_95;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_;
wire pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_;
wire pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_0__153;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_1__192;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_2__231;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_3__270;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q;
wire pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q;
wire pci_target_unit_fifos_pciw_inTransactionCount_0_;
wire pci_target_unit_fifos_pciw_inTransactionCount_1_;
wire pci_target_unit_fifos_pciw_inTransactionCount_reg_1__Q;
wire pci_target_unit_fifos_pciw_outTransactionCount_1_;
wire pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q;
wire pci_target_unit_fifos_pciw_outTransactionCount_reg_1__Q;
wire pci_target_unit_fifos_pciw_wenable_in;
wire pci_target_unit_fifos_pciw_whole_waddr;
wire pci_target_unit_fifos_pciw_whole_waddr_47;
wire pci_target_unit_fifos_wb_clk_inGreyCount_0_;
wire pci_target_unit_fifos_wb_clk_inGreyCount_1_;
wire pci_target_unit_fifos_wb_clk_sync_inGreyCount;
wire pci_target_unit_fifos_wb_clk_sync_inGreyCount_36;
wire pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_Q;
wire pci_target_unit_pci_target_if_keep_desconnect_wo_data_set;
wire pci_target_unit_pci_target_if_norm_address_reg_0__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_1__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_2__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_3__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_4__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_5__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_6__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_7__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_8__Q;
wire pci_target_unit_pci_target_if_norm_address_reg_9__Q;
wire pci_target_unit_pci_target_if_norm_prf_en;
wire pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q;
wire pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q;
wire pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__Q;
wire pci_target_unit_pci_target_if_same_read_reg;
wire pci_target_unit_pci_target_if_target_rd_completed;
wire pci_target_unit_pci_target_sm_backoff;
wire pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_Q;
wire pci_target_unit_pci_target_sm_cnf_progress;
wire pci_target_unit_pci_target_sm_master_will_request_read;
wire pci_target_unit_pci_target_sm_n_2;
wire pci_target_unit_pci_target_sm_n_3;
wire pci_target_unit_pci_target_sm_previous_frame;
wire pci_target_unit_pci_target_sm_rd_from_fifo;
wire pci_target_unit_pci_target_sm_rd_progress;
wire pci_target_unit_pci_target_sm_rd_request;
wire pci_target_unit_pci_target_sm_rd_request_reg_Q;
wire pci_target_unit_pci_target_sm_read_completed_reg;
wire pci_target_unit_pci_target_sm_read_completed_reg_reg_Q;
wire pci_target_unit_pci_target_sm_same_read_reg;
wire pci_target_unit_pci_target_sm_state_backoff_reg_reg_Q;
wire pci_target_unit_pci_target_sm_state_transfere_reg;
wire pci_target_unit_pci_target_sm_state_transfere_reg_reg_Q;
wire pci_target_unit_pci_target_sm_wr_progress;
wire pci_target_unit_pci_target_sm_wr_to_fifo;
wire pci_target_unit_pcit_if_comp_flush_in;
wire pci_target_unit_pcit_if_pcir_fifo_control_in_637;
wire pci_target_unit_pcit_if_pcir_fifo_data_in;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_766;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_767;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_768;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_769;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_770;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_771;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_772;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_773;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_774;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_775;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_776;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_777;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_778;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_779;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_780;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_781;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_782;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_783;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_784;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_785;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_786;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_787;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_788;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_789;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_790;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_791;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_792;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_793;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_794;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_795;
wire pci_target_unit_pcit_if_pcir_fifo_data_in_796;
wire pci_target_unit_pcit_if_req_req_pending_in;
wire pci_target_unit_pcit_if_strd_addr_in;
wire pci_target_unit_pcit_if_strd_addr_in_686;
wire pci_target_unit_pcit_if_strd_addr_in_687;
wire pci_target_unit_pcit_if_strd_addr_in_688;
wire pci_target_unit_pcit_if_strd_addr_in_689;
wire pci_target_unit_pcit_if_strd_addr_in_690;
wire pci_target_unit_pcit_if_strd_addr_in_691;
wire pci_target_unit_pcit_if_strd_addr_in_692;
wire pci_target_unit_pcit_if_strd_addr_in_693;
wire pci_target_unit_pcit_if_strd_addr_in_694;
wire pci_target_unit_pcit_if_strd_addr_in_695;
wire pci_target_unit_pcit_if_strd_addr_in_696;
wire pci_target_unit_pcit_if_strd_addr_in_697;
wire pci_target_unit_pcit_if_strd_addr_in_698;
wire pci_target_unit_pcit_if_strd_addr_in_699;
wire pci_target_unit_pcit_if_strd_addr_in_700;
wire pci_target_unit_pcit_if_strd_addr_in_701;
wire pci_target_unit_pcit_if_strd_addr_in_702;
wire pci_target_unit_pcit_if_strd_addr_in_703;
wire pci_target_unit_pcit_if_strd_addr_in_704;
wire pci_target_unit_pcit_if_strd_addr_in_705;
wire pci_target_unit_pcit_if_strd_addr_in_706;
wire pci_target_unit_pcit_if_strd_addr_in_707;
wire pci_target_unit_pcit_if_strd_addr_in_708;
wire pci_target_unit_pcit_if_strd_addr_in_709;
wire pci_target_unit_pcit_if_strd_addr_in_710;
wire pci_target_unit_pcit_if_strd_addr_in_711;
wire pci_target_unit_pcit_if_strd_addr_in_712;
wire pci_target_unit_pcit_if_strd_addr_in_713;
wire pci_target_unit_pcit_if_strd_addr_in_714;
wire pci_target_unit_pcit_if_strd_addr_in_715;
wire pci_target_unit_pcit_if_strd_addr_in_716;
wire pci_target_unit_pcit_if_strd_bc_in;
wire pci_target_unit_pcit_if_strd_bc_in_717;
wire pci_target_unit_pcit_if_strd_bc_in_718;
wire pci_target_unit_pcit_if_strd_bc_in_719;
wire pci_target_unit_wbm_sm_pci_tar_burst_ok;
wire pci_target_unit_wbm_sm_pci_tar_read_request;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79;
wire pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80;
wire pci_target_unit_wbm_sm_pciw_fifo_cbe_in;
wire pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81;
wire pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82;
wire pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83;
wire pci_target_unit_wbm_sm_pciw_fifo_control_in;
wire pci_target_unit_wbm_sm_pciw_fifo_control_in_84;
wire pci_target_unit_wbm_sm_pciw_fifo_control_in_85;
wire pci_target_unit_wbm_sm_pciw_fifo_control_in_86;
wire pci_target_unit_wishbone_master_addr_into_cnt_reg;
wire pci_target_unit_wishbone_master_bc_register_reg_0__Q;
wire pci_target_unit_wishbone_master_bc_register_reg_1__Q;
wire pci_target_unit_wishbone_master_bc_register_reg_2__Q;
wire pci_target_unit_wishbone_master_bc_register_reg_3__Q;
wire pci_target_unit_wishbone_master_burst_chopped;
wire pci_target_unit_wishbone_master_burst_chopped_delayed;
wire pci_target_unit_wishbone_master_burst_chopped_delayed_reg_Q;
wire pci_target_unit_wishbone_master_c_state_0_;
wire pci_target_unit_wishbone_master_c_state_1_;
wire pci_target_unit_wishbone_master_c_state_2_;
wire pci_target_unit_wishbone_master_first_data_is_burst_reg;
wire pci_target_unit_wishbone_master_first_wb_data_access;
wire pci_target_unit_wishbone_master_read_bound;
wire pci_target_unit_wishbone_master_read_count_0_;
wire pci_target_unit_wishbone_master_read_count_1_;
wire pci_target_unit_wishbone_master_read_count_reg_2__Q;
wire pci_target_unit_wishbone_master_reset_rty_cnt;
wire pci_target_unit_wishbone_master_reset_rty_cnt_reg_Q;
wire pci_target_unit_wishbone_master_retried;
wire pci_target_unit_wishbone_master_rty_counter_0_;
wire pci_target_unit_wishbone_master_rty_counter_1_;
wire pci_target_unit_wishbone_master_rty_counter_3_;
wire pci_target_unit_wishbone_master_rty_counter_4_;
wire pci_target_unit_wishbone_master_rty_counter_5_;
wire pci_target_unit_wishbone_master_rty_counter_6_;
wire pci_target_unit_wishbone_master_rty_counter_7_;
wire pci_target_unit_wishbone_master_wb_cyc_o_reg_Q;
wire pciu_am1_in;
wire pciu_am1_in_518;
wire pciu_am1_in_519;
wire pciu_am1_in_520;
wire pciu_am1_in_521;
wire pciu_am1_in_522;
wire pciu_am1_in_523;
wire pciu_am1_in_524;
wire pciu_am1_in_525;
wire pciu_am1_in_526;
wire pciu_am1_in_527;
wire pciu_am1_in_528;
wire pciu_am1_in_529;
wire pciu_am1_in_530;
wire pciu_am1_in_531;
wire pciu_am1_in_532;
wire pciu_am1_in_533;
wire pciu_am1_in_534;
wire pciu_am1_in_535;
wire pciu_am1_in_536;
wire pciu_am1_in_537;
wire pciu_am1_in_538;
wire pciu_am1_in_539;
wire pciu_am1_in_540;
wire pciu_bar0_in;
wire pciu_bar0_in_361;
wire pciu_bar0_in_362;
wire pciu_bar0_in_363;
wire pciu_bar0_in_364;
wire pciu_bar0_in_365;
wire pciu_bar0_in_366;
wire pciu_bar0_in_367;
wire pciu_bar0_in_368;
wire pciu_bar0_in_369;
wire pciu_bar0_in_370;
wire pciu_bar0_in_371;
wire pciu_bar0_in_372;
wire pciu_bar0_in_373;
wire pciu_bar0_in_374;
wire pciu_bar0_in_375;
wire pciu_bar0_in_376;
wire pciu_bar0_in_377;
wire pciu_bar0_in_378;
wire pciu_bar0_in_379;
wire pciu_bar1_in;
wire pciu_bar1_in_380;
wire pciu_bar1_in_381;
wire pciu_bar1_in_382;
wire pciu_bar1_in_383;
wire pciu_bar1_in_384;
wire pciu_bar1_in_385;
wire pciu_bar1_in_386;
wire pciu_bar1_in_387;
wire pciu_bar1_in_388;
wire pciu_bar1_in_389;
wire pciu_bar1_in_390;
wire pciu_bar1_in_391;
wire pciu_bar1_in_392;
wire pciu_bar1_in_393;
wire pciu_bar1_in_394;
wire pciu_bar1_in_395;
wire pciu_bar1_in_396;
wire pciu_bar1_in_397;
wire pciu_bar1_in_398;
wire pciu_bar1_in_399;
wire pciu_bar1_in_400;
wire pciu_bar1_in_401;
wire pciu_bar1_in_402;
wire pciu_cache_line_size_in_775;
wire pciu_cache_line_size_in_776;
wire pciu_cache_line_size_in_777;
wire pciu_cache_lsize_not_zero_in;
wire pciu_pciif_bckp_stop_in;
wire pciu_pciif_idsel_reg_in;
wire pciu_pciif_stop_reg_in;
wire pciu_pref_en_in_320;
wire wbm_cyc_o_1378;
wire wbs_ack_o_1307;
wire wbs_err_o_1309;
wire wbs_rty_o_1308;
wire wbs_wbb3_2_wbb2_dat_o_i;
wire wbs_wbb3_2_wbb2_dat_o_i_100;
wire wbs_wbb3_2_wbb2_dat_o_i_101;
wire wbs_wbb3_2_wbb2_dat_o_i_102;
wire wbs_wbb3_2_wbb2_dat_o_i_103;
wire wbs_wbb3_2_wbb2_dat_o_i_104;
wire wbs_wbb3_2_wbb2_dat_o_i_105;
wire wbs_wbb3_2_wbb2_dat_o_i_106;
wire wbs_wbb3_2_wbb2_dat_o_i_107;
wire wbs_wbb3_2_wbb2_dat_o_i_108;
wire wbs_wbb3_2_wbb2_dat_o_i_109;
wire wbs_wbb3_2_wbb2_dat_o_i_110;
wire wbs_wbb3_2_wbb2_dat_o_i_111;
wire wbs_wbb3_2_wbb2_dat_o_i_112;
wire wbs_wbb3_2_wbb2_dat_o_i_113;
wire wbs_wbb3_2_wbb2_dat_o_i_114;
wire wbs_wbb3_2_wbb2_dat_o_i_115;
wire wbs_wbb3_2_wbb2_dat_o_i_116;
wire wbs_wbb3_2_wbb2_dat_o_i_117;
wire wbs_wbb3_2_wbb2_dat_o_i_118;
wire wbs_wbb3_2_wbb2_dat_o_i_119;
wire wbs_wbb3_2_wbb2_dat_o_i_120;
wire wbs_wbb3_2_wbb2_dat_o_i_121;
wire wbs_wbb3_2_wbb2_dat_o_i_122;
wire wbs_wbb3_2_wbb2_dat_o_i_123;
wire wbs_wbb3_2_wbb2_dat_o_i_124;
wire wbs_wbb3_2_wbb2_dat_o_i_125;
wire wbs_wbb3_2_wbb2_dat_o_i_126;
wire wbs_wbb3_2_wbb2_dat_o_i_127;
wire wbs_wbb3_2_wbb2_dat_o_i_128;
wire wbs_wbb3_2_wbb2_dat_o_i_129;
wire wbs_wbb3_2_wbb2_dat_o_i_130;
wire wbu_addr_in;
wire wbu_addr_in_250;
wire wbu_addr_in_251;
wire wbu_addr_in_252;
wire wbu_addr_in_253;
wire wbu_addr_in_254;
wire wbu_addr_in_255;
wire wbu_addr_in_256;
wire wbu_addr_in_257;
wire wbu_addr_in_258;
wire wbu_addr_in_259;
wire wbu_addr_in_260;
wire wbu_addr_in_261;
wire wbu_addr_in_262;
wire wbu_addr_in_263;
wire wbu_addr_in_264;
wire wbu_addr_in_265;
wire wbu_addr_in_266;
wire wbu_addr_in_267;
wire wbu_addr_in_268;
wire wbu_addr_in_269;
wire wbu_addr_in_270;
wire wbu_addr_in_271;
wire wbu_addr_in_272;
wire wbu_addr_in_273;
wire wbu_addr_in_274;
wire wbu_addr_in_275;
wire wbu_addr_in_276;
wire wbu_addr_in_277;
wire wbu_addr_in_278;
wire wbu_addr_in_279;
wire wbu_addr_in_280;
wire wbu_am1_in;
wire wbu_am2_in;
wire wbu_bar1_in;
wire wbu_bar2_in;
wire wbu_cache_line_size_in_206;
wire wbu_cache_line_size_in_207;
wire wbu_cache_line_size_in_208;
wire wbu_cache_line_size_in_209;
wire wbu_cache_line_size_in_210;
wire wbu_cache_line_size_in_211;
wire wbu_latency_tim_val_in;
wire wbu_latency_tim_val_in_243;
wire wbu_latency_tim_val_in_244;
wire wbu_latency_tim_val_in_245;
wire wbu_latency_tim_val_in_246;
wire wbu_latency_tim_val_in_247;
wire wbu_latency_tim_val_in_248;
wire wbu_latency_tim_val_in_249;
wire wbu_map_in_131;
wire wbu_map_in_132;
wire wbu_mrl_en_in_141;
wire wbu_mrl_en_in_142;
wire wbu_pci_drcomp_pending_in;
wire wbu_pciif_devsel_reg_in;
wire wbu_pciif_frame_out_in;
wire wbu_pref_en_in_136;
wire wbu_pref_en_in_137;
wire wbu_sel_in;
wire wbu_sel_in_312;
wire wbu_sel_in_313;
wire wbu_sel_in_314;
wire wbu_wb_init_complete_in;
wire wbu_we_in;
wire wishbone_slave_unit_del_sync_addr_out_reg_0__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_10__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_11__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_12__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_13__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_14__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_15__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_16__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_17__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_18__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_19__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_1__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_20__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_21__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_22__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_23__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_24__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_25__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_26__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_27__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_28__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_29__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_2__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_30__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_31__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_3__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_4__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_5__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_6__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_7__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_8__Q;
wire wishbone_slave_unit_del_sync_addr_out_reg_9__Q;
wire wishbone_slave_unit_del_sync_bc_out_reg_0__Q;
wire wishbone_slave_unit_del_sync_bc_out_reg_1__Q;
wire wishbone_slave_unit_del_sync_bc_out_reg_2__Q;
wire wishbone_slave_unit_del_sync_bc_out_reg_3__Q;
wire wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_0_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_10_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_11_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_12_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_1_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_2_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_3_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_4_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_5_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_6_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_7_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_8_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_9_;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__Q;
wire wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__Q;
wire wishbone_slave_unit_del_sync_comp_done_reg_clr;
wire wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_Q;
wire wishbone_slave_unit_del_sync_comp_done_reg_main;
wire wishbone_slave_unit_del_sync_comp_flush_out;
wire wishbone_slave_unit_del_sync_comp_req_pending_reg_Q;
wire wishbone_slave_unit_del_sync_comp_rty_exp_clr;
wire wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_Q;
wire wishbone_slave_unit_del_sync_comp_rty_exp_reg;
wire wishbone_slave_unit_del_sync_req_comp_pending;
wire wishbone_slave_unit_del_sync_req_comp_pending_sample;
wire wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_Q;
wire wishbone_slave_unit_del_sync_req_done_reg;
wire wishbone_slave_unit_del_sync_req_done_reg_reg_Q;
wire wishbone_slave_unit_del_sync_req_rty_exp_clr;
wire wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_Q;
wire wishbone_slave_unit_del_sync_req_rty_exp_reg;
wire wishbone_slave_unit_del_sync_sync_comp_done;
wire wishbone_slave_unit_del_sync_sync_comp_req_pending;
wire wishbone_slave_unit_del_sync_sync_comp_rty_exp_clr;
wire wishbone_slave_unit_del_sync_sync_req_comp_pending;
wire wishbone_slave_unit_del_sync_sync_req_rty_exp;
wire wishbone_slave_unit_del_sync_we_out_reg_Q;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_100;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_101;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_70;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_71;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_72;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_73;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_74;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_75;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_76;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_77;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_78;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_79;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_80;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_81;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_82;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_83;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_84;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_85;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_86;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_87;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_88;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_89;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_90;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_91;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_92;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_93;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_94;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_95;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_96;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_97;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_98;
wire wishbone_slave_unit_delayed_write_data_comp_wdata_out_99;
wire wishbone_slave_unit_fifos_inGreyCount_0_;
wire wishbone_slave_unit_fifos_inGreyCount_reg_0__Q;
wire wishbone_slave_unit_fifos_inGreyCount_reg_1__Q;
wire wishbone_slave_unit_fifos_inGreyCount_reg_2__Q;
wire wishbone_slave_unit_fifos_outGreyCount_0_;
wire wishbone_slave_unit_fifos_outGreyCount_1_;
wire wishbone_slave_unit_fifos_outGreyCount_2_;
wire wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_;
wire wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_;
wire wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_;
wire wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__Q;
wire wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount;
wire wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_49;
wire wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_50;
wire wishbone_slave_unit_fifos_wbr_be_in;
wire wishbone_slave_unit_fifos_wbr_be_in_264;
wire wishbone_slave_unit_fifos_wbr_be_in_265;
wire wishbone_slave_unit_fifos_wbr_be_in_266;
wire wishbone_slave_unit_fifos_wbr_control_in;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_45;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_46;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_47;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__531;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__248;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__265;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__363;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__365;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__379;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__Q;
wire wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__Q;
wire wishbone_slave_unit_fifos_wbr_whole_waddr;
wire wishbone_slave_unit_fifos_wbr_whole_waddr_104;
wire wishbone_slave_unit_fifos_wbr_whole_waddr_105;
wire wishbone_slave_unit_fifos_wbr_whole_waddr_106;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_70;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_71;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_72;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus1;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_93;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_94;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_95;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_;
wire wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_4__213;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q;
wire wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_0_;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_1_;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__Q;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__Q;
wire wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_0_;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_1_;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__Q;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__Q;
wire wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q;
wire wishbone_slave_unit_fifos_wbw_whole_waddr;
wire wishbone_slave_unit_fifos_wbw_whole_waddr_55;
wire wishbone_slave_unit_fifos_wbw_whole_waddr_56;
wire wishbone_slave_unit_fifos_wbw_whole_waddr_57;
wire wishbone_slave_unit_pci_initiator_if_current_byte_address;
wire wishbone_slave_unit_pci_initiator_if_current_byte_address_36;
wire wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q;
wire wishbone_slave_unit_pci_initiator_if_data_source;
wire wishbone_slave_unit_pci_initiator_if_del_read_req;
wire wishbone_slave_unit_pci_initiator_if_del_write_req;
wire wishbone_slave_unit_pci_initiator_if_err_recovery;
wire wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q;
wire wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q;
wire wishbone_slave_unit_pci_initiator_if_posted_write_req;
wire wishbone_slave_unit_pci_initiator_if_read_bound;
wire wishbone_slave_unit_pci_initiator_if_read_count_0_;
wire wishbone_slave_unit_pci_initiator_if_read_count_1_;
wire wishbone_slave_unit_pci_initiator_if_read_count_2_;
wire wishbone_slave_unit_pci_initiator_if_read_count_3_;
wire wishbone_slave_unit_pci_initiator_if_read_count_reg_3__Q;
wire wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_Q;
wire wishbone_slave_unit_pci_initiator_if_write_req_int;
wire wishbone_slave_unit_pci_initiator_sm_cur_state_0_;
wire wishbone_slave_unit_pci_initiator_sm_cur_state_1_;
wire wishbone_slave_unit_pci_initiator_sm_cur_state_2_;
wire wishbone_slave_unit_pci_initiator_sm_cur_state_3_;
wire wishbone_slave_unit_pci_initiator_sm_decode_count_0_;
wire wishbone_slave_unit_pci_initiator_sm_decode_count_1_;
wire wishbone_slave_unit_pci_initiator_sm_decode_count_2_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_0_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_1_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_2_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_3_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_4_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_5_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_6_;
wire wishbone_slave_unit_pci_initiator_sm_latency_timer_7_;
wire wishbone_slave_unit_pci_initiator_sm_mabort1;
wire wishbone_slave_unit_pci_initiator_sm_mabort2;
wire wishbone_slave_unit_pci_initiator_sm_rdata_selector;
wire wishbone_slave_unit_pci_initiator_sm_rdata_selector_14;
wire wishbone_slave_unit_pci_initiator_sm_timeout;
wire wishbone_slave_unit_pci_initiator_sm_transfer;
wire wishbone_slave_unit_pcim_if_del_bc_in;
wire wishbone_slave_unit_pcim_if_del_bc_in_382;
wire wishbone_slave_unit_pcim_if_del_bc_in_383;
wire wishbone_slave_unit_pcim_if_del_burst_in;
wire wishbone_slave_unit_pcim_if_del_req_in;
wire wishbone_slave_unit_pcim_if_del_we_in;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_384;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_385;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_386;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_387;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_388;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_389;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_390;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_391;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_392;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_393;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_394;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_395;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_396;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_397;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_398;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_399;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_400;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_401;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_402;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_403;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_404;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_405;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_406;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_407;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_408;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_409;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_410;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_411;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_412;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_413;
wire wishbone_slave_unit_pcim_if_wbw_addr_data_in_414;
wire wishbone_slave_unit_pcim_if_wbw_cbe_in;
wire wishbone_slave_unit_pcim_if_wbw_cbe_in_416;
wire wishbone_slave_unit_pcim_if_wbw_cbe_in_417;
wire wishbone_slave_unit_pcim_sm_be_in_557;
wire wishbone_slave_unit_pcim_sm_be_in_558;
wire wishbone_slave_unit_pcim_sm_be_in_559;
wire wishbone_slave_unit_pcim_sm_data_in;
wire wishbone_slave_unit_pcim_sm_data_in_635;
wire wishbone_slave_unit_pcim_sm_data_in_636;
wire wishbone_slave_unit_pcim_sm_data_in_637;
wire wishbone_slave_unit_pcim_sm_data_in_638;
wire wishbone_slave_unit_pcim_sm_data_in_639;
wire wishbone_slave_unit_pcim_sm_data_in_640;
wire wishbone_slave_unit_pcim_sm_data_in_641;
wire wishbone_slave_unit_pcim_sm_data_in_642;
wire wishbone_slave_unit_pcim_sm_data_in_643;
wire wishbone_slave_unit_pcim_sm_data_in_644;
wire wishbone_slave_unit_pcim_sm_data_in_645;
wire wishbone_slave_unit_pcim_sm_data_in_646;
wire wishbone_slave_unit_pcim_sm_data_in_647;
wire wishbone_slave_unit_pcim_sm_data_in_648;
wire wishbone_slave_unit_pcim_sm_data_in_649;
wire wishbone_slave_unit_pcim_sm_data_in_650;
wire wishbone_slave_unit_pcim_sm_data_in_651;
wire wishbone_slave_unit_pcim_sm_data_in_652;
wire wishbone_slave_unit_pcim_sm_data_in_653;
wire wishbone_slave_unit_pcim_sm_data_in_654;
wire wishbone_slave_unit_pcim_sm_data_in_655;
wire wishbone_slave_unit_pcim_sm_data_in_656;
wire wishbone_slave_unit_pcim_sm_data_in_657;
wire wishbone_slave_unit_pcim_sm_data_in_658;
wire wishbone_slave_unit_pcim_sm_data_in_659;
wire wishbone_slave_unit_pcim_sm_data_in_660;
wire wishbone_slave_unit_pcim_sm_data_in_661;
wire wishbone_slave_unit_pcim_sm_data_in_662;
wire wishbone_slave_unit_pcim_sm_data_in_663;
wire wishbone_slave_unit_pcim_sm_data_in_664;
wire wishbone_slave_unit_pcim_sm_data_in_665;
wire wishbone_slave_unit_pcim_sm_last_in;
wire wishbone_slave_unit_pcim_sm_rdy_in;
wire wishbone_slave_unit_wbs_sm_del_req_pending_in;
wire wishbone_slave_unit_wbs_sm_wbr_control_in;
wire wishbone_slave_unit_wbs_sm_wbr_control_in_190;
wire wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_Q;
wire wishbone_slave_unit_wishbone_slave_c_state;
wire wishbone_slave_unit_wishbone_slave_c_state_1;
wire wishbone_slave_unit_wishbone_slave_c_state_2;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q;
wire wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q;
wire wishbone_slave_unit_wishbone_slave_del_addr_hit;
wire wishbone_slave_unit_wishbone_slave_del_completion_allow;
wire wishbone_slave_unit_wishbone_slave_do_del_request;
wire wishbone_slave_unit_wishbone_slave_img_hit_0_;
wire wishbone_slave_unit_wishbone_slave_img_hit_1_;
wire wishbone_slave_unit_wishbone_slave_img_hit_2_;
wire wishbone_slave_unit_wishbone_slave_img_hit_3_;
wire wishbone_slave_unit_wishbone_slave_img_hit_4_;
wire wishbone_slave_unit_wishbone_slave_img_wallow;
wire wishbone_slave_unit_wishbone_slave_map;
wire wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q;
wire wishbone_slave_unit_wishbone_slave_pref_en_reg_Q;
wire wishbone_slave_unit_wishbone_slave_wb_conf_hit;
wire wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_Q;
wire TIMEBOOST_net_0;
wire TIMEBOOST_net_1;
wire TIMEBOOST_net_2;
wire TIMEBOOST_net_3;
wire TIMEBOOST_net_4;
wire TIMEBOOST_net_5;

// Start cells
in01f08 FE_OCPC1822_n_16560 ( .a(n_16560), .o(FE_OCPN1822_n_16560) );
in01f10 FE_OCPC1823_n_16560 ( .a(FE_OCPN1822_n_16560), .o(FE_OCPN1823_n_16560) );
in01f04 FE_OCPC1824_n_12030 ( .a(FE_OCP_RBN2284_FE_RN_494_0), .o(FE_OCPN1824_n_12030) );
in01f08 FE_OCPC1825_n_12030 ( .a(FE_OCPN1824_n_12030), .o(FE_OCPN1825_n_12030) );
in01f08 FE_OCPC1827_n_14995 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCPN1827_n_14995) );
in01f10 FE_OCPC1831_n_16949 ( .a(n_16949), .o(FE_OCPN1831_n_16949) );
in01f10 FE_OCPC1832_n_16949 ( .a(FE_OCPN1831_n_16949), .o(FE_OCPN1832_n_16949) );
in01f02 FE_OCPC1833_n_11884 ( .a(n_11884), .o(FE_OCPN1833_n_11884) );
in01f04 FE_OCPC1834_n_11884 ( .a(FE_OCPN1833_n_11884), .o(FE_OCPN1834_n_11884) );
in01f08 FE_OCPC1835_n_16798 ( .a(n_16798), .o(FE_OCPN1835_n_16798) );
in01f10 FE_OCPC1836_n_16798 ( .a(FE_OCPN1835_n_16798), .o(FE_OCPN1836_n_16798) );
in01f40 FE_OCPC1837_n_1238 ( .a(n_1238), .o(FE_OCPN1837_n_1238) );
in01m20 FE_OCPC1838_n_1238 ( .a(FE_OCPN1837_n_1238), .o(FE_OCPN1838_n_1238) );
in01f02 FE_OCPC1839_n_1238 ( .a(FE_OCPN1837_n_1238), .o(FE_OCPN1839_n_1238) );
in01f10 FE_OCPC1840_n_16089 ( .a(n_16089), .o(FE_OCPN1840_n_16089) );
in01f20 FE_OCPC1841_n_16089 ( .a(FE_OCPN1840_n_16089), .o(FE_OCPN1841_n_16089) );
in01f20 FE_OCPC1842_n_16033 ( .a(n_16033), .o(FE_OCPN1842_n_16033) );
in01f20 FE_OCPC1843_n_16033 ( .a(FE_OCPN1842_n_16033), .o(FE_OCPN1843_n_16033) );
in01f06 FE_OCPC1844_n_16427 ( .a(n_16427), .o(FE_OCPN1844_n_16427) );
in01f06 FE_OCPC1845_n_16427 ( .a(FE_OCPN1844_n_16427), .o(TIMEBOOST_net_1) );
in01f10 FE_OCPC1846_n_14981 ( .a(n_14981), .o(FE_OCPN1846_n_14981) );
in01f20 FE_OCPC1847_n_14981 ( .a(FE_OCPN1846_n_14981), .o(FE_OCPN1847_n_14981) );
in01f02 FE_OCPC1848_n_15998 ( .a(n_15998), .o(FE_OCPN1848_n_15998) );
in01f02 FE_OCPC1849_n_15998 ( .a(FE_OCPN1848_n_15998), .o(FE_OCPN1849_n_15998) );
in01f02 FE_OCPC1850_n_15998 ( .a(FE_OCPN1848_n_15998), .o(FE_OCPN1850_n_15998) );
in01f20 FE_OCPC1851_n_16538 ( .a(n_16538), .o(FE_OCPN1851_n_16538) );
in01f20 FE_OCPC1852_n_16538 ( .a(FE_OCPN1851_n_16538), .o(FE_OCPN1852_n_16538) );
in01f20 FE_OCPC1853_n_2071 ( .a(n_2071), .o(FE_OCPN1853_n_2071) );
in01f20 FE_OCPC1854_n_2071 ( .a(FE_OCPN1853_n_2071), .o(FE_OCPN1854_n_2071) );
in01f01 FE_OCPC1855_n_2071 ( .a(FE_OCPN1853_n_2071), .o(FE_OCPN1855_n_2071) );
in01f02 FE_OCPC1856_FE_OFN1774_n_13800 ( .a(FE_OFN1774_n_13800), .o(FE_OCPN1856_FE_OFN1774_n_13800) );
in01f10 FE_OCPC1860_FE_OFN468_n_15534 ( .a(FE_OFN2137_n_15534), .o(FE_OCPN1860_FE_OFN468_n_15534) );
in01f10 FE_OCPC1861_FE_OFN468_n_15534 ( .a(FE_OCPN1860_FE_OFN468_n_15534), .o(FE_OCPN1861_FE_OFN468_n_15534) );
in01f04 FE_OCPC1862_FE_OFN474_n_16992 ( .a(FE_OFN2142_n_16992), .o(FE_OCPN1862_FE_OFN474_n_16992) );
in01f06 FE_OCPC1863_FE_OFN474_n_16992 ( .a(FE_OCPN1862_FE_OFN474_n_16992), .o(FE_OCPN1863_FE_OFN474_n_16992) );
in01f02 FE_OCPC1865_n_12377 ( .a(n_12381), .o(FE_OCPN1865_n_12377) );
in01f04 FE_OCPC1866_n_12377 ( .a(n_12381), .o(FE_OCPN1866_n_12377) );
in01f10 FE_OCPC1871_FE_OFN474_n_16992 ( .a(FE_OFN2142_n_16992), .o(FE_OCPN1871_FE_OFN474_n_16992) );
in01f06 FE_OCPC1872_FE_OFN474_n_16992 ( .a(FE_OCPN1871_FE_OFN474_n_16992), .o(FE_OCPN1872_FE_OFN474_n_16992) );
in01f10 FE_OCPC1873_FE_OFN474_n_16992 ( .a(FE_OCPN1871_FE_OFN474_n_16992), .o(FE_OCPN1873_FE_OFN474_n_16992) );
in01f08 FE_OCPC1875_n_14526 ( .a(n_16460), .o(FE_OCPN1875_n_14526) );
in01f04 FE_OCPC1876_n_13903 ( .a(n_13903), .o(FE_OCPN1876_n_13903) );
in01f04 FE_OCPC1877_n_13903 ( .a(FE_OCPN1876_n_13903), .o(FE_OCPN1877_n_13903) );
in01f06 FE_OCPC1878_FE_OFN470_n_10588 ( .a(FE_OFN2131_n_10588), .o(FE_OCPN1878_FE_OFN470_n_10588) );
in01f06 FE_OCPC1879_FE_OFN470_n_10588 ( .a(FE_OCPN1878_FE_OFN470_n_10588), .o(FE_OCPN1879_FE_OFN470_n_10588) );
in01f08 FE_OCPC1880_n_9991 ( .a(n_9991), .o(FE_OCPN1880_n_9991) );
in01f08 FE_OCPC1881_n_9991 ( .a(FE_OCPN1880_n_9991), .o(FE_OCPN1881_n_9991) );
in01f06 FE_OCPC1882_n_9991 ( .a(FE_OCPN1880_n_9991), .o(FE_OCPN1882_n_9991) );
in01f08 FE_OCPC1883_n_15566 ( .a(n_15566), .o(FE_OCPN1883_n_15566) );
in01f10 FE_OCPC1884_n_15566 ( .a(FE_OCPN1883_n_15566), .o(FE_OCPN1884_n_15566) );
in01f04 FE_OCPC1885_FE_OFN1508_n_15587 ( .a(FE_OFN1508_n_15587), .o(FE_OCPN1885_FE_OFN1508_n_15587) );
in01f06 FE_OCPC1886_FE_OFN1508_n_15587 ( .a(FE_OCPN1885_FE_OFN1508_n_15587), .o(FE_OCPN1886_FE_OFN1508_n_15587) );
in01f08 FE_OCPC1887_FE_OFN473_n_16992 ( .a(FE_OFN2139_n_16992), .o(FE_OCPN1887_FE_OFN473_n_16992) );
in01f10 FE_OCPC1888_FE_OFN473_n_16992 ( .a(FE_OCPN1887_FE_OFN473_n_16992), .o(FE_OCPN1888_FE_OFN473_n_16992) );
in01f02 FE_OCPC1889_n_16553 ( .a(n_16553), .o(FE_OCPN1889_n_16553) );
in01f04 FE_OCPC1890_n_16553 ( .a(FE_OCPN1889_n_16553), .o(FE_OCPN1890_n_16553) );
in01f08 FE_OCPC1891_FE_OFN1727_n_9975 ( .a(FE_OFN1727_n_9975), .o(FE_OCPN1891_FE_OFN1727_n_9975) );
in01f08 FE_OCPC1892_FE_OFN1727_n_9975 ( .a(FE_OCPN1891_FE_OFN1727_n_9975), .o(FE_OCPN1892_FE_OFN1727_n_9975) );
in01f08 FE_OCPC1895_FE_OFN1559_n_12042 ( .a(FE_OFN1559_n_12042), .o(FE_OCPN1895_FE_OFN1559_n_12042) );
in01f08 FE_OCPC1897_n_3231 ( .a(n_3231), .o(FE_OCPN1897_n_3231) );
in01f10 FE_OCPC1898_n_3231 ( .a(FE_OCPN1897_n_3231), .o(FE_OCPN1898_n_3231) );
in01f04 FE_OCPC1899_n_16810 ( .a(n_16810), .o(FE_OCPN1899_n_16810) );
in01f02 FE_OCPC1900_n_16810 ( .a(FE_OCPN1899_n_16810), .o(FE_OCPN1900_n_16810) );
in01f04 FE_OCPC1901_n_16810 ( .a(FE_OCPN1899_n_16810), .o(FE_OCPN1901_n_16810) );
in01f06 FE_OCPC1902_FE_OFN1061_n_16720 ( .a(FE_OFN1061_n_16720), .o(FE_OCPN1902_FE_OFN1061_n_16720) );
in01f06 FE_OCPC1903_FE_OFN1061_n_16720 ( .a(FE_OCPN1902_FE_OFN1061_n_16720), .o(FE_OCPN1903_FE_OFN1061_n_16720) );
in01f04 FE_OCPC1904_n_8927 ( .a(n_8927), .o(FE_OCPN1904_n_8927) );
in01f08 FE_OCPC1905_n_8927 ( .a(FE_OCPN1904_n_8927), .o(FE_OCPN1905_n_8927) );
in01f02 FE_OCPC1907_n_11767 ( .a(FE_OCP_RBN1970_n_11767), .o(FE_OCPN1907_n_11767) );
in01f08 FE_OCPC1908_n_16497 ( .a(FE_OFN2127_n_16497), .o(FE_OCPN1908_n_16497) );
in01f10 FE_OCPC1909_n_16497 ( .a(FE_OCPN1908_n_16497), .o(FE_OCPN1909_n_16497) );
in01f10 FE_OCPC1910_FE_OFN1152_n_13249 ( .a(FE_OFN1152_n_13249), .o(FE_OCPN1910_FE_OFN1152_n_13249) );
in01f10 FE_OCPC1911_FE_OFN1152_n_13249 ( .a(FE_OCPN1910_FE_OFN1152_n_13249), .o(FE_OCPN1911_FE_OFN1152_n_13249) );
in01f04 FE_OCPC1912_FE_OFN1150_n_13249 ( .a(FE_OFN1150_n_13249), .o(FE_OCPN1912_FE_OFN1150_n_13249) );
in01f06 FE_OCPC1913_FE_OFN1150_n_13249 ( .a(FE_OCPN1912_FE_OFN1150_n_13249), .o(FE_OCPN1913_FE_OFN1150_n_13249) );
in01f06 FE_OCPC1914_FE_OFN1522_n_10892 ( .a(FE_OFN1522_n_10892), .o(FE_OCPN1914_FE_OFN1522_n_10892) );
in01f08 FE_OCPC1915_FE_OFN1522_n_10892 ( .a(FE_OCPN1914_FE_OFN1522_n_10892), .o(FE_OCPN1915_FE_OFN1522_n_10892) );
in01f02 FE_OCPC2014_n_10195 ( .a(n_10195), .o(FE_OCPN2014_n_10195) );
in01f04 FE_OCPC2015_n_10195 ( .a(FE_OCPN2014_n_10195), .o(FE_OCPN2015_n_10195) );
in01f06 FE_OCPC2217_n_13997 ( .a(n_13997), .o(FE_OCPN2217_n_13997) );
in01f08 FE_OCPC2218_n_13997 ( .a(FE_OCPN2217_n_13997), .o(FE_OCPN2218_n_13997) );
in01f02 FE_OCPC2219_n_13997 ( .a(FE_OCPN2217_n_13997), .o(FE_OCPN2219_n_13997) );
in01f08 FE_OCPUNCOC1951_FE_OFN697_n_16760 ( .a(FE_OFN697_n_16760), .o(FE_OCPUNCON1951_FE_OFN697_n_16760) );
in01f10 FE_OCPUNCOC1952_FE_OFN697_n_16760 ( .a(FE_OCPUNCON1951_FE_OFN697_n_16760), .o(FE_OCPUNCON1952_FE_OFN697_n_16760) );
in01f08 FE_OCP_DRV_C1949_n_8660 ( .a(FE_OCP_DRV_N2262_n_8660), .o(FE_OCP_DRV_N1949_n_8660) );
in01f10 FE_OCP_DRV_C1950_n_8660 ( .a(FE_OCP_DRV_N1949_n_8660), .o(FE_OCP_DRV_N1950_n_8660) );
in01f04 FE_OCP_DRV_C2261_n_8660 ( .a(n_8660), .o(FE_OCP_DRV_N2261_n_8660) );
in01f06 FE_OCP_DRV_C2262_n_8660 ( .a(FE_OCP_DRV_N2261_n_8660), .o(FE_OCP_DRV_N2262_n_8660) );
in01m01 FE_OCP_RBC1917_wbs_cti_i_1_ ( .a(FE_OCP_RBN1918_wbs_cti_i_1_), .o(FE_OCP_RBN1917_wbs_cti_i_1_) );
in01f80 FE_OCP_RBC1918_wbs_cti_i_1_ ( .a(wbs_cti_i_1_), .o(FE_OCP_RBN1918_wbs_cti_i_1_) );
in01f04 FE_OCP_RBC1921_n_10273 ( .a(n_10273), .o(FE_OCP_RBN1921_n_10273) );
in01f08 FE_OCP_RBC1922_n_10273 ( .a(FE_OCP_RBN1921_n_10273), .o(FE_OCP_RBN1922_n_10273) );
in01f02 FE_OCP_RBC1923_n_10273 ( .a(FE_OCP_RBN1921_n_10273), .o(FE_OCP_RBN1923_n_10273) );
in01f01 FE_OCP_RBC1924_n_10273 ( .a(FE_OCP_RBN1923_n_10273), .o(FE_OCP_RBN1924_n_10273) );
in01f03 FE_OCP_RBC1925_n_10259 ( .a(n_10259), .o(FE_OCP_RBN1925_n_10259) );
in01f02 FE_OCP_RBC1926_n_10259 ( .a(FE_OCP_RBN1925_n_10259), .o(FE_OCP_RBN1926_n_10259) );
in01f02 FE_OCP_RBC1927_n_10259 ( .a(FE_OCP_RBN1925_n_10259), .o(FE_OCP_RBN1927_n_10259) );
in01f04 FE_OCP_RBC1928_n_10259 ( .a(FE_OCP_RBN1925_n_10259), .o(FE_OCP_RBN1928_n_10259) );
in01f10 FE_OCP_RBC1929_parchk_pci_trdy_reg_in ( .a(parchk_pci_trdy_reg_in), .o(FE_OCP_RBN1929_parchk_pci_trdy_reg_in) );
in01m10 FE_OCP_RBC1930_parchk_pci_trdy_reg_in ( .a(FE_OCP_RBN1929_parchk_pci_trdy_reg_in), .o(FE_OCP_RBN1930_parchk_pci_trdy_reg_in) );
in01f08 FE_OCP_RBC1932_FE_OFN1515_n_10538 ( .a(FE_OCP_RBN1966_FE_RN_459_0), .o(FE_OCP_RBN1932_FE_OFN1515_n_10538) );
in01f06 FE_OCP_RBC1933_FE_OFN1515_n_10538 ( .a(FE_OCP_RBN1966_FE_RN_459_0), .o(FE_OCP_RBN1933_FE_OFN1515_n_10538) );
in01f06 FE_OCP_RBC1934_FE_OFN1515_n_10538 ( .a(FE_OCP_RBN1966_FE_RN_459_0), .o(FE_OCP_RBN1934_FE_OFN1515_n_10538) );
in01f08 FE_OCP_RBC1954_FE_RN_462_0 ( .a(FE_RN_462_0), .o(FE_OCP_RBN1954_FE_RN_462_0) );
in01f03 FE_OCP_RBC1955_n_16981 ( .a(n_16981), .o(FE_OCP_RBN1955_n_16981) );
in01f06 FE_OCP_RBC1956_n_16981 ( .a(n_16981), .o(FE_OCP_RBN1956_n_16981) );
in01f04 FE_OCP_RBC1961_FE_OFN1591_n_13741 ( .a(FE_OFN1591_n_13741), .o(FE_OCP_RBN1961_FE_OFN1591_n_13741) );
in01f03 FE_OCP_RBC1962_FE_OFN1591_n_13741 ( .a(FE_OFN1591_n_13741), .o(FE_OCP_RBN1962_FE_OFN1591_n_13741) );
in01f06 FE_OCP_RBC1963_FE_OFN1591_n_13741 ( .a(FE_OFN1591_n_13741), .o(FE_OCP_RBN1963_FE_OFN1591_n_13741) );
in01f08 FE_OCP_RBC1964_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1963_FE_OFN1591_n_13741), .o(FE_OCP_RBN1964_FE_OFN1591_n_13741) );
in01f08 FE_OCP_RBC1965_FE_RN_459_0 ( .a(FE_RN_459_0), .o(FE_OCP_RBN1965_FE_RN_459_0) );
in01f08 FE_OCP_RBC1966_FE_RN_459_0 ( .a(FE_OCP_RBN1965_FE_RN_459_0), .o(FE_OCP_RBN1966_FE_RN_459_0) );
in01f06 FE_OCP_RBC1967_FE_RN_459_0 ( .a(FE_OCP_RBN1965_FE_RN_459_0), .o(FE_OCP_RBN1967_FE_RN_459_0) );
in01f08 FE_OCP_RBC1968_FE_OFN1532_n_10143 ( .a(FE_OFN1532_n_10143), .o(FE_OCP_RBN1968_FE_OFN1532_n_10143) );
in01f08 FE_OCP_RBC1969_FE_OFN1532_n_10143 ( .a(FE_OFN1532_n_10143), .o(FE_OCP_RBN1969_FE_OFN1532_n_10143) );
in01f04 FE_OCP_RBC1970_n_11767 ( .a(n_11767), .o(FE_OCP_RBN1970_n_11767) );
in01f04 FE_OCP_RBC1971_n_11767 ( .a(FE_OCP_RBN1970_n_11767), .o(FE_OCP_RBN1971_n_11767) );
in01f04 FE_OCP_RBC1972_n_11767 ( .a(FE_OCP_RBN1970_n_11767), .o(FE_OCP_RBN1972_n_11767) );
in01f06 FE_OCP_RBC1973_n_12381 ( .a(n_12381), .o(FE_OCP_RBN1973_n_12381) );
in01f01 FE_OCP_RBC1974_n_12381 ( .a(n_12381), .o(FE_OCP_RBN1974_n_12381) );
in01f02 FE_OCP_RBC1975_n_12381 ( .a(n_12381), .o(FE_OCP_RBN1975_n_12381) );
in01f04 FE_OCP_RBC1976_n_12381 ( .a(n_12381), .o(FE_OCP_RBN1976_n_12381) );
in01f01 FE_OCP_RBC1977_n_10273 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCP_RBN1977_n_10273) );
in01f01 FE_OCP_RBC1978_n_10273 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCP_RBN1978_n_10273) );
in01f04 FE_OCP_RBC1979_n_10273 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCP_RBN1979_n_10273) );
in01f02 FE_OCP_RBC1980_n_10273 ( .a(FE_OCP_RBN1922_n_10273), .o(FE_OCP_RBN1980_n_10273) );
in01f02 FE_OCP_RBC1981_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(FE_OCP_RBN1981_FE_OFN1591_n_13741) );
in01f02 FE_OCP_RBC1983_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(FE_OCP_RBN1983_FE_OFN1591_n_13741) );
in01f04 FE_OCP_RBC1984_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(FE_OCP_RBN1984_FE_OFN1591_n_13741) );
in01f06 FE_OCP_RBC1985_FE_OFN1591_n_13741 ( .a(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(FE_OCP_RBN1985_FE_OFN1591_n_13741) );
in01f10 FE_OCP_RBC1994_n_13971 ( .a(n_13971), .o(FE_OCP_RBN1994_n_13971) );
in01f06 FE_OCP_RBC1995_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1995_n_13971) );
in01f06 FE_OCP_RBC1996_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1996_n_13971) );
in01f08 FE_OCP_RBC1997_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1997_n_13971) );
in01f08 FE_OCP_RBC1998_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1998_n_13971) );
in01f04 FE_OCP_RBC1999_n_13971 ( .a(FE_OCP_RBN1994_n_13971), .o(FE_OCP_RBN1999_n_13971) );
in01f08 FE_OCP_RBC2000_n_1403 ( .a(n_1403), .o(FE_OCP_RBN2000_n_1403) );
in01f10 FE_OCP_RBC2003_FE_OFN1026_n_16760 ( .a(FE_OFN1026_n_16760), .o(FE_OCP_RBN2003_FE_OFN1026_n_16760) );
in01f04 FE_OCP_RBC2004_FE_OFN1026_n_16760 ( .a(FE_OFN1026_n_16760), .o(FE_OCP_RBN2004_FE_OFN1026_n_16760) );
in01f08 FE_OCP_RBC2005_FE_RN_459_0 ( .a(FE_OCP_RBN1967_FE_RN_459_0), .o(FE_OCP_RBN2005_FE_RN_459_0) );
in01f06 FE_OCP_RBC2006_FE_RN_459_0 ( .a(FE_OCP_RBN1967_FE_RN_459_0), .o(FE_OCP_RBN2006_FE_RN_459_0) );
in01f02 FE_OCP_RBC2007_n_16698 ( .a(n_16698), .o(FE_OCP_RBN2007_n_16698) );
in01f10 FE_OCP_RBC2008_n_16698 ( .a(n_16698), .o(FE_OCP_RBN2008_n_16698) );
in01f08 FE_OCP_RBC2009_n_16698 ( .a(FE_OCP_RBN2008_n_16698), .o(FE_OCP_RBN2009_n_16698) );
in01f08 FE_OCP_RBC2010_n_16698 ( .a(FE_OCP_RBN2008_n_16698), .o(FE_OCP_RBN2010_n_16698) );
in01f08 FE_OCP_RBC2011_n_16698 ( .a(FE_OCP_RBN2008_n_16698), .o(FE_OCP_RBN2011_n_16698) );
in01f08 FE_OCP_RBC2012_n_16698 ( .a(FE_OCP_RBN2008_n_16698), .o(FE_OCP_RBN2012_n_16698) );
in01f08 FE_OCP_RBC2013_FE_OCPN1895_FE_OFN1559_n_12042 ( .a(FE_OCPN1895_FE_OFN1559_n_12042), .o(FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042) );
in01f04 FE_OCP_RBC2016_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2016_n_16970) );
in01f02 FE_OCP_RBC2017_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2017_n_16970) );
in01f01 FE_OCP_RBC2018_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2018_n_16970) );
in01f01 FE_OCP_RBC2019_n_16970 ( .a(n_16970), .o(FE_OCP_RBN2019_n_16970) );
in01f02 FE_OCP_RBC2220_n_15347 ( .a(n_15347), .o(FE_OCP_RBN2220_n_15347) );
in01f02 FE_OCP_RBC2221_n_15347 ( .a(n_15347), .o(FE_OCP_RBN2221_n_15347) );
in01f08 FE_OCP_RBC2222_n_15347 ( .a(n_15347), .o(FE_OCP_RBN2222_n_15347) );
in01f06 FE_OCP_RBC2223_n_15347 ( .a(n_15347), .o(FE_OCP_RBN2223_n_15347) );
in01f06 FE_OCP_RBC2224_n_16322 ( .a(n_16322), .o(FE_OCP_RBN2224_n_16322) );
in01f06 FE_OCP_RBC2225_n_16322 ( .a(n_16322), .o(FE_OCP_RBN2225_n_16322) );
in01f06 FE_OCP_RBC2226_g75174_p ( .a(g75174_p), .o(FE_OCP_RBN2226_g75174_p) );
in01f02 FE_OCP_RBC2227_g75174_p ( .a(g75174_p), .o(FE_OCP_RBN2227_g75174_p) );
in01f02 FE_OCP_RBC2228_n_15969 ( .a(n_15969), .o(FE_OCP_RBN2228_n_15969) );
in01f04 FE_OCP_RBC2229_n_15969 ( .a(FE_OCP_RBN2228_n_15969), .o(FE_OCP_RBN2229_n_15969) );
in01f02 FE_OCP_RBC2231_FE_RN_390_0 ( .a(FE_RN_390_0), .o(FE_OCP_RBN2231_FE_RN_390_0) );
in01f03 FE_OCP_RBC2232_n_16273 ( .a(n_16273), .o(FE_OCP_RBN2232_n_16273) );
in01f02 FE_OCP_RBC2233_n_16273 ( .a(n_16273), .o(FE_OCP_RBN2233_n_16273) );
in01f02 FE_OCP_RBC2237_g74749_p ( .a(g74749_p), .o(FE_OCP_RBN2237_g74749_p) );
in01f06 FE_OCP_RBC2238_g74749_p ( .a(g74749_p), .o(FE_OCP_RBN2238_g74749_p) );
in01f06 FE_OCP_RBC2239_g74749_p ( .a(g74749_p), .o(FE_OCP_RBN2239_g74749_p) );
in01s01 FE_OCP_RBC2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_ ( .a(FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .o(FE_OCP_RBN2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_) );
in01f80 FE_OCP_RBC2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_ ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .o(FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_) );
in01f40 FE_OCP_RBC2270_g75061_p ( .a(g75061_p), .o(FE_OCP_RBN2270_g75061_p) );
in01f08 FE_OCP_RBC2271_g75061_p ( .a(g75061_p), .o(FE_OCP_RBN2271_g75061_p) );
in01f01 FE_OCP_RBC2272_n_10268 ( .a(n_10268), .o(FE_OCP_RBN2272_n_10268) );
in01f04 FE_OCP_RBC2273_n_10268 ( .a(n_10268), .o(FE_OCP_RBN2273_n_10268) );
in01f08 FE_OCP_RBC2274_n_10268 ( .a(FE_OCP_RBN2273_n_10268), .o(FE_OCP_RBN2274_n_10268) );
in01f02 FE_OCP_RBC2275_n_10268 ( .a(FE_OCP_RBN2273_n_10268), .o(FE_OCP_RBN2275_n_10268) );
in01f80 FE_OCP_RBC2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_ ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_), .o(FE_OCP_RBN2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_) );
in01f04 FE_OCP_RBC2278_n_16974 ( .a(n_16974), .o(FE_OCP_RBN2278_n_16974) );
in01f02 FE_OCP_RBC2279_n_16974 ( .a(n_16974), .o(FE_OCP_RBN2279_n_16974) );
in01f02 FE_OCP_RBC2280_g74996_p ( .a(g74996_p), .o(FE_OCP_RBN2280_g74996_p) );
in01f02 FE_OCP_RBC2281_g74996_p ( .a(g74996_p), .o(FE_OCP_RBN2281_g74996_p) );
in01f02 FE_OCP_RBC2282_g74996_p ( .a(g74996_p), .o(FE_OCP_RBN2282_g74996_p) );
in01f02 FE_OCP_RBC2283_g74996_p ( .a(g74996_p), .o(FE_OCP_RBN2283_g74996_p) );
in01f02 FE_OCP_RBC2284_FE_RN_494_0 ( .a(FE_RN_494_0), .o(FE_OCP_RBN2284_FE_RN_494_0) );
in01f04 FE_OCP_RBC2285_FE_RN_494_0 ( .a(FE_RN_494_0), .o(FE_OCP_RBN2285_FE_RN_494_0) );
in01f08 FE_OCP_RBC2286_FE_RN_494_0 ( .a(FE_OCP_RBN2285_FE_RN_494_0), .o(FE_OCP_RBN2286_FE_RN_494_0) );
in01s01 FE_OCP_RBC2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_ ( .a(FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .o(FE_OCP_RBN2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_) );
in01f40 FE_OCP_RBC2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_ ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .o(FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_) );
in01f06 FE_OCP_RBC2291_FE_OFN1575_n_12028 ( .a(FE_OFN1575_n_12028), .o(FE_OCP_RBN2291_FE_OFN1575_n_12028) );
in01f06 FE_OCP_RBC2292_FE_OFN1575_n_12028 ( .a(FE_OFN1575_n_12028), .o(FE_OCP_RBN2292_FE_OFN1575_n_12028) );
in01f04 FE_OCP_RBC2293_FE_OFN1581_n_12306 ( .a(FE_OFN1581_n_12306), .o(FE_OCP_RBN2293_FE_OFN1581_n_12306) );
in01f08 FE_OFC1001_n_15978 ( .a(FE_OFN997_n_15978), .o(FE_OFN1001_n_15978) );
in01f02 FE_OFC1002_n_2047 ( .a(n_2047), .o(FE_OFN1002_n_2047) );
in01f08 FE_OFC1003_n_2047 ( .a(FE_OFN1002_n_2047), .o(FE_OFN1003_n_2047) );
in01f08 FE_OFC1004_n_16288 ( .a(n_16288), .o(FE_OFN1004_n_16288) );
in01f10 FE_OFC1005_n_16288 ( .a(FE_OFN1004_n_16288), .o(FE_OFN1005_n_16288) );
in01f10 FE_OFC1006_n_16288 ( .a(FE_OFN1004_n_16288), .o(FE_OFN1006_n_16288) );
in01f02 FE_OFC1007_n_4734 ( .a(n_4734), .o(FE_OFN1007_n_4734) );
in01f03 FE_OFC1008_n_4734 ( .a(n_4734), .o(FE_OFN1008_n_4734) );
in01f08 FE_OFC1009_n_4734 ( .a(n_4734), .o(FE_OFN1009_n_4734) );
in01f06 FE_OFC1010_n_4734 ( .a(FE_OFN1008_n_4734), .o(FE_OFN1010_n_4734) );
in01f04 FE_OFC1011_n_4734 ( .a(FE_OFN1008_n_4734), .o(FE_OFN1011_n_4734) );
in01f08 FE_OFC1012_n_4734 ( .a(FE_OFN1009_n_4734), .o(FE_OFN1012_n_4734) );
in01f10 FE_OFC1013_n_4734 ( .a(FE_OFN1009_n_4734), .o(FE_OFN1013_n_4734) );
in01f08 FE_OFC1014_n_2053 ( .a(n_2053), .o(FE_OFN1014_n_2053) );
in01f06 FE_OFC1015_n_2053 ( .a(FE_OFN1014_n_2053), .o(FE_OFN1015_n_2053) );
in01f10 FE_OFC1016_n_2053 ( .a(FE_OFN1014_n_2053), .o(FE_OFN1016_n_2053) );
in01f06 FE_OFC1017_n_2053 ( .a(FE_OFN1014_n_2053), .o(FE_OFN1017_n_2053) );
in01f08 FE_OFC1018_n_11877 ( .a(n_11877), .o(FE_OFN1018_n_11877) );
in01f04 FE_OFC1019_n_11877 ( .a(n_11877), .o(FE_OFN1019_n_11877) );
in01f10 FE_OFC1020_n_11877 ( .a(n_11877), .o(FE_OFN1020_n_11877) );
in01f06 FE_OFC1021_n_11877 ( .a(FE_OFN1018_n_11877), .o(FE_OFN1021_n_11877) );
in01f10 FE_OFC1022_n_11877 ( .a(FE_OFN1018_n_11877), .o(FE_OFN1022_n_11877) );
in01m08 FE_OFC1023_n_11877 ( .a(FE_OFN1019_n_11877), .o(FE_OFN1023_n_11877) );
in01f01 FE_OFC1024_n_11877 ( .a(FE_OFN1019_n_11877), .o(FE_OFN1024_n_11877) );
in01f08 FE_OFC1025_n_11877 ( .a(FE_OFN1020_n_11877), .o(FE_OFN1025_n_11877) );
in01f08 FE_OFC1028_n_4732 ( .a(n_4732), .o(FE_OFN1028_n_4732) );
in01f20 FE_OFC1029_n_4732 ( .a(n_4732), .o(FE_OFN1029_n_4732) );
in01f10 FE_OFC1030_n_4732 ( .a(n_4732), .o(FE_OFN1030_n_4732) );
in01f08 FE_OFC1031_n_4732 ( .a(FE_OFN1028_n_4732), .o(FE_OFN1031_n_4732) );
in01f08 FE_OFC1032_n_4732 ( .a(FE_OFN1029_n_4732), .o(FE_OFN1032_n_4732) );
in01f06 FE_OFC1033_n_4732 ( .a(FE_OFN1030_n_4732), .o(FE_OFN1033_n_4732) );
in01f10 FE_OFC1034_n_4732 ( .a(FE_OFN1030_n_4732), .o(FE_OFN1034_n_4732) );
in01f01 FE_OFC1035_n_4732 ( .a(FE_OFN1028_n_4732), .o(FE_OFN1035_n_4732) );
in01m08 FE_OFC1036_n_4732 ( .a(FE_OFN1028_n_4732), .o(FE_OFN1036_n_4732) );
in01m20 FE_OFC1037_n_4732 ( .a(FE_OFN1029_n_4732), .o(FE_OFN1037_n_4732) );
in01f04 FE_OFC1038_n_2037 ( .a(n_2037), .o(FE_OFN1038_n_2037) );
in01f01 FE_OFC1039_n_2037 ( .a(n_2037), .o(FE_OFN1039_n_2037) );
in01m01 FE_OFC1040_n_2037 ( .a(n_2037), .o(FE_OFN1040_n_2037) );
in01m08 FE_OFC1041_n_2037 ( .a(FE_OFN1038_n_2037), .o(FE_OFN1041_n_2037) );
in01f04 FE_OFC1042_n_2037 ( .a(FE_OFN1038_n_2037), .o(FE_OFN1042_n_2037) );
in01f04 FE_OFC1043_n_2037 ( .a(FE_OFN1039_n_2037), .o(FE_OFN1043_n_2037) );
in01f04 FE_OFC1044_n_2037 ( .a(FE_OFN1040_n_2037), .o(FE_OFN1044_n_2037) );
in01f20 FE_OFC1045_n_16657 ( .a(n_16657), .o(FE_OFN1045_n_16657) );
in01f40 FE_OFC1046_n_16657 ( .a(FE_OFN1045_n_16657), .o(FE_OFN1046_n_16657) );
in01m10 FE_OFC1047_n_16657 ( .a(n_16657), .o(FE_OFN1047_n_16657) );
in01f06 FE_OFC1048_n_16657 ( .a(n_16657), .o(FE_OFN1048_n_16657) );
in01f10 FE_OFC1049_n_16657 ( .a(FE_OFN1048_n_16657), .o(FE_OFN1049_n_16657) );
in01m10 FE_OFC1050_n_16657 ( .a(FE_OFN1047_n_16657), .o(FE_OFN1050_n_16657) );
in01f10 FE_OFC1051_n_16657 ( .a(FE_OFN1047_n_16657), .o(FE_OFN1051_n_16657) );
in01f10 FE_OFC1052_n_4727 ( .a(n_4727), .o(FE_OFN1052_n_4727) );
in01f08 FE_OFC1053_n_4727 ( .a(n_4727), .o(FE_OFN1053_n_4727) );
in01f10 FE_OFC1054_n_4727 ( .a(n_4727), .o(FE_OFN1054_n_4727) );
in01f06 FE_OFC1055_n_4727 ( .a(FE_OFN1053_n_4727), .o(FE_OFN1055_n_4727) );
in01f10 FE_OFC1056_n_4727 ( .a(FE_OFN1053_n_4727), .o(FE_OFN1056_n_4727) );
in01f20 FE_OFC1057_n_4727 ( .a(FE_OFN1054_n_4727), .o(FE_OFN1057_n_4727) );
in01m04 FE_OFC1058_n_4727 ( .a(FE_OFN1054_n_4727), .o(FE_OFN1058_n_4727) );
in01f04 FE_OFC1059_n_4727 ( .a(FE_OFN1054_n_4727), .o(FE_OFN1059_n_4727) );
in01f08 FE_OFC1061_n_16720 ( .a(FE_OFN1060_n_16720), .o(TIMEBOOST_net_5) );
in01f10 FE_OFC1062_n_15808 ( .a(n_15808), .o(FE_OFN1062_n_15808) );
in01f20 FE_OFC1063_n_15808 ( .a(FE_OFN1062_n_15808), .o(FE_OFN1063_n_15808) );
in01f10 FE_OFC1064_n_15808 ( .a(n_15808), .o(FE_OFN1064_n_15808) );
in01f08 FE_OFC1065_n_15808 ( .a(FE_OFN1064_n_15808), .o(FE_OFN1065_n_15808) );
in01f10 FE_OFC1066_n_15808 ( .a(FE_OFN1064_n_15808), .o(FE_OFN1066_n_15808) );
in01f10 FE_OFC1067_n_15729 ( .a(n_15729), .o(FE_OFN1067_n_15729) );
in01f04 FE_OFC1068_n_15729 ( .a(FE_OFN1067_n_15729), .o(FE_OFN1068_n_15729) );
in01f10 FE_OFC1069_n_15729 ( .a(FE_OFN1067_n_15729), .o(FE_OFN1069_n_15729) );
in01f10 FE_OFC1070_n_15729 ( .a(FE_OFN1067_n_15729), .o(FE_OFN1070_n_15729) );
in01f08 FE_OFC1071_n_15729 ( .a(FE_OFN1067_n_15729), .o(FE_OFN1071_n_15729) );
in01f10 FE_OFC1072_n_4740 ( .a(n_4740), .o(FE_OFN1072_n_4740) );
in01f40 FE_OFC1073_n_4740 ( .a(n_4740), .o(FE_OFN1073_n_4740) );
in01f20 FE_OFC1074_n_4740 ( .a(FE_OFN1073_n_4740), .o(FE_OFN1074_n_4740) );
in01f10 FE_OFC1075_n_4740 ( .a(FE_OFN1073_n_4740), .o(FE_OFN1075_n_4740) );
in01f20 FE_OFC1076_n_4740 ( .a(FE_OFN1073_n_4740), .o(FE_OFN1076_n_4740) );
in01f20 FE_OFC1077_n_4740 ( .a(FE_OFN1073_n_4740), .o(FE_OFN1077_n_4740) );
in01f06 FE_OFC1078_n_4778 ( .a(n_4778), .o(FE_OFN1078_n_4778) );
in01f10 FE_OFC1079_n_4778 ( .a(FE_OFN1078_n_4778), .o(FE_OFN1079_n_4778) );
in01f10 FE_OFC1080_n_13221 ( .a(n_13221), .o(FE_OFN1080_n_13221) );
in01f10 FE_OFC1081_n_13221 ( .a(n_13221), .o(FE_OFN1081_n_13221) );
in01f08 FE_OFC1082_n_13221 ( .a(FE_OFN1080_n_13221), .o(FE_OFN1082_n_13221) );
in01f10 FE_OFC1083_n_13221 ( .a(FE_OFN1080_n_13221), .o(FE_OFN1083_n_13221) );
in01f10 FE_OFC1084_n_13221 ( .a(FE_OFN1081_n_13221), .o(FE_OFN1084_n_13221) );
in01f10 FE_OFC1085_n_13221 ( .a(FE_OFN1081_n_13221), .o(FE_OFN1085_n_13221) );
in01f04 FE_OFC1086_g64577_p ( .a(g64577_p), .o(FE_OFN1086_g64577_p) );
in01f20 FE_OFC1087_g64577_p ( .a(g64577_p), .o(FE_OFN1087_g64577_p) );
in01f08 FE_OFC1088_g64577_p ( .a(g64577_p), .o(FE_OFN1088_g64577_p) );
in01f08 FE_OFC1089_g64577_p ( .a(g64577_p), .o(FE_OFN1089_g64577_p) );
in01f06 FE_OFC1090_g64577_p ( .a(FE_OFN1086_g64577_p), .o(FE_OFN1090_g64577_p) );
in01f10 FE_OFC1091_g64577_p ( .a(FE_OFN1087_g64577_p), .o(FE_OFN1091_g64577_p) );
in01f20 FE_OFC1092_g64577_p ( .a(FE_OFN1087_g64577_p), .o(FE_OFN1092_g64577_p) );
in01f08 FE_OFC1093_g64577_p ( .a(FE_OFN1087_g64577_p), .o(FE_OFN1093_g64577_p) );
in01f03 FE_OFC1094_g64577_p ( .a(FE_OFN1087_g64577_p), .o(FE_OFN1094_g64577_p) );
in01f03 FE_OFC1095_g64577_p ( .a(FE_OFN1089_g64577_p), .o(FE_OFN1095_g64577_p) );
in01f08 FE_OFC1096_g64577_p ( .a(FE_OFN1089_g64577_p), .o(FE_OFN1096_g64577_p) );
in01f10 FE_OFC1097_g64577_p ( .a(FE_OFN1089_g64577_p), .o(FE_OFN1097_g64577_p) );
in01f08 FE_OFC1098_g64577_p ( .a(FE_OFN1090_g64577_p), .o(FE_OFN1098_g64577_p) );
in01f03 FE_OFC1099_g64577_p ( .a(FE_OFN1090_g64577_p), .o(FE_OFN1099_g64577_p) );
in01f02 FE_OFC1100_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1100_g64577_p) );
in01f20 FE_OFC1101_g64577_p ( .a(FE_OFN1091_g64577_p), .o(FE_OFN1101_g64577_p) );
in01f08 FE_OFC1102_g64577_p ( .a(FE_OFN1091_g64577_p), .o(FE_OFN1102_g64577_p) );
in01f08 FE_OFC1103_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1103_g64577_p) );
in01f06 FE_OFC1104_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1104_g64577_p) );
in01f20 FE_OFC1105_g64577_p ( .a(FE_OFN1092_g64577_p), .o(FE_OFN1105_g64577_p) );
in01f08 FE_OFC1106_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1106_g64577_p) );
in01f03 FE_OFC1107_g64577_p ( .a(FE_OFN1088_g64577_p), .o(FE_OFN1107_g64577_p) );
in01f10 FE_OFC1108_g64577_p ( .a(FE_OFN1096_g64577_p), .o(FE_OFN1108_g64577_p) );
in01f10 FE_OFC1109_g64577_p ( .a(FE_OFN1097_g64577_p), .o(FE_OFN1109_g64577_p) );
in01f10 FE_OFC1110_g64577_p ( .a(FE_OFN1093_g64577_p), .o(FE_OFN1110_g64577_p) );
in01f06 FE_OFC1111_g64577_p ( .a(FE_OFN1093_g64577_p), .o(FE_OFN1111_g64577_p) );
in01f06 FE_OFC1112_g64577_p ( .a(FE_OFN1102_g64577_p), .o(FE_OFN1112_g64577_p) );
in01f08 FE_OFC1113_g64577_p ( .a(FE_OFN1103_g64577_p), .o(FE_OFN1113_g64577_p) );
in01f06 FE_OFC1114_g64577_p ( .a(FE_OFN1103_g64577_p), .o(FE_OFN1114_g64577_p) );
in01f08 FE_OFC1115_g64577_p ( .a(FE_OFN1101_g64577_p), .o(FE_OFN1115_g64577_p) );
in01f06 FE_OFC1116_g64577_p ( .a(FE_OFN1102_g64577_p), .o(FE_OFN1116_g64577_p) );
in01f20 FE_OFC1117_g64577_p ( .a(FE_OFN1105_g64577_p), .o(FE_OFN1117_g64577_p) );
in01f08 FE_OFC1118_g64577_p ( .a(FE_OFN1108_g64577_p), .o(FE_OFN1118_g64577_p) );
in01f10 FE_OFC1119_g64577_p ( .a(FE_OFN1109_g64577_p), .o(FE_OFN1119_g64577_p) );
in01f10 FE_OFC1120_g64577_p ( .a(FE_OFN1109_g64577_p), .o(FE_OFN1120_g64577_p) );
in01f10 FE_OFC1121_g64577_p ( .a(FE_OFN1101_g64577_p), .o(FE_OFN1121_g64577_p) );
in01f06 FE_OFC1122_g64577_p ( .a(FE_OFN1102_g64577_p), .o(FE_OFN1122_g64577_p) );
in01f08 FE_OFC1123_g64577_p ( .a(FE_OFN1102_g64577_p), .o(FE_OFN1123_g64577_p) );
in01f08 FE_OFC1124_g64577_p ( .a(FE_OFN1105_g64577_p), .o(FE_OFN1124_g64577_p) );
in01f10 FE_OFC1125_g64577_p ( .a(FE_OFN1105_g64577_p), .o(FE_OFN1125_g64577_p) );
in01f10 FE_OFC1126_g64577_p ( .a(FE_OFN1110_g64577_p), .o(FE_OFN1126_g64577_p) );
in01f02 FE_OFC1127_g64577_p ( .a(FE_OFN1111_g64577_p), .o(FE_OFN1127_g64577_p) );
in01f08 FE_OFC1128_g64577_p ( .a(FE_OFN1111_g64577_p), .o(FE_OFN1128_g64577_p) );
in01f08 FE_OFC1129_g64577_p ( .a(FE_OFN1108_g64577_p), .o(FE_OFN1129_g64577_p) );
in01f06 FE_OFC1130_g64577_p ( .a(FE_OFN1101_g64577_p), .o(FE_OFN1130_g64577_p) );
in01f10 FE_OFC1131_g64577_p ( .a(FE_OFN1101_g64577_p), .o(FE_OFN1131_g64577_p) );
in01f08 FE_OFC1132_g64577_p ( .a(FE_OFN1110_g64577_p), .o(FE_OFN1132_g64577_p) );
in01f10 FE_OFC1133_g64577_p ( .a(FE_OFN1110_g64577_p), .o(FE_OFN1133_g64577_p) );
in01f10 FE_OFC1134_g64577_p ( .a(FE_OFN1113_g64577_p), .o(FE_OFN1134_g64577_p) );
in01f10 FE_OFC1135_g64577_p ( .a(FE_OFN1114_g64577_p), .o(FE_OFN1135_g64577_p) );
in01f10 FE_OFC1136_g64577_p ( .a(FE_OFN1108_g64577_p), .o(FE_OFN1136_g64577_p) );
in01f06 FE_OFC1137_g64577_p ( .a(FE_OFN1108_g64577_p), .o(FE_OFN1137_g64577_p) );
in01f08 FE_OFC1138_g64577_p ( .a(FE_OFN1107_g64577_p), .o(FE_OFN1138_g64577_p) );
in01f08 FE_OFC1139_g64577_p ( .a(FE_OFN1138_g64577_p), .o(FE_OFN1139_g64577_p) );
in01f08 FE_OFC1140_g64577_p ( .a(FE_OFN1138_g64577_p), .o(FE_OFN1140_g64577_p) );
in01m20 FE_OFC1141_n_15261 ( .a(n_15261), .o(FE_OFN1141_n_15261) );
in01f10 FE_OFC1142_n_15261 ( .a(FE_OFN1141_n_15261), .o(FE_OFN1142_n_15261) );
in01f10 FE_OFC1143_n_15261 ( .a(FE_OFN1141_n_15261), .o(FE_OFN1143_n_15261) );
in01f08 FE_OFC1144_n_15261 ( .a(FE_OFN1141_n_15261), .o(FE_OFN1144_n_15261) );
in01f08 FE_OFC1145_n_15261 ( .a(FE_OFN1141_n_15261), .o(FE_OFN1145_n_15261) );
in01f40 FE_OFC1146_n_13249 ( .a(n_13249), .o(FE_OFN1146_n_13249) );
in01f20 FE_OFC1147_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1147_n_13249) );
in01f20 FE_OFC1148_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1148_n_13249) );
in01f08 FE_OFC1149_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1149_n_13249) );
in01f10 FE_OFC1150_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1150_n_13249) );
in01m10 FE_OFC1151_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1151_n_13249) );
in01f10 FE_OFC1152_n_13249 ( .a(FE_OFN1146_n_13249), .o(FE_OFN1152_n_13249) );
in01f10 FE_OFC1153_n_3464 ( .a(n_3464), .o(FE_OFN1153_n_3464) );
in01f10 FE_OFC1154_n_3464 ( .a(FE_OFN1153_n_3464), .o(FE_OFN1154_n_3464) );
in01f20 FE_OFC1155_n_3464 ( .a(FE_OFN1153_n_3464), .o(FE_OFN1155_n_3464) );
in01f04 FE_OFC1156_n_7498 ( .a(n_7498), .o(FE_OFN1156_n_7498) );
in01f20 FE_OFC1157_n_15325 ( .a(n_15325), .o(FE_OFN1157_n_15325) );
in01f10 FE_OFC1158_n_15325 ( .a(FE_OFN1157_n_15325), .o(FE_OFN1158_n_15325) );
in01f20 FE_OFC1159_n_15325 ( .a(FE_OFN1157_n_15325), .o(FE_OFN1159_n_15325) );
in01f06 FE_OFC1160_n_5615 ( .a(n_5592), .o(FE_OFN1160_n_5615) );
in01f08 FE_OFC1161_n_5615 ( .a(n_5592), .o(FE_OFN1161_n_5615) );
in01f06 FE_OFC1162_n_5615 ( .a(n_5592), .o(FE_OFN1162_n_5615) );
in01f08 FE_OFC1163_n_5615 ( .a(FE_OFN1160_n_5615), .o(FE_OFN1163_n_5615) );
in01f08 FE_OFC1164_n_5615 ( .a(FE_OFN1161_n_5615), .o(FE_OFN1164_n_5615) );
in01f06 FE_OFC1165_n_5615 ( .a(FE_OFN1161_n_5615), .o(FE_OFN1165_n_5615) );
in01f08 FE_OFC1166_n_5615 ( .a(FE_OFN1162_n_5615), .o(FE_OFN1166_n_5615) );
in01f40 FE_OFC1167_n_5592 ( .a(n_5592), .o(FE_OFN1167_n_5592) );
in01f10 FE_OFC1168_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1168_n_5592) );
in01f10 FE_OFC1169_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1169_n_5592) );
in01f10 FE_OFC1170_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1170_n_5592) );
in01f20 FE_OFC1171_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1171_n_5592) );
in01f04 FE_OFC1172_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1172_n_5592) );
in01f10 FE_OFC1173_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1173_n_5592) );
in01f20 FE_OFC1174_n_5592 ( .a(FE_OFN1167_n_5592), .o(FE_OFN1174_n_5592) );
in01f08 FE_OFC1175_n_3476 ( .a(n_3476), .o(FE_OFN1175_n_3476) );
in01f08 FE_OFC1176_n_3476 ( .a(n_3476), .o(FE_OFN1176_n_3476) );
in01f10 FE_OFC1177_n_3476 ( .a(n_3476), .o(FE_OFN1177_n_3476) );
in01f08 FE_OFC1178_n_3476 ( .a(n_3476), .o(FE_OFN1178_n_3476) );
in01f10 FE_OFC1179_n_3476 ( .a(FE_OFN1178_n_3476), .o(FE_OFN1179_n_3476) );
in01f08 FE_OFC1180_n_3476 ( .a(FE_OFN1175_n_3476), .o(FE_OFN1180_n_3476) );
in01f10 FE_OFC1181_n_3476 ( .a(FE_OFN1175_n_3476), .o(FE_OFN1181_n_3476) );
in01f08 FE_OFC1182_n_3476 ( .a(FE_OFN1176_n_3476), .o(FE_OFN1182_n_3476) );
in01f10 FE_OFC1183_n_3476 ( .a(FE_OFN1176_n_3476), .o(FE_OFN1183_n_3476) );
in01f10 FE_OFC1184_n_3476 ( .a(FE_OFN1177_n_3476), .o(FE_OFN1184_n_3476) );
in01f10 FE_OFC1185_n_3476 ( .a(FE_OFN1177_n_3476), .o(FE_OFN1185_n_3476) );
in01f06 FE_OFC1186_n_3476 ( .a(FE_OFN1178_n_3476), .o(FE_OFN1186_n_3476) );
in01f08 FE_OFC1187_n_5742 ( .a(n_5742), .o(FE_OFN1187_n_5742) );
in01f06 FE_OFC1188_n_5742 ( .a(FE_OFN1187_n_5742), .o(FE_OFN1188_n_5742) );
in01f10 FE_OFC1189_n_5742 ( .a(FE_OFN1187_n_5742), .o(FE_OFN1189_n_5742) );
in01f04 FE_OFC1190_n_6935 ( .a(n_6935), .o(FE_OFN1190_n_6935) );
in01f20 FE_OFC1191_n_6935 ( .a(n_6935), .o(FE_OFN1191_n_6935) );
in01f40 FE_OFC1192_n_6935 ( .a(FE_OFN1191_n_6935), .o(FE_OFN1192_n_6935) );
in01f08 FE_OFC1193_n_6935 ( .a(FE_OFN1190_n_6935), .o(FE_OFN1193_n_6935) );
in01f04 FE_OFC1194_n_6935 ( .a(FE_OFN1190_n_6935), .o(FE_OFN1194_n_6935) );
in01f02 FE_OFC1195_n_4090 ( .a(n_4090), .o(FE_OFN1195_n_4090) );
in01f02 FE_OFC1196_n_4090 ( .a(FE_OFN1195_n_4090), .o(FE_OFN1196_n_4090) );
in01f02 FE_OFC1197_n_4090 ( .a(FE_OFN1195_n_4090), .o(FE_OFN1197_n_4090) );
in01f02 FE_OFC1198_n_4090 ( .a(n_4090), .o(FE_OFN1198_n_4090) );
in01f04 FE_OFC1199_n_4090 ( .a(n_4090), .o(FE_OFN1199_n_4090) );
in01f06 FE_OFC1200_n_4090 ( .a(FE_OFN1198_n_4090), .o(FE_OFN1200_n_4090) );
in01f04 FE_OFC1201_n_4090 ( .a(n_4090), .o(FE_OFN1201_n_4090) );
in01f08 FE_OFC1202_n_4090 ( .a(FE_OFN1201_n_4090), .o(FE_OFN1202_n_4090) );
in01f04 FE_OFC1203_n_4090 ( .a(FE_OFN1199_n_4090), .o(FE_OFN1203_n_4090) );
in01f04 FE_OFC1204_n_4090 ( .a(FE_OFN1199_n_4090), .o(FE_OFN1204_n_4090) );
in01f08 FE_OFC1205_n_6356 ( .a(n_6356), .o(FE_OFN1205_n_6356) );
in01f06 FE_OFC1206_n_6356 ( .a(FE_OFN1205_n_6356), .o(FE_OFN1206_n_6356) );
in01f08 FE_OFC1207_n_6356 ( .a(FE_OFN1205_n_6356), .o(FE_OFN1207_n_6356) );
in01f08 FE_OFC1208_n_6356 ( .a(FE_OFN1205_n_6356), .o(FE_OFN1208_n_6356) );
in01f02 FE_OFC1209_n_4151 ( .a(n_4151), .o(FE_OFN1209_n_4151) );
in01f08 FE_OFC1210_n_4151 ( .a(n_4151), .o(FE_OFN1210_n_4151) );
in01f04 FE_OFC1211_n_4151 ( .a(n_4151), .o(FE_OFN1211_n_4151) );
in01f08 FE_OFC1212_n_4151 ( .a(FE_OFN1210_n_4151), .o(FE_OFN1212_n_4151) );
in01f08 FE_OFC1213_n_4151 ( .a(FE_OFN1210_n_4151), .o(FE_OFN1213_n_4151) );
in01f06 FE_OFC1214_n_4151 ( .a(FE_OFN1209_n_4151), .o(FE_OFN1214_n_4151) );
in01f06 FE_OFC1215_n_4151 ( .a(FE_OFN1211_n_4151), .o(FE_OFN1215_n_4151) );
in01f04 FE_OFC1216_n_4151 ( .a(FE_OFN1211_n_4151), .o(FE_OFN1216_n_4151) );
in01f08 FE_OFC1217_n_6886 ( .a(n_6886), .o(FE_OFN1217_n_6886) );
in01f08 FE_OFC1218_n_6886 ( .a(FE_OFN1217_n_6886), .o(FE_OFN1218_n_6886) );
in01m08 FE_OFC1219_n_6886 ( .a(FE_OFN1217_n_6886), .o(FE_OFN1219_n_6886) );
in01f40 FE_OFC1220_n_6391 ( .a(n_6391), .o(FE_OFN1220_n_6391) );
in01f40 FE_OFC1221_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1221_n_6391) );
in01f20 FE_OFC1222_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1222_n_6391) );
in01f20 FE_OFC1223_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1223_n_6391) );
in01f08 FE_OFC1224_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1224_n_6391) );
in01f06 FE_OFC1225_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1225_n_6391) );
in01f02 FE_OFC1226_n_6391 ( .a(FE_OFN1220_n_6391), .o(FE_OFN1226_n_6391) );
in01f20 FE_OFC1227_n_6391 ( .a(FE_OFN1221_n_6391), .o(FE_OFN1227_n_6391) );
in01f20 FE_OFC1228_n_6391 ( .a(FE_OFN1221_n_6391), .o(FE_OFN1228_n_6391) );
in01f20 FE_OFC1229_n_6391 ( .a(FE_OFN1222_n_6391), .o(FE_OFN1229_n_6391) );
in01f10 FE_OFC1230_n_6391 ( .a(FE_OFN1227_n_6391), .o(FE_OFN1230_n_6391) );
in01f10 FE_OFC1231_n_6391 ( .a(FE_OFN1227_n_6391), .o(FE_OFN1231_n_6391) );
in01f10 FE_OFC1232_n_6391 ( .a(FE_OFN1227_n_6391), .o(FE_OFN1232_n_6391) );
in01f10 FE_OFC1233_n_6391 ( .a(FE_OFN1228_n_6391), .o(FE_OFN1233_n_6391) );
in01f20 FE_OFC1234_n_6391 ( .a(FE_OFN1229_n_6391), .o(FE_OFN1234_n_6391) );
in01f10 FE_OFC1235_n_6391 ( .a(FE_OFN1228_n_6391), .o(FE_OFN1235_n_6391) );
in01f10 FE_OFC1236_n_6391 ( .a(FE_OFN1228_n_6391), .o(FE_OFN1236_n_6391) );
in01m01 FE_OFC1237_n_4092 ( .a(n_4092), .o(FE_OFN1237_n_4092) );
in01f08 FE_OFC1238_n_4092 ( .a(n_4092), .o(FE_OFN1238_n_4092) );
in01f04 FE_OFC1239_n_4092 ( .a(n_4092), .o(FE_OFN1239_n_4092) );
in01f04 FE_OFC1240_n_4092 ( .a(n_4092), .o(FE_OFN1240_n_4092) );
in01f08 FE_OFC1241_n_4092 ( .a(FE_OFN1238_n_4092), .o(FE_OFN1241_n_4092) );
in01f08 FE_OFC1242_n_4092 ( .a(FE_OFN1238_n_4092), .o(FE_OFN1242_n_4092) );
in01f08 FE_OFC1243_n_4092 ( .a(FE_OFN1240_n_4092), .o(FE_OFN1243_n_4092) );
in01f08 FE_OFC1244_n_4092 ( .a(FE_OFN1239_n_4092), .o(FE_OFN1244_n_4092) );
in01f10 FE_OFC1245_n_4093 ( .a(n_4093), .o(FE_OFN1245_n_4093) );
in01f06 FE_OFC1246_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1246_n_4093) );
in01f02 FE_OFC1247_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1247_n_4093) );
in01f10 FE_OFC1248_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1248_n_4093) );
in01f08 FE_OFC1249_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1249_n_4093) );
in01f10 FE_OFC1250_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN1250_n_4093) );
in01f04 FE_OFC1251_n_4143 ( .a(n_4143), .o(FE_OFN1251_n_4143) );
in01f04 FE_OFC1252_n_4143 ( .a(FE_OFN1251_n_4143), .o(FE_OFN1252_n_4143) );
in01f08 FE_OFC1253_n_4143 ( .a(FE_OFN1251_n_4143), .o(FE_OFN1253_n_4143) );
in01f03 FE_OFC1254_n_4143 ( .a(n_4143), .o(FE_OFN1254_n_4143) );
in01f04 FE_OFC1255_n_4143 ( .a(n_4143), .o(FE_OFN1255_n_4143) );
in01f04 FE_OFC1256_n_4143 ( .a(n_4143), .o(FE_OFN1256_n_4143) );
in01f02 FE_OFC1257_n_4143 ( .a(FE_OFN1254_n_4143), .o(FE_OFN1257_n_4143) );
in01f08 FE_OFC1258_n_4143 ( .a(FE_OFN1254_n_4143), .o(FE_OFN1258_n_4143) );
in01m02 FE_OFC1259_n_4143 ( .a(FE_OFN1255_n_4143), .o(FE_OFN1259_n_4143) );
in01f08 FE_OFC1260_n_4143 ( .a(FE_OFN1255_n_4143), .o(FE_OFN1260_n_4143) );
in01f08 FE_OFC1261_n_4143 ( .a(FE_OFN1256_n_4143), .o(FE_OFN1261_n_4143) );
in01f02 FE_OFC1262_n_4095 ( .a(n_4095), .o(FE_OFN1262_n_4095) );
in01f04 FE_OFC1263_n_4095 ( .a(n_4095), .o(FE_OFN1263_n_4095) );
in01f04 FE_OFC1264_n_4095 ( .a(FE_OFN1262_n_4095), .o(FE_OFN1264_n_4095) );
in01f02 FE_OFC1265_n_4095 ( .a(FE_OFN1262_n_4095), .o(FE_OFN1265_n_4095) );
in01f06 FE_OFC1266_n_4095 ( .a(n_4095), .o(FE_OFN1266_n_4095) );
in01f02 FE_OFC1267_n_4095 ( .a(n_4095), .o(FE_OFN1267_n_4095) );
in01f08 FE_OFC1268_n_4095 ( .a(FE_OFN1263_n_4095), .o(FE_OFN1268_n_4095) );
in01f08 FE_OFC1269_n_4095 ( .a(FE_OFN1267_n_4095), .o(FE_OFN1269_n_4095) );
in01f08 FE_OFC1270_n_4095 ( .a(FE_OFN1266_n_4095), .o(FE_OFN1270_n_4095) );
in01f08 FE_OFC1271_n_4096 ( .a(n_4096), .o(FE_OFN1271_n_4096) );
in01f08 FE_OFC1272_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1272_n_4096) );
in01f02 FE_OFC1273_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1273_n_4096) );
in01f06 FE_OFC1274_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1274_n_4096) );
in01f04 FE_OFC1275_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1275_n_4096) );
in01f08 FE_OFC1276_n_4096 ( .a(FE_OFN1271_n_4096), .o(FE_OFN1276_n_4096) );
in01f06 FE_OFC1277_n_4097 ( .a(n_4097), .o(FE_OFN1277_n_4097) );
in01f08 FE_OFC1278_n_4097 ( .a(FE_OFN1277_n_4097), .o(FE_OFN1278_n_4097) );
in01f04 FE_OFC1279_n_4097 ( .a(FE_OFN1277_n_4097), .o(FE_OFN1279_n_4097) );
in01f04 FE_OFC1280_n_4097 ( .a(n_4097), .o(FE_OFN1280_n_4097) );
in01f08 FE_OFC1281_n_4097 ( .a(n_4097), .o(FE_OFN1281_n_4097) );
in01f04 FE_OFC1282_n_4097 ( .a(FE_OFN1280_n_4097), .o(FE_OFN1282_n_4097) );
in01f06 FE_OFC1283_n_4097 ( .a(FE_OFN1280_n_4097), .o(FE_OFN1283_n_4097) );
in01f08 FE_OFC1284_n_4097 ( .a(FE_OFN1281_n_4097), .o(FE_OFN1284_n_4097) );
in01f08 FE_OFC1285_n_4097 ( .a(FE_OFN1281_n_4097), .o(FE_OFN1285_n_4097) );
in01f02 FE_OFC1286_n_4098 ( .a(n_4098), .o(FE_OFN1286_n_4098) );
in01m02 FE_OFC1287_n_4098 ( .a(n_4098), .o(FE_OFN1287_n_4098) );
in01f06 FE_OFC1288_n_4098 ( .a(FE_OFN1286_n_4098), .o(FE_OFN1288_n_4098) );
in01f04 FE_OFC1289_n_4098 ( .a(FE_OFN1287_n_4098), .o(FE_OFN1289_n_4098) );
in01f04 FE_OFC1290_n_4098 ( .a(n_4098), .o(FE_OFN1290_n_4098) );
in01f04 FE_OFC1291_n_4098 ( .a(n_4098), .o(FE_OFN1291_n_4098) );
in01f04 FE_OFC1292_n_4098 ( .a(n_4098), .o(FE_OFN1292_n_4098) );
in01f08 FE_OFC1293_n_4098 ( .a(FE_OFN1290_n_4098), .o(FE_OFN1293_n_4098) );
in01f08 FE_OFC1294_n_4098 ( .a(FE_OFN1291_n_4098), .o(FE_OFN1294_n_4098) );
in01f08 FE_OFC1295_n_4098 ( .a(FE_OFN1292_n_4098), .o(FE_OFN1295_n_4098) );
in01f04 FE_OFC1296_n_5763 ( .a(n_5763), .o(FE_OFN1296_n_5763) );
in01f08 FE_OFC1297_n_5763 ( .a(n_5763), .o(FE_OFN1297_n_5763) );
in01s02 FE_OFC1298_n_5763 ( .a(n_5763), .o(FE_OFN1298_n_5763) );
in01f08 FE_OFC1299_n_5763 ( .a(FE_OFN1297_n_5763), .o(FE_OFN1299_n_5763) );
in01f04 FE_OFC1300_n_5763 ( .a(FE_OFN1298_n_5763), .o(FE_OFN1300_n_5763) );
in01f10 FE_OFC1301_n_5763 ( .a(FE_OFN1297_n_5763), .o(FE_OFN1301_n_5763) );
in01f08 FE_OFC1302_n_5763 ( .a(FE_OFN1296_n_5763), .o(FE_OFN1302_n_5763) );
in01f08 FE_OFC1303_n_13124 ( .a(n_13124), .o(FE_OFN1303_n_13124) );
in01f08 FE_OFC1304_n_13124 ( .a(FE_OFN1303_n_13124), .o(FE_OFN1304_n_13124) );
in01f08 FE_OFC1305_n_13124 ( .a(FE_OFN1303_n_13124), .o(FE_OFN1305_n_13124) );
in01m08 FE_OFC1306_n_13124 ( .a(FE_OFN1303_n_13124), .o(FE_OFN1306_n_13124) );
in01f40 FE_OFC1307_n_6624 ( .a(n_6624), .o(FE_OFN1307_n_6624) );
in01f80 FE_OFC1308_n_6624 ( .a(n_6624), .o(FE_OFN1308_n_6624) );
in01f40 FE_OFC1309_n_6624 ( .a(n_6624), .o(FE_OFN1309_n_6624) );
in01f20 FE_OFC1310_n_6624 ( .a(FE_OFN1308_n_6624), .o(FE_OFN1310_n_6624) );
in01f20 FE_OFC1311_n_6624 ( .a(FE_OFN1307_n_6624), .o(FE_OFN1311_n_6624) );
in01f20 FE_OFC1312_n_6624 ( .a(FE_OFN1307_n_6624), .o(FE_OFN1312_n_6624) );
in01f20 FE_OFC1313_n_6624 ( .a(FE_OFN1308_n_6624), .o(FE_OFN1313_n_6624) );
in01f20 FE_OFC1314_n_6624 ( .a(FE_OFN1308_n_6624), .o(FE_OFN1314_n_6624) );
in01f20 FE_OFC1315_n_6624 ( .a(FE_OFN1308_n_6624), .o(FE_OFN1315_n_6624) );
in01f20 FE_OFC1316_n_6624 ( .a(FE_OFN1309_n_6624), .o(FE_OFN1316_n_6624) );
in01f20 FE_OFC1317_n_6624 ( .a(FE_OFN1309_n_6624), .o(FE_OFN1317_n_6624) );
in01f10 FE_OFC1318_n_6436 ( .a(n_6436), .o(FE_OFN1318_n_6436) );
in01f04 FE_OFC1319_n_6436 ( .a(FE_OFN1318_n_6436), .o(FE_OFN1319_n_6436) );
in01f10 FE_OFC1320_n_6436 ( .a(FE_OFN1318_n_6436), .o(FE_OFN1320_n_6436) );
in01f20 FE_OFC1321_n_6436 ( .a(n_6436), .o(FE_OFN1321_n_6436) );
in01f10 FE_OFC1322_n_6436 ( .a(FE_OFN1321_n_6436), .o(FE_OFN1322_n_6436) );
in01f20 FE_OFC1323_n_6436 ( .a(FE_OFN1321_n_6436), .o(FE_OFN1323_n_6436) );
in01f04 FE_OFC1324_n_13547 ( .a(n_13547), .o(FE_OFN1324_n_13547) );
in01f02 FE_OFC1325_n_13547 ( .a(n_13547), .o(FE_OFN1325_n_13547) );
in01f06 FE_OFC1326_n_13547 ( .a(FE_OFN1324_n_13547), .o(FE_OFN1326_n_13547) );
in01f08 FE_OFC1327_n_13547 ( .a(FE_OFN1324_n_13547), .o(FE_OFN1327_n_13547) );
in01f04 FE_OFC1328_n_13547 ( .a(n_13547), .o(FE_OFN1328_n_13547) );
in01f01 FE_OFC1329_n_13547 ( .a(n_13547), .o(FE_OFN1329_n_13547) );
in01f06 FE_OFC1330_n_13547 ( .a(FE_OFN1325_n_13547), .o(FE_OFN1330_n_13547) );
in01f08 FE_OFC1331_n_13547 ( .a(FE_OFN1328_n_13547), .o(FE_OFN1331_n_13547) );
in01f04 FE_OFC1332_n_13547 ( .a(FE_OFN1328_n_13547), .o(FE_OFN1332_n_13547) );
in01f04 FE_OFC1333_n_13547 ( .a(FE_OFN1329_n_13547), .o(FE_OFN1333_n_13547) );
in01f02 FE_OFC1334_n_13720 ( .a(n_13720), .o(FE_OFN1334_n_13720) );
in01f02 FE_OFC1335_n_13720 ( .a(FE_OFN1334_n_13720), .o(FE_OFN1335_n_13720) );
in01f10 FE_OFC1336_n_16439 ( .a(n_16439), .o(FE_OFN1336_n_16439) );
in01f20 FE_OFC1337_n_16439 ( .a(FE_OFN1336_n_16439), .o(FE_OFN1337_n_16439) );
in01f80 FE_OFC1338_n_8567 ( .a(n_8567), .o(FE_OFN1338_n_8567) );
in01f40 FE_OFC1339_n_8567 ( .a(n_8567), .o(FE_OFN1339_n_8567) );
in01f40 FE_OFC1340_n_8567 ( .a(n_8567), .o(FE_OFN1340_n_8567) );
in01f40 FE_OFC1341_n_8567 ( .a(FE_OFN1339_n_8567), .o(FE_OFN1341_n_8567) );
in01f40 FE_OFC1342_n_8567 ( .a(FE_OFN1339_n_8567), .o(FE_OFN1342_n_8567) );
in01f40 FE_OFC1343_n_8567 ( .a(FE_OFN1340_n_8567), .o(FE_OFN1343_n_8567) );
in01f20 FE_OFC1344_n_8567 ( .a(FE_OFN1340_n_8567), .o(FE_OFN1344_n_8567) );
in01f80 FE_OFC1345_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1345_n_8567) );
in01f40 FE_OFC1346_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1346_n_8567) );
in01f40 FE_OFC1347_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1347_n_8567) );
in01f80 FE_OFC1348_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1348_n_8567) );
in01f20 FE_OFC1349_n_8567 ( .a(FE_OFN1338_n_8567), .o(FE_OFN1349_n_8567) );
in01f40 FE_OFC1350_n_8567 ( .a(FE_OFN1341_n_8567), .o(FE_OFN1350_n_8567) );
in01f40 FE_OFC1351_n_8567 ( .a(FE_OFN1342_n_8567), .o(FE_OFN1351_n_8567) );
in01f40 FE_OFC1352_n_8567 ( .a(FE_OFN1343_n_8567), .o(FE_OFN1352_n_8567) );
in01f40 FE_OFC1353_n_8567 ( .a(FE_OFN1343_n_8567), .o(FE_OFN1353_n_8567) );
in01f40 FE_OFC1354_n_8567 ( .a(FE_OFN1346_n_8567), .o(FE_OFN1354_n_8567) );
in01f40 FE_OFC1355_n_8567 ( .a(FE_OFN1347_n_8567), .o(FE_OFN1355_n_8567) );
in01f20 FE_OFC1356_n_8567 ( .a(FE_OFN1347_n_8567), .o(FE_OFN1356_n_8567) );
in01f40 FE_OFC1357_n_8567 ( .a(FE_OFN1348_n_8567), .o(FE_OFN1357_n_8567) );
in01f20 FE_OFC1358_n_8567 ( .a(FE_OFN1341_n_8567), .o(FE_OFN1358_n_8567) );
in01f10 FE_OFC1359_n_8567 ( .a(FE_OFN1345_n_8567), .o(FE_OFN1359_n_8567) );
in01f40 FE_OFC1360_n_8567 ( .a(FE_OFN1345_n_8567), .o(FE_OFN1360_n_8567) );
in01f80 FE_OFC1361_n_8567 ( .a(FE_OFN1348_n_8567), .o(FE_OFN1361_n_8567) );
in01f40 FE_OFC1362_n_8567 ( .a(FE_OFN1348_n_8567), .o(FE_OFN1362_n_8567) );
in01f20 FE_OFC1363_n_8567 ( .a(FE_OFN1342_n_8567), .o(FE_OFN1363_n_8567) );
in01f10 FE_OFC1364_n_8567 ( .a(FE_OFN1342_n_8567), .o(FE_OFN1364_n_8567) );
in01f10 FE_OFC1365_n_8567 ( .a(FE_OFN1344_n_8567), .o(FE_OFN1365_n_8567) );
in01f20 FE_OFC1366_n_8567 ( .a(FE_OFN1344_n_8567), .o(FE_OFN1366_n_8567) );
in01f40 FE_OFC1367_n_8567 ( .a(FE_OFN1345_n_8567), .o(FE_OFN1367_n_8567) );
in01f20 FE_OFC1368_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1368_n_8567) );
in01f10 FE_OFC1369_n_8567 ( .a(FE_OFN1352_n_8567), .o(FE_OFN1369_n_8567) );
in01f20 FE_OFC1370_n_8567 ( .a(FE_OFN1353_n_8567), .o(FE_OFN1370_n_8567) );
in01m20 FE_OFC1371_n_8567 ( .a(FE_OFN1345_n_8567), .o(FE_OFN1371_n_8567) );
in01f20 FE_OFC1372_n_8567 ( .a(FE_OFN1354_n_8567), .o(FE_OFN1372_n_8567) );
in01f20 FE_OFC1373_n_8567 ( .a(FE_OFN1354_n_8567), .o(FE_OFN1373_n_8567) );
in01f20 FE_OFC1374_n_8567 ( .a(FE_OFN1356_n_8567), .o(FE_OFN1374_n_8567) );
in01f20 FE_OFC1376_n_8567 ( .a(FE_OFN1357_n_8567), .o(FE_OFN1376_n_8567) );
in01f20 FE_OFC1377_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1377_n_8567) );
in01f20 FE_OFC1378_n_8567 ( .a(FE_OFN1358_n_8567), .o(FE_OFN1378_n_8567) );
in01f10 FE_OFC1379_n_8567 ( .a(FE_OFN1358_n_8567), .o(FE_OFN1379_n_8567) );
in01f10 FE_OFC1380_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1380_n_8567) );
in01f20 FE_OFC1381_n_8567 ( .a(FE_OFN1352_n_8567), .o(FE_OFN1381_n_8567) );
in01f20 FE_OFC1382_n_8567 ( .a(FE_OFN1353_n_8567), .o(FE_OFN1382_n_8567) );
in01f10 FE_OFC1383_n_8567 ( .a(FE_OFN1359_n_8567), .o(FE_OFN1383_n_8567) );
in01f20 FE_OFC1384_n_8567 ( .a(FE_OFN1360_n_8567), .o(FE_OFN1384_n_8567) );
in01f20 FE_OFC1385_n_8567 ( .a(FE_OFN1355_n_8567), .o(FE_OFN1385_n_8567) );
in01f08 FE_OFC1386_n_8567 ( .a(FE_OFN1355_n_8567), .o(FE_OFN1386_n_8567) );
in01f20 FE_OFC1387_n_8567 ( .a(FE_OFN1355_n_8567), .o(FE_OFN1387_n_8567) );
in01f20 FE_OFC1388_n_8567 ( .a(FE_OFN1355_n_8567), .o(FE_OFN1388_n_8567) );
in01f20 FE_OFC1389_n_8567 ( .a(FE_OFN1357_n_8567), .o(FE_OFN1389_n_8567) );
in01f20 FE_OFC1390_n_8567 ( .a(FE_OFN1362_n_8567), .o(FE_OFN1390_n_8567) );
in01f10 FE_OFC1391_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1391_n_8567) );
in01f20 FE_OFC1392_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1392_n_8567) );
in01f20 FE_OFC1394_n_8567 ( .a(FE_OFN1363_n_8567), .o(FE_OFN1394_n_8567) );
in01f20 FE_OFC1396_n_8567 ( .a(FE_OFN1364_n_8567), .o(FE_OFN1396_n_8567) );
in01f20 FE_OFC1397_n_8567 ( .a(FE_OFN1352_n_8567), .o(FE_OFN1397_n_8567) );
in01f20 FE_OFC1398_n_8567 ( .a(FE_OFN1352_n_8567), .o(FE_OFN1398_n_8567) );
in01f20 FE_OFC1399_n_8567 ( .a(FE_OFN1353_n_8567), .o(FE_OFN1399_n_8567) );
in01f20 FE_OFC1400_n_8567 ( .a(FE_OFN1353_n_8567), .o(FE_OFN1400_n_8567) );
in01f20 FE_OFC1401_n_8567 ( .a(FE_OFN1365_n_8567), .o(FE_OFN1401_n_8567) );
in01f20 FE_OFC1402_n_8567 ( .a(FE_OFN1366_n_8567), .o(FE_OFN1402_n_8567) );
in01f20 FE_OFC1403_n_8567 ( .a(FE_OFN1366_n_8567), .o(FE_OFN1403_n_8567) );
in01f20 FE_OFC1404_n_8567 ( .a(FE_OFN1367_n_8567), .o(FE_OFN1404_n_8567) );
in01f20 FE_OFC1405_n_8567 ( .a(FE_OFN1360_n_8567), .o(FE_OFN1405_n_8567) );
in01f20 FE_OFC1406_n_8567 ( .a(FE_OFN1357_n_8567), .o(FE_OFN1406_n_8567) );
in01f20 FE_OFC1407_n_8567 ( .a(FE_OFN1357_n_8567), .o(FE_OFN1407_n_8567) );
in01f20 FE_OFC1408_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1408_n_8567) );
in01f20 FE_OFC1409_n_8567 ( .a(FE_OFN1362_n_8567), .o(FE_OFN1409_n_8567) );
in01f20 FE_OFC1410_n_8567 ( .a(FE_OFN1362_n_8567), .o(FE_OFN1410_n_8567) );
in01f20 FE_OFC1411_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1411_n_8567) );
in01f10 FE_OFC1412_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1412_n_8567) );
in01f10 FE_OFC1413_n_8567 ( .a(FE_OFN1351_n_8567), .o(FE_OFN1413_n_8567) );
in01f20 FE_OFC1414_n_8567 ( .a(FE_OFN1367_n_8567), .o(FE_OFN1414_n_8567) );
in01f20 FE_OFC1415_n_8567 ( .a(FE_OFN1367_n_8567), .o(FE_OFN1415_n_8567) );
in01f20 FE_OFC1416_n_8567 ( .a(FE_OFN1360_n_8567), .o(FE_OFN1416_n_8567) );
in01f20 FE_OFC1417_n_8567 ( .a(FE_OFN1360_n_8567), .o(FE_OFN1417_n_8567) );
in01f20 FE_OFC1419_n_8567 ( .a(FE_OFN1371_n_8567), .o(FE_OFN1419_n_8567) );
in01f20 FE_OFC1420_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1420_n_8567) );
in01f20 FE_OFC1421_n_8567 ( .a(FE_OFN1350_n_8567), .o(FE_OFN1421_n_8567) );
in01f20 FE_OFC1422_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1422_n_8567) );
in01f20 FE_OFC1423_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1423_n_8567) );
in01f20 FE_OFC1424_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1424_n_8567) );
in01f20 FE_OFC1425_n_8567 ( .a(FE_OFN1361_n_8567), .o(FE_OFN1425_n_8567) );
in01f10 FE_OFC1426_n_8567 ( .a(FE_OFN1379_n_8567), .o(FE_OFN1426_n_8567) );
in01f08 FE_OFC1427_n_8567 ( .a(FE_OFN1426_n_8567), .o(FE_OFN1427_n_8567) );
in01f08 FE_OFC1428_n_8567 ( .a(FE_OFN1426_n_8567), .o(FE_OFN1428_n_8567) );
in01f08 FE_OFC1429_n_16779 ( .a(n_16779), .o(FE_OFN1429_n_16779) );
in01f06 FE_OFC1430_n_16779 ( .a(n_16779), .o(FE_OFN1430_n_16779) );
in01f04 FE_OFC1431_n_16779 ( .a(FE_OFN1429_n_16779), .o(FE_OFN1431_n_16779) );
in01f10 FE_OFC1432_n_16779 ( .a(FE_OFN1429_n_16779), .o(FE_OFN1432_n_16779) );
in01f08 FE_OFC1433_n_16779 ( .a(FE_OFN1430_n_16779), .o(FE_OFN1433_n_16779) );
in01f01 FE_OFC1434_n_9372 ( .a(n_9372), .o(FE_OFN1434_n_9372) );
in01f20 FE_OFC1435_n_9372 ( .a(n_9372), .o(FE_OFN1435_n_9372) );
in01f10 FE_OFC1436_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1436_n_9372) );
in01f08 FE_OFC1437_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1437_n_9372) );
in01f10 FE_OFC1438_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1438_n_9372) );
in01f08 FE_OFC1439_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1439_n_9372) );
in01f10 FE_OFC1440_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1440_n_9372) );
in01f06 FE_OFC1441_n_9372 ( .a(FE_OFN1435_n_9372), .o(FE_OFN1441_n_9372) );
in01f06 FE_OFC1442_n_11125 ( .a(n_11125), .o(FE_OFN1442_n_11125) );
in01f08 FE_OFC1443_n_11125 ( .a(n_11125), .o(FE_OFN1443_n_11125) );
in01f04 FE_OFC1444_n_11125 ( .a(FE_OFN1442_n_11125), .o(FE_OFN1444_n_11125) );
in01f10 FE_OFC1445_n_11125 ( .a(FE_OFN1443_n_11125), .o(FE_OFN1445_n_11125) );
in01f08 FE_OFC1446_n_11125 ( .a(FE_OFN1442_n_11125), .o(FE_OFN1446_n_11125) );
in01f06 FE_OFC1447_n_9163 ( .a(n_9163), .o(FE_OFN1447_n_9163) );
in01f02 FE_OFC1448_n_9163 ( .a(n_9163), .o(FE_OFN1448_n_9163) );
in01f04 FE_OFC1449_n_9163 ( .a(FE_OFN1448_n_9163), .o(FE_OFN1449_n_9163) );
in01f02 FE_OFC1450_n_9163 ( .a(FE_OFN1448_n_9163), .o(FE_OFN1450_n_9163) );
in01f08 FE_OFC1451_n_10588 ( .a(n_10588), .o(FE_OFN1451_n_10588) );
in01f04 FE_OFC1452_n_10588 ( .a(n_10588), .o(FE_OFN1452_n_10588) );
in01f08 FE_OFC1453_n_10588 ( .a(FE_OFN1452_n_10588), .o(FE_OFN1453_n_10588) );
in01f10 FE_OFC1454_n_11138 ( .a(n_11138), .o(FE_OFN1454_n_11138) );
in01f08 FE_OFC1455_n_11138 ( .a(FE_OFN1454_n_11138), .o(FE_OFN1455_n_11138) );
in01f08 FE_OFC1456_n_11138 ( .a(FE_OFN1454_n_11138), .o(FE_OFN1456_n_11138) );
in01f08 FE_OFC1457_n_11138 ( .a(FE_OFN1454_n_11138), .o(FE_OFN1457_n_11138) );
in01f08 FE_OFC1458_n_11138 ( .a(FE_OFN1454_n_11138), .o(FE_OFN1458_n_11138) );
in01f10 FE_OFC1459_n_11795 ( .a(n_11795), .o(FE_OFN1459_n_11795) );
in01f10 FE_OFC1460_n_11795 ( .a(FE_OFN1459_n_11795), .o(FE_OFN1460_n_11795) );
in01f06 FE_OFC1461_n_11795 ( .a(FE_OFN1459_n_11795), .o(FE_OFN1461_n_11795) );
in01f08 FE_OFC1462_n_11795 ( .a(FE_OFN1459_n_11795), .o(FE_OFN1462_n_11795) );
in01f08 FE_OFC1463_n_10789 ( .a(n_10789), .o(FE_OFN1463_n_10789) );
in01f08 FE_OFC1464_n_10789 ( .a(n_10789), .o(FE_OFN1464_n_10789) );
in01f08 FE_OFC1465_n_10789 ( .a(FE_OFN1463_n_10789), .o(FE_OFN1465_n_10789) );
in01f08 FE_OFC1466_n_10789 ( .a(FE_OFN1464_n_10789), .o(FE_OFN1466_n_10789) );
in01f08 FE_OFC1467_n_10789 ( .a(FE_OFN1464_n_10789), .o(FE_OFN1467_n_10789) );
in01f08 FE_OFC1468_n_10789 ( .a(FE_OFN1463_n_10789), .o(FE_OFN1468_n_10789) );
in01f08 FE_OFC1469_g52675_p ( .a(g52675_p), .o(FE_OFN1469_g52675_p) );
in01f02 FE_OFC146_g65530_p ( .a(g65530_p), .o(FE_OFN146_g65530_p) );
in01f08 FE_OFC1470_g52675_p ( .a(FE_OFN1469_g52675_p), .o(FE_OFN1470_g52675_p) );
in01f08 FE_OFC1471_g52675_p ( .a(FE_OFN1469_g52675_p), .o(FE_OFN1471_g52675_p) );
in01f06 FE_OFC1472_g52675_p ( .a(FE_OFN1469_g52675_p), .o(FE_OFN1472_g52675_p) );
in01f06 FE_OFC1473_n_16637 ( .a(n_16637), .o(FE_OFN1473_n_16637) );
in01f08 FE_OFC1474_n_16637 ( .a(n_16637), .o(FE_OFN1474_n_16637) );
in01f08 FE_OFC1475_n_16637 ( .a(n_16637), .o(FE_OFN1475_n_16637) );
in01f08 FE_OFC1477_n_16637 ( .a(FE_OFN1473_n_16637), .o(FE_OFN1477_n_16637) );
in01f08 FE_OFC1478_n_16637 ( .a(FE_OFN1474_n_16637), .o(FE_OFN1478_n_16637) );
in01f10 FE_OFC1479_n_16637 ( .a(FE_OFN1475_n_16637), .o(FE_OFN1479_n_16637) );
in01f02 FE_OFC147_g65530_p ( .a(FE_OFN146_g65530_p), .o(FE_OFN147_g65530_p) );
in01f03 FE_OFC1480_n_15534 ( .a(n_15534), .o(FE_OFN1480_n_15534) );
in01f06 FE_OFC1481_n_15534 ( .a(n_15534), .o(FE_OFN1481_n_15534) );
in01f03 FE_OFC1483_n_15534 ( .a(n_15534), .o(FE_OFN1483_n_15534) );
in01f06 FE_OFC1484_n_15534 ( .a(FE_OFN1480_n_15534), .o(FE_OFN1484_n_15534) );
in01f08 FE_OFC1485_n_15534 ( .a(FE_OFN1483_n_15534), .o(FE_OFN1485_n_15534) );
in01f10 FE_OFC1486_n_16992 ( .a(n_16992), .o(FE_OFN1486_n_16992) );
in01f08 FE_OFC1487_n_9320 ( .a(n_9320), .o(FE_OFN1487_n_9320) );
in01f02 FE_OFC1488_n_9320 ( .a(n_9320), .o(FE_OFN1488_n_9320) );
in01f08 FE_OFC1489_n_9320 ( .a(FE_OFN1487_n_9320), .o(FE_OFN1489_n_9320) );
in01f08 FE_OFC1490_n_9320 ( .a(FE_OFN1487_n_9320), .o(FE_OFN1490_n_9320) );
in01f02 FE_OFC1491_n_9320 ( .a(FE_OFN1487_n_9320), .o(FE_OFN1491_n_9320) );
in01f08 FE_OFC1492_n_9320 ( .a(FE_OFN1490_n_9320), .o(FE_OFN1492_n_9320) );
in01f08 FE_OFC1493_n_9320 ( .a(FE_OFN1492_n_9320), .o(FE_OFN1493_n_9320) );
in01f08 FE_OFC1495_n_15558 ( .a(n_15558), .o(FE_OFN1495_n_15558) );
in01f04 FE_OFC1496_n_15558 ( .a(n_15558), .o(FE_OFN1496_n_15558) );
in01f06 FE_OFC1497_n_15558 ( .a(n_15558), .o(FE_OFN1497_n_15558) );
in01f06 FE_OFC1498_n_15558 ( .a(FE_OFN1495_n_15558), .o(FE_OFN1498_n_15558) );
in01f10 FE_OFC1499_n_15558 ( .a(FE_OFN1495_n_15558), .o(FE_OFN1499_n_15558) );
in01f04 FE_OFC1500_n_15558 ( .a(FE_OFN1496_n_15558), .o(FE_OFN1500_n_15558) );
in01f04 FE_OFC1501_n_15558 ( .a(FE_OFN1496_n_15558), .o(FE_OFN1501_n_15558) );
in01f08 FE_OFC1502_n_15558 ( .a(FE_OFN1497_n_15558), .o(FE_OFN1502_n_15558) );
in01f08 FE_OFC1505_n_15768 ( .a(FE_OFN1503_n_15768), .o(FE_OFN1505_n_15768) );
in01f01 FE_OFC1506_n_15768 ( .a(FE_OFN1503_n_15768), .o(FE_OFN1506_n_15768) );
in01f08 FE_OFC1507_n_15587 ( .a(n_15587), .o(FE_OFN1507_n_15587) );
in01f08 FE_OFC1508_n_15587 ( .a(FE_OFN1507_n_15587), .o(FE_OFN1508_n_15587) );
in01f04 FE_OFC1509_n_15587 ( .a(FE_OFN1507_n_15587), .o(FE_OFN1509_n_15587) );
in01f04 FE_OFC1510_n_15587 ( .a(FE_OFN1507_n_15587), .o(FE_OFN1510_n_15587) );
in01f04 FE_OFC1511_n_15587 ( .a(FE_OFN1507_n_15587), .o(FE_OFN1511_n_15587) );
in01f04 FE_OFC1513_n_14987 ( .a(FE_OCP_RBN1923_n_10273), .o(FE_OFN1513_n_14987) );
in01f04 FE_OFC1514_n_10538 ( .a(FE_OCP_RBN1965_FE_RN_459_0), .o(FE_OFN1514_n_10538) );
in01f06 FE_OFC1519_n_10892 ( .a(n_10892), .o(FE_OFN1519_n_10892) );
in01f06 FE_OFC1520_n_10892 ( .a(n_10892), .o(FE_OFN1520_n_10892) );
in01f04 FE_OFC1521_n_10892 ( .a(FE_OFN1519_n_10892), .o(FE_OFN1521_n_10892) );
in01f08 FE_OFC1522_n_10892 ( .a(FE_OFN1519_n_10892), .o(FE_OFN1522_n_10892) );
in01f08 FE_OFC1523_n_10892 ( .a(FE_OFN1520_n_10892), .o(FE_OFN1523_n_10892) );
in01f04 FE_OFC1524_n_10853 ( .a(n_10853), .o(FE_OFN1524_n_10853) );
in01f04 FE_OFC1525_n_10853 ( .a(n_10853), .o(FE_OFN1525_n_10853) );
in01f08 FE_OFC1526_n_10853 ( .a(n_10853), .o(FE_OFN1526_n_10853) );
in01f08 FE_OFC1527_n_10853 ( .a(FE_OFN1524_n_10853), .o(FE_OFN1527_n_10853) );
in01f08 FE_OFC1528_n_10853 ( .a(FE_OFN1526_n_10853), .o(FE_OFN1528_n_10853) );
in01f08 FE_OFC1529_n_10853 ( .a(FE_OFN1525_n_10853), .o(FE_OFN1529_n_10853) );
in01f10 FE_OFC1530_n_10853 ( .a(FE_OFN1526_n_10853), .o(FE_OFN1530_n_10853) );
in01f04 FE_OFC1531_n_10143 ( .a(n_10143), .o(FE_OFN1531_n_10143) );
in01f08 FE_OFC1532_n_10143 ( .a(n_10143), .o(FE_OFN1532_n_10143) );
in01f06 FE_OFC1533_n_10143 ( .a(n_10143), .o(FE_OFN1533_n_10143) );
in01f04 FE_OFC1535_n_10143 ( .a(FE_OFN1533_n_10143), .o(FE_OFN1535_n_10143) );
in01f08 FE_OFC1536_n_10143 ( .a(FE_OFN1533_n_10143), .o(FE_OFN1536_n_10143) );
in01f02 FE_OFC1537_n_10595 ( .a(n_10595), .o(FE_OFN1537_n_10595) );
in01f02 FE_OFC1538_n_10595 ( .a(FE_OFN1537_n_10595), .o(FE_OFN1538_n_10595) );
in01f04 FE_OFC1539_n_10595 ( .a(FE_OFN1537_n_10595), .o(FE_OFN1539_n_10595) );
in01f03 FE_OFC1540_n_10595 ( .a(n_10595), .o(FE_OFN1540_n_10595) );
in01f06 FE_OFC1541_n_10595 ( .a(n_10595), .o(FE_OFN1541_n_10595) );
in01f04 FE_OFC1542_n_10566 ( .a(n_10566), .o(FE_OFN1542_n_10566) );
in01f08 FE_OFC1543_n_10566 ( .a(n_10566), .o(FE_OFN1543_n_10566) );
in01f06 FE_OFC1544_n_10566 ( .a(n_10566), .o(FE_OFN1544_n_10566) );
in01f04 FE_OFC1545_n_10566 ( .a(FE_OFN1543_n_10566), .o(FE_OFN1545_n_10566) );
in01f10 FE_OFC1546_n_10566 ( .a(FE_OFN1543_n_10566), .o(FE_OFN1546_n_10566) );
in01f08 FE_OFC1547_n_10566 ( .a(FE_OFN1542_n_10566), .o(FE_OFN1547_n_10566) );
in01f08 FE_OFC1548_n_10566 ( .a(FE_OFN1544_n_10566), .o(FE_OFN1548_n_10566) );
in01f06 FE_OFC1549_n_12104 ( .a(n_12104), .o(FE_OFN1549_n_12104) );
in01f02 FE_OFC1550_n_12104 ( .a(n_12104), .o(FE_OFN1550_n_12104) );
in01f04 FE_OFC1551_n_12104 ( .a(FE_OFN1549_n_12104), .o(FE_OFN1551_n_12104) );
in01f06 FE_OFC1552_n_12104 ( .a(FE_OFN1549_n_12104), .o(FE_OFN1552_n_12104) );
in01f06 FE_OFC1553_n_12104 ( .a(FE_OFN1550_n_12104), .o(FE_OFN1553_n_12104) );
in01f06 FE_OFC1554_n_12104 ( .a(FE_OFN1549_n_12104), .o(FE_OFN1554_n_12104) );
in01f06 FE_OFC1556_n_12042 ( .a(FE_OCP_RBN2229_n_15969), .o(FE_OFN1556_n_12042) );
in01f04 FE_OFC1558_n_12042 ( .a(FE_OCP_RBN2229_n_15969), .o(FE_OFN1558_n_12042) );
in01f10 FE_OFC1559_n_12042 ( .a(FE_OFN2203_n_12042), .o(FE_OFN1559_n_12042) );
in01f06 FE_OFC1560_n_12502 ( .a(n_12502), .o(FE_OFN1560_n_12502) );
in01f02 FE_OFC1561_n_12502 ( .a(n_12502), .o(FE_OFN1561_n_12502) );
in01f02 FE_OFC1562_n_12502 ( .a(FE_OFN1561_n_12502), .o(FE_OFN1562_n_12502) );
in01f04 FE_OFC1563_n_12502 ( .a(FE_OFN1560_n_12502), .o(FE_OFN1563_n_12502) );
in01f04 FE_OFC1564_n_12502 ( .a(FE_OFN1561_n_12502), .o(FE_OFN1564_n_12502) );
in01f06 FE_OFC1565_n_12502 ( .a(FE_OFN1560_n_12502), .o(FE_OFN1565_n_12502) );
in01f08 FE_OFC1566_n_12502 ( .a(FE_OFN1560_n_12502), .o(FE_OFN1566_n_12502) );
in01f04 FE_OFC1568_n_11027 ( .a(FE_OCP_RBN2275_n_10268), .o(FE_OFN1568_n_11027) );
in01f06 FE_OFC1572_n_11027 ( .a(FE_OCP_RBN2274_n_10268), .o(FE_OFN1572_n_11027) );
in01f04 FE_OFC1573_n_12028 ( .a(n_12028), .o(FE_OFN1573_n_12028) );
in01f02 FE_OFC1574_n_12028 ( .a(FE_OFN1573_n_12028), .o(FE_OFN1574_n_12028) );
in01f08 FE_OFC1575_n_12028 ( .a(FE_OFN1573_n_12028), .o(FE_OFN1575_n_12028) );
in01f02 FE_OFC1576_n_12028 ( .a(n_12028), .o(FE_OFN1576_n_12028) );
in01f06 FE_OFC1577_n_12028 ( .a(FE_OFN1576_n_12028), .o(FE_OFN1577_n_12028) );
in01f06 FE_OFC1579_n_12306 ( .a(FE_OCP_RBN1928_n_10259), .o(FE_OFN1579_n_12306) );
in01f06 FE_OFC1581_n_12306 ( .a(FE_OCP_RBN1928_n_10259), .o(FE_OFN1581_n_12306) );
in01f06 FE_OFC1583_n_12306 ( .a(FE_OCP_RBN1927_n_10259), .o(FE_OFN1583_n_12306) );
in01f06 FE_OFC1584_n_12306 ( .a(FE_OCP_RBN1926_n_10259), .o(FE_OFN1584_n_12306) );
in01f08 FE_OFC1585_n_13736 ( .a(n_13736), .o(FE_OFN1585_n_13736) );
in01f06 FE_OFC1586_n_13736 ( .a(FE_OFN1585_n_13736), .o(FE_OFN1586_n_13736) );
in01f08 FE_OFC1587_n_13736 ( .a(FE_OFN1585_n_13736), .o(FE_OFN1587_n_13736) );
in01f06 FE_OFC1588_n_13736 ( .a(FE_OFN1585_n_13736), .o(FE_OFN1588_n_13736) );
in01f08 FE_OFC1589_n_13736 ( .a(FE_OFN1585_n_13736), .o(FE_OFN1589_n_13736) );
in01f02 FE_OFC1590_n_13741 ( .a(n_13741), .o(FE_OFN1590_n_13741) );
in01f06 FE_OFC1591_n_13741 ( .a(n_13741), .o(FE_OFN1591_n_13741) );
in01f02 FE_OFC1592_n_13741 ( .a(n_13741), .o(FE_OFN1592_n_13741) );
in01f06 FE_OFC1593_n_13741 ( .a(FE_OFN1590_n_13741), .o(FE_OFN1593_n_13741) );
in01f06 FE_OFC1596_n_13741 ( .a(FE_OFN1592_n_13741), .o(FE_OFN1596_n_13741) );
in01f08 FE_OFC1598_n_13995 ( .a(n_13995), .o(FE_OFN1598_n_13995) );
in01f06 FE_OFC1599_n_13995 ( .a(FE_OFN1598_n_13995), .o(FE_OFN1599_n_13995) );
in01f06 FE_OFC1600_n_13995 ( .a(FE_OFN1598_n_13995), .o(FE_OFN1600_n_13995) );
in01f06 FE_OFC1601_n_13995 ( .a(FE_OFN1598_n_13995), .o(FE_OFN1601_n_13995) );
in01f06 FE_OFC1602_n_13995 ( .a(FE_OFN1598_n_13995), .o(FE_OFN1602_n_13995) );
in01f04 FE_OFC1603_n_13997 ( .a(n_13997), .o(FE_OFN1603_n_13997) );
in01f04 FE_OFC1604_n_13997 ( .a(n_13997), .o(FE_OFN1604_n_13997) );
in01f08 FE_OFC1605_n_13997 ( .a(FE_OFN1603_n_13997), .o(FE_OFN1605_n_13997) );
in01f08 FE_OFC1606_n_13997 ( .a(FE_OFN1604_n_13997), .o(FE_OFN1606_n_13997) );
in01f10 FE_OFC1607_n_2122 ( .a(n_2122), .o(FE_OFN1607_n_2122) );
in01f20 FE_OFC1608_n_2122 ( .a(n_2122), .o(FE_OFN1608_n_2122) );
in01f10 FE_OFC1609_n_2122 ( .a(FE_OFN1607_n_2122), .o(FE_OFN1609_n_2122) );
in01f10 FE_OFC1610_n_2122 ( .a(FE_OFN1607_n_2122), .o(FE_OFN1610_n_2122) );
in01f08 FE_OFC1611_n_2122 ( .a(FE_OFN1608_n_2122), .o(FE_OFN1611_n_2122) );
in01f10 FE_OFC1612_n_2122 ( .a(FE_OFN1608_n_2122), .o(FE_OFN1612_n_2122) );
in01f08 FE_OFC1613_n_1787 ( .a(n_1787), .o(FE_OFN1613_n_1787) );
in01f10 FE_OFC1614_n_1787 ( .a(n_1787), .o(FE_OFN1614_n_1787) );
in01f10 FE_OFC1615_n_1787 ( .a(n_1787), .o(FE_OFN1615_n_1787) );
in01f10 FE_OFC1616_n_1787 ( .a(n_1787), .o(FE_OFN1616_n_1787) );
in01f10 FE_OFC1617_n_1787 ( .a(FE_OFN1613_n_1787), .o(FE_OFN1617_n_1787) );
in01m02 FE_OFC1618_n_1787 ( .a(FE_OFN1614_n_1787), .o(FE_OFN1618_n_1787) );
in01f10 FE_OFC1619_n_1787 ( .a(FE_OFN1614_n_1787), .o(FE_OFN1619_n_1787) );
in01f10 FE_OFC1620_n_1787 ( .a(FE_OFN1615_n_1787), .o(FE_OFN1620_n_1787) );
in01f10 FE_OFC1621_n_1787 ( .a(FE_OFN1616_n_1787), .o(FE_OFN1621_n_1787) );
in01f20 FE_OFC1622_n_4438 ( .a(n_4438), .o(FE_OFN1622_n_4438) );
in01m06 FE_OFC1623_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN1623_n_4438) );
in01m10 FE_OFC1624_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN1624_n_4438) );
in01m06 FE_OFC1625_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN1625_n_4438) );
in01f20 FE_OFC1626_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN1626_n_4438) );
in01m08 FE_OFC1627_n_4438 ( .a(FE_OFN1626_n_4438), .o(FE_OFN1627_n_4438) );
in01m10 FE_OFC1628_n_4438 ( .a(FE_OFN1627_n_4438), .o(FE_OFN1628_n_4438) );
in01f04 FE_OFC1629_n_9531 ( .a(n_9531), .o(FE_OFN1629_n_9531) );
in01f08 FE_OFC1630_n_9531 ( .a(n_9531), .o(FE_OFN1630_n_9531) );
in01f10 FE_OFC1631_n_9531 ( .a(FE_OFN1630_n_9531), .o(FE_OFN1631_n_9531) );
in01f04 FE_OFC1632_n_9531 ( .a(FE_OFN1630_n_9531), .o(FE_OFN1632_n_9531) );
in01f10 FE_OFC1633_n_9531 ( .a(FE_OFN1631_n_9531), .o(FE_OFN1633_n_9531) );
in01f03 FE_OFC1634_n_9531 ( .a(FE_OFN1633_n_9531), .o(FE_OFN1634_n_9531) );
in01f10 FE_OFC1635_n_9531 ( .a(FE_OFN1633_n_9531), .o(FE_OFN1635_n_9531) );
in01f20 FE_OFC1636_n_4460 ( .a(n_4460), .o(FE_OFN1636_n_4460) );
in01m10 FE_OFC1637_n_4671 ( .a(n_4671), .o(FE_OFN1637_n_4671) );
in01m10 FE_OFC1638_n_4671 ( .a(n_4671), .o(FE_OFN1638_n_4671) );
in01m10 FE_OFC1639_n_4671 ( .a(n_4671), .o(FE_OFN1639_n_4671) );
in01m20 FE_OFC1640_n_4671 ( .a(FE_OFN1638_n_4671), .o(FE_OFN1640_n_4671) );
in01m08 FE_OFC1641_n_4671 ( .a(n_4671), .o(FE_OFN1641_n_4671) );
in01m20 FE_OFC1642_n_4671 ( .a(FE_OFN1637_n_4671), .o(FE_OFN1642_n_4671) );
in01m20 FE_OFC1643_n_4671 ( .a(FE_OFN1639_n_4671), .o(FE_OFN1643_n_4671) );
in01m10 FE_OFC1644_n_4671 ( .a(FE_OFN1641_n_4671), .o(FE_OFN1644_n_4671) );
in01m01 FE_OFC1645_n_4671 ( .a(FE_OFN1641_n_4671), .o(FE_OFN1645_n_4671) );
in01s02 FE_OFC1646_n_9428 ( .a(n_9428), .o(FE_OFN1646_n_9428) );
in01f20 FE_OFC1647_n_9428 ( .a(n_9428), .o(FE_OFN1647_n_9428) );
in01f20 FE_OFC1648_n_9428 ( .a(FE_OFN1647_n_9428), .o(FE_OFN1648_n_9428) );
in01m03 FE_OFC1649_n_9428 ( .a(FE_OFN1647_n_9428), .o(FE_OFN1649_n_9428) );
in01m02 FE_OFC1650_n_9428 ( .a(FE_OFN1647_n_9428), .o(FE_OFN1650_n_9428) );
in01s03 FE_OFC1651_n_9428 ( .a(FE_OFN1647_n_9428), .o(FE_OFN1651_n_9428) );
in01f04 FE_OFC1652_n_9502 ( .a(n_9502), .o(FE_OFN1652_n_9502) );
in01f06 FE_OFC1653_n_9502 ( .a(n_9502), .o(FE_OFN1653_n_9502) );
in01f06 FE_OFC1654_n_9502 ( .a(FE_OFN1653_n_9502), .o(FE_OFN1654_n_9502) );
in01f06 FE_OFC1655_n_9502 ( .a(FE_OFN1653_n_9502), .o(FE_OFN1655_n_9502) );
in01m04 FE_OFC1656_n_9502 ( .a(FE_OFN1653_n_9502), .o(FE_OFN1656_n_9502) );
in01f04 FE_OFC1657_n_9502 ( .a(FE_OFN1653_n_9502), .o(FE_OFN1657_n_9502) );
in01f08 FE_OFC1658_n_4490 ( .a(n_4490), .o(FE_OFN1658_n_4490) );
in01f01 FE_OFC1659_n_4490 ( .a(FE_OFN1658_n_4490), .o(FE_OFN1659_n_4490) );
in01m10 FE_OFC1660_n_4490 ( .a(FE_OFN1658_n_4490), .o(FE_OFN1660_n_4490) );
in01f10 FE_OFC1661_n_4490 ( .a(n_4490), .o(FE_OFN1661_n_4490) );
in01m10 FE_OFC1662_n_4490 ( .a(n_4490), .o(FE_OFN1662_n_4490) );
in01m20 FE_OFC1663_n_4490 ( .a(FE_OFN1662_n_4490), .o(FE_OFN1663_n_4490) );
in01s02 FE_OFC1664_n_9477 ( .a(n_9477), .o(FE_OFN1664_n_9477) );
in01f20 FE_OFC1665_n_9477 ( .a(n_9477), .o(FE_OFN1665_n_9477) );
in01f20 FE_OFC1666_n_9477 ( .a(FE_OFN1665_n_9477), .o(FE_OFN1666_n_9477) );
in01f01 FE_OFC1667_n_9477 ( .a(FE_OFN1665_n_9477), .o(FE_OFN1667_n_9477) );
in01f02 FE_OFC1668_n_9477 ( .a(FE_OFN1665_n_9477), .o(FE_OFN1668_n_9477) );
in01f04 FE_OFC1669_n_9477 ( .a(FE_OFN1667_n_9477), .o(FE_OFN1669_n_9477) );
in01f08 FE_OFC1670_n_9477 ( .a(FE_OFN1669_n_9477), .o(FE_OFN1670_n_9477) );
in01f02 FE_OFC1671_n_9477 ( .a(FE_OFN1669_n_9477), .o(FE_OFN1671_n_9477) );
in01m20 FE_OFC1672_n_4655 ( .a(n_4655), .o(FE_OFN1672_n_4655) );
in01f10 FE_OFC1673_n_4655 ( .a(n_4655), .o(FE_OFN1673_n_4655) );
in01f20 FE_OFC1674_n_4655 ( .a(n_4655), .o(FE_OFN1674_n_4655) );
in01m06 FE_OFC1675_n_4655 ( .a(n_4655), .o(FE_OFN1675_n_4655) );
in01f20 FE_OFC1676_n_4655 ( .a(FE_OFN1673_n_4655), .o(FE_OFN1676_n_4655) );
in01f20 FE_OFC1677_n_4655 ( .a(FE_OFN1674_n_4655), .o(FE_OFN1677_n_4655) );
in01m10 FE_OFC1678_n_4655 ( .a(FE_OFN1675_n_4655), .o(FE_OFN1678_n_4655) );
in01m04 FE_OFC1679_n_4655 ( .a(FE_OFN1672_n_4655), .o(FE_OFN1679_n_4655) );
in01m20 FE_OFC1680_n_4655 ( .a(FE_OFN1672_n_4655), .o(FE_OFN1680_n_4655) );
in01m10 FE_OFC1681_n_4669 ( .a(n_4669), .o(FE_OFN1681_n_4669) );
in01f20 FE_OFC1682_n_4669 ( .a(n_4669), .o(FE_OFN1682_n_4669) );
in01f02 FE_OFC1683_n_9528 ( .a(n_9528), .o(FE_OFN1683_n_9528) );
in01f02 FE_OFC1684_n_9528 ( .a(n_9528), .o(FE_OFN1684_n_9528) );
in01f04 FE_OFC1685_n_9528 ( .a(n_9528), .o(FE_OFN1685_n_9528) );
in01f04 FE_OFC1686_n_9528 ( .a(n_9528), .o(FE_OFN1686_n_9528) );
in01f06 FE_OFC1687_n_9528 ( .a(FE_OFN1684_n_9528), .o(FE_OFN1687_n_9528) );
in01f02 FE_OFC1688_n_9528 ( .a(FE_OFN1686_n_9528), .o(FE_OFN1688_n_9528) );
in01f06 FE_OFC1689_n_9528 ( .a(FE_OFN1686_n_9528), .o(FE_OFN1689_n_9528) );
in01f08 FE_OFC1690_n_9528 ( .a(FE_OFN1685_n_9528), .o(FE_OFN1690_n_9528) );
in01f02 FE_OFC1691_n_9528 ( .a(FE_OFN1686_n_9528), .o(FE_OFN1691_n_9528) );
in01f02 FE_OFC1692_n_9528 ( .a(FE_OFN1686_n_9528), .o(FE_OFN1692_n_9528) );
in01f06 FE_OFC1693_n_3368 ( .a(n_3368), .o(FE_OFN1693_n_3368) );
in01f08 FE_OFC1694_n_3368 ( .a(FE_OFN1693_n_3368), .o(FE_OFN1694_n_3368) );
in01f06 FE_OFC1695_n_3368 ( .a(FE_OFN1693_n_3368), .o(FE_OFN1695_n_3368) );
in01f08 FE_OFC1696_n_5751 ( .a(n_5751), .o(FE_OFN1696_n_5751) );
in01f08 FE_OFC1697_n_5751 ( .a(FE_OFN1696_n_5751), .o(FE_OFN1697_n_5751) );
in01f06 FE_OFC1698_n_5751 ( .a(FE_OFN1696_n_5751), .o(FE_OFN1698_n_5751) );
in01f08 FE_OFC1699_n_5751 ( .a(FE_OFN1696_n_5751), .o(FE_OFN1699_n_5751) );
in01f08 FE_OFC1700_n_5751 ( .a(FE_OFN1696_n_5751), .o(FE_OFN1700_n_5751) );
in01f04 FE_OFC1701_n_4868 ( .a(n_4868), .o(FE_OFN1701_n_4868) );
in01f08 FE_OFC1702_n_4868 ( .a(n_4868), .o(FE_OFN1702_n_4868) );
in01f08 FE_OFC1703_n_4868 ( .a(n_4868), .o(FE_OFN1703_n_4868) );
in01f06 FE_OFC1704_n_4868 ( .a(n_4868), .o(FE_OFN1704_n_4868) );
in01f08 FE_OFC1705_n_4868 ( .a(FE_OFN1701_n_4868), .o(FE_OFN1705_n_4868) );
in01f08 FE_OFC1706_n_4868 ( .a(FE_OFN1703_n_4868), .o(FE_OFN1706_n_4868) );
in01f08 FE_OFC1707_n_4868 ( .a(FE_OFN1703_n_4868), .o(FE_OFN1707_n_4868) );
in01f08 FE_OFC1708_n_4868 ( .a(FE_OFN1704_n_4868), .o(FE_OFN1708_n_4868) );
in01f10 FE_OFC1709_n_4868 ( .a(FE_OFN1702_n_4868), .o(FE_OFN1709_n_4868) );
in01f10 FE_OFC1710_n_4868 ( .a(FE_OFN1702_n_4868), .o(FE_OFN1710_n_4868) );
in01f02 FE_OFC1711_n_13563 ( .a(n_13563), .o(FE_OFN1711_n_13563) );
in01f02 FE_OFC1712_n_13563 ( .a(FE_OFN1711_n_13563), .o(FE_OFN1712_n_13563) );
in01f02 FE_OFC1713_n_13650 ( .a(n_13650), .o(FE_OFN1713_n_13650) );
in01f02 FE_OFC1714_n_13650 ( .a(FE_OFN1713_n_13650), .o(FE_OFN1714_n_13650) );
in01f02 FE_OFC1716_n_16698 ( .a(FE_OCP_RBN2007_n_16698), .o(FE_OFN1716_n_16698) );
in01f06 FE_OFC1719_n_16891 ( .a(n_16891), .o(FE_OFN1719_n_16891) );
in01f10 FE_OFC1720_n_16891 ( .a(FE_OFN1719_n_16891), .o(FE_OFN1720_n_16891) );
in01f04 FE_OFC1721_n_16891 ( .a(n_16891), .o(FE_OFN1721_n_16891) );
in01f04 FE_OFC1722_n_16891 ( .a(n_16891), .o(FE_OFN1722_n_16891) );
in01f04 FE_OFC1723_n_16891 ( .a(FE_OFN1719_n_16891), .o(FE_OFN1723_n_16891) );
in01f08 FE_OFC1724_n_16891 ( .a(FE_OFN1722_n_16891), .o(FE_OFN1724_n_16891) );
in01f08 FE_OFC1725_n_16891 ( .a(FE_OFN1721_n_16891), .o(FE_OFN1725_n_16891) );
in01f08 FE_OFC1726_n_9975 ( .a(n_9975), .o(FE_OFN1726_n_9975) );
in01f10 FE_OFC1727_n_9975 ( .a(FE_OFN1726_n_9975), .o(FE_OFN1727_n_9975) );
in01f04 FE_OFC1728_n_9975 ( .a(FE_OFN1726_n_9975), .o(FE_OFN1728_n_9975) );
in01f06 FE_OFC1729_n_9975 ( .a(n_9975), .o(FE_OFN1729_n_9975) );
in01f06 FE_OFC1730_n_9975 ( .a(FE_OFN1729_n_9975), .o(FE_OFN1730_n_9975) );
in01f08 FE_OFC1731_n_9975 ( .a(FE_OFN1729_n_9975), .o(FE_OFN1731_n_9975) );
in01f06 FE_OFC1732_n_16317 ( .a(n_16317), .o(FE_OFN1732_n_16317) );
in01f04 FE_OFC1733_n_16317 ( .a(FE_OFN1732_n_16317), .o(FE_OFN1733_n_16317) );
in01f06 FE_OFC1734_n_16317 ( .a(FE_OFN1732_n_16317), .o(FE_OFN1734_n_16317) );
in01f06 FE_OFC1735_n_16317 ( .a(FE_OFN1732_n_16317), .o(FE_OFN1735_n_16317) );
in01f04 FE_OFC1736_n_16317 ( .a(FE_OFN1732_n_16317), .o(FE_OFN1736_n_16317) );
in01f08 FE_OFC1737_n_11019 ( .a(n_11019), .o(FE_OFN1737_n_11019) );
in01f04 FE_OFC1738_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1738_n_11019) );
in01f08 FE_OFC1739_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1739_n_11019) );
in01f02 FE_OFC1740_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1740_n_11019) );
in01f06 FE_OFC1741_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1741_n_11019) );
in01f04 FE_OFC1742_n_11019 ( .a(FE_OFN1737_n_11019), .o(FE_OFN1742_n_11019) );
in01f02 FE_OFC1743_n_12004 ( .a(n_12004), .o(FE_OFN1743_n_12004) );
in01f02 FE_OFC1744_n_12004 ( .a(n_12004), .o(FE_OFN1744_n_12004) );
in01f08 FE_OFC1745_n_12004 ( .a(n_12004), .o(FE_OFN1745_n_12004) );
in01f04 FE_OFC1746_n_12004 ( .a(FE_OFN1744_n_12004), .o(FE_OFN1746_n_12004) );
in01f04 FE_OFC1747_n_12004 ( .a(FE_OFN1743_n_12004), .o(FE_OFN1747_n_12004) );
in01f06 FE_OFC1748_n_12004 ( .a(FE_OFN1745_n_12004), .o(FE_OFN1748_n_12004) );
in01f10 FE_OFC1749_n_12004 ( .a(FE_OFN1745_n_12004), .o(FE_OFN1749_n_12004) );
in01f02 FE_OFC1751_n_12086 ( .a(FE_OCP_RBN1972_n_11767), .o(FE_OFN1751_n_12086) );
in01f06 FE_OFC1752_n_12086 ( .a(FE_OCP_RBN1972_n_11767), .o(FE_OFN1752_n_12086) );
in01f08 FE_OFC1753_n_12086 ( .a(FE_OCP_RBN1971_n_11767), .o(FE_OFN1753_n_12086) );
in01f08 FE_OFC1754_n_12681 ( .a(n_12681), .o(FE_OFN1754_n_12681) );
in01f02 FE_OFC1755_n_12681 ( .a(FE_OFN1754_n_12681), .o(FE_OFN1755_n_12681) );
in01f04 FE_OFC1756_n_12681 ( .a(FE_OFN1754_n_12681), .o(FE_OFN1756_n_12681) );
in01f08 FE_OFC1757_n_12681 ( .a(FE_OFN1754_n_12681), .o(FE_OFN1757_n_12681) );
in01f06 FE_OFC1758_n_10780 ( .a(n_10780), .o(FE_OFN1758_n_10780) );
in01f06 FE_OFC1759_n_10780 ( .a(FE_OFN1758_n_10780), .o(FE_OFN1759_n_10780) );
in01f06 FE_OFC1760_n_10780 ( .a(FE_OFN1758_n_10780), .o(FE_OFN1760_n_10780) );
in01f06 FE_OFC1761_n_10780 ( .a(FE_OFN1758_n_10780), .o(FE_OFN1761_n_10780) );
in01f06 FE_OFC1762_n_10780 ( .a(FE_OFN1758_n_10780), .o(FE_OFN1762_n_10780) );
in01f08 FE_OFC1767_n_14054 ( .a(n_14054), .o(FE_OFN1767_n_14054) );
in01f06 FE_OFC1768_n_14054 ( .a(FE_OFN1767_n_14054), .o(FE_OFN1768_n_14054) );
in01f06 FE_OFC1769_n_14054 ( .a(FE_OFN1767_n_14054), .o(FE_OFN1769_n_14054) );
in01f06 FE_OFC1770_n_14054 ( .a(FE_OFN1767_n_14054), .o(FE_OFN1770_n_14054) );
in01f06 FE_OFC1771_n_14054 ( .a(FE_OFN1767_n_14054), .o(FE_OFN1771_n_14054) );
in01f04 FE_OFC1773_n_13800 ( .a(FE_OFN1772_n_13800), .o(FE_OFN1773_n_13800) );
in01f08 FE_OFC1775_n_13800 ( .a(FE_OFN1772_n_13800), .o(FE_OFN1775_n_13800) );
in01f80 FE_OFC1776_parchk_pci_ad_reg_in_1222 ( .a(parchk_pci_ad_reg_in_1222), .o(FE_OFN1776_parchk_pci_ad_reg_in_1222) );
in01f40 FE_OFC1777_parchk_pci_ad_reg_in_1222 ( .a(FE_OFN1776_parchk_pci_ad_reg_in_1222), .o(FE_OFN1777_parchk_pci_ad_reg_in_1222) );
in01f20 FE_OFC1778_parchk_pci_ad_reg_in_1222 ( .a(FE_OFN1776_parchk_pci_ad_reg_in_1222), .o(FE_OFN1778_parchk_pci_ad_reg_in_1222) );
in01f40 FE_OFC1779_parchk_pci_ad_reg_in_1221 ( .a(parchk_pci_ad_reg_in_1221), .o(FE_OFN1779_parchk_pci_ad_reg_in_1221) );
in01f20 FE_OFC1780_parchk_pci_ad_reg_in_1221 ( .a(FE_OFN1779_parchk_pci_ad_reg_in_1221), .o(FE_OFN1780_parchk_pci_ad_reg_in_1221) );
in01f20 FE_OFC1781_parchk_pci_ad_reg_in_1221 ( .a(FE_OFN1779_parchk_pci_ad_reg_in_1221), .o(FE_OFN1781_parchk_pci_ad_reg_in_1221) );
in01f06 FE_OFC1782_n_1699 ( .a(n_1699), .o(FE_OFN1782_n_1699) );
in01f08 FE_OFC1783_n_1699 ( .a(FE_OFN1782_n_1699), .o(FE_OFN1783_n_1699) );
in01f02 FE_OFC1784_n_1699 ( .a(FE_OFN1782_n_1699), .o(FE_OFN1784_n_1699) );
in01f02 FE_OFC1785_n_1699 ( .a(FE_OFN1782_n_1699), .o(FE_OFN1785_n_1699) );
in01m04 FE_OFC1786_n_1699 ( .a(FE_OFN1782_n_1699), .o(FE_OFN1786_n_1699) );
in01f01 FE_OFC1789_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN1789_n_9823) );
in01f08 FE_OFC1790_n_2687 ( .a(n_2687), .o(FE_OFN1790_n_2687) );
in01f10 FE_OFC1791_n_9904 ( .a(FE_OFN607_n_9904), .o(FE_OFN1791_n_9904) );
in01m01 FE_OFC1792_n_9904 ( .a(FE_OFN607_n_9904), .o(FE_OFN1792_n_9904) );
in01f01 FE_OFC1793_n_9904 ( .a(FE_OFN1791_n_9904), .o(FE_OFN1793_n_9904) );
in01f10 FE_OFC1794_n_9904 ( .a(FE_OFN1791_n_9904), .o(FE_OFN1794_n_9904) );
in01s04 FE_OFC1795_n_9904 ( .a(FE_OFN1792_n_9904), .o(FE_OFN1795_n_9904) );
in01f08 FE_OFC1796_n_2299 ( .a(FE_OFN958_n_2299), .o(FE_OFN1796_n_2299) );
in01f10 FE_OFC1797_n_2299 ( .a(FE_OFN1796_n_2299), .o(FE_OFN1797_n_2299) );
in01s06 FE_OFC1798_n_9690 ( .a(FE_OFN541_n_9690), .o(FE_OFN1798_n_9690) );
in01f10 FE_OFC1799_n_9690 ( .a(FE_OFN541_n_9690), .o(FE_OFN1799_n_9690) );
in01s01 FE_OFC1800_n_9690 ( .a(FE_OFN1798_n_9690), .o(FE_OFN1800_n_9690) );
in01s04 FE_OFC1801_n_9690 ( .a(FE_OFN1798_n_9690), .o(FE_OFN1801_n_9690) );
in01s01 FE_OFC1802_n_9690 ( .a(FE_OFN1799_n_9690), .o(FE_OFN1802_n_9690) );
in01f10 FE_OFC1803_n_9690 ( .a(FE_OFN1799_n_9690), .o(FE_OFN1803_n_9690) );
in01m04 FE_OFC1804_n_4501 ( .a(FE_OFN613_n_4501), .o(FE_OFN1804_n_4501) );
in01m10 FE_OFC1805_n_4501 ( .a(FE_OFN613_n_4501), .o(FE_OFN1805_n_4501) );
in01m08 FE_OFC1806_n_4501 ( .a(FE_OFN1804_n_4501), .o(FE_OFN1806_n_4501) );
in01f10 FE_OFC1807_n_4501 ( .a(FE_OFN1805_n_4501), .o(FE_OFN1807_n_4501) );
in01f10 FE_OFC1808_n_4454 ( .a(FE_OFN632_n_4454), .o(FE_OFN1808_n_4454) );
in01f02 FE_OFC1809_n_4454 ( .a(FE_OFN1808_n_4454), .o(FE_OFN1809_n_4454) );
in01f10 FE_OFC1810_n_4454 ( .a(FE_OFN1808_n_4454), .o(FE_OFN1810_n_4454) );
in01f08 FE_OFC1811_n_7845 ( .a(FE_OFN700_n_7845), .o(FE_OFN1811_n_7845) );
in01f10 FE_OFC1812_n_7845 ( .a(FE_OFN1811_n_7845), .o(FE_OFN1812_n_7845) );
in01f02 FE_OFC1813_n_2919 ( .a(FE_OFN1819_n_2919), .o(FE_OFN1813_n_2919) );
in01f01 FE_OFC1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(FE_OFN1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid) );
in01m04 FE_OFC1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid ( .a(FE_OFN1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid) );
in01f02 FE_OFC1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid ( .a(FE_OFN1814_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid) );
in01f02 FE_OFC1819_n_2919 ( .a(n_2919), .o(FE_OFN1819_n_2919) );
in01f01 FE_OFC186_n_15768 ( .a(FE_OFN1503_n_15768), .o(FE_OFN186_n_15768) );
in01f20 FE_OFC190_n_1193 ( .a(n_1193), .o(FE_OFN190_n_1193) );
in01f20 FE_OFC191_n_1193 ( .a(FE_OFN190_n_1193), .o(FE_OFN191_n_1193) );
in01f02 FE_OFC1935_n_1781 ( .a(n_1781), .o(FE_OFN1935_n_1781) );
in01f02 FE_OFC1936_n_1781 ( .a(FE_OFN1935_n_1781), .o(FE_OFN1936_n_1781) );
in01m02 FE_OFC1937_g66085_p ( .a(g66085_p), .o(FE_OFN1937_g66085_p) );
in01f06 FE_OFC1938_g66085_p ( .a(FE_OFN1937_g66085_p), .o(FE_OFN1938_g66085_p) );
in01m02 FE_OFC1939_g66095_p ( .a(g66095_p), .o(FE_OFN1939_g66095_p) );
in01f04 FE_OFC1940_g66095_p ( .a(FE_OFN1939_g66095_p), .o(FE_OFN1940_g66095_p) );
in01f02 FE_OFC1941_n_3241 ( .a(n_3241), .o(FE_OFN1941_n_3241) );
in01f02 FE_OFC1942_n_3241 ( .a(FE_OFN1941_n_3241), .o(FE_OFN1942_n_3241) );
in01f02 FE_OFC1943_n_15813 ( .a(n_15813), .o(FE_OFN1943_n_15813) );
in01f02 FE_OFC1944_n_15813 ( .a(FE_OFN1943_n_15813), .o(FE_OFN1944_n_15813) );
in01f40 FE_OFC1945_n_13784 ( .a(n_13784), .o(FE_OFN1945_n_13784) );
in01f40 FE_OFC1946_n_13784 ( .a(FE_OFN1945_n_13784), .o(FE_OFN1946_n_13784) );
in01f04 FE_OFC196_n_2683 ( .a(n_2683), .o(FE_OFN196_n_2683) );
in01f06 FE_OFC197_n_2683 ( .a(FE_OFN196_n_2683), .o(FE_OFN197_n_2683) );
in01f02 FE_OFC198_n_3298 ( .a(n_3298), .o(FE_OFN198_n_3298) );
in01f02 FE_OFC199_n_3298 ( .a(FE_OFN198_n_3298), .o(FE_OFN199_n_3298) );
in01f08 FE_OFC1_n_4778 ( .a(FE_OFN1079_n_4778), .o(FE_OFN1_n_4778) );
in01m02 FE_OFC200_n_9230 ( .a(n_9230), .o(FE_OFN200_n_9230) );
in01s06 FE_OFC201_n_9230 ( .a(FE_OFN200_n_9230), .o(FE_OFN201_n_9230) );
in01f01 FE_OFC2020_n_4778 ( .a(FE_OFN1079_n_4778), .o(FE_OFN2020_n_4778) );
in01m04 FE_OFC2021_n_4778 ( .a(FE_OFN2020_n_4778), .o(FE_OFN2021_n_4778) );
in01f03 FE_OFC2022_n_4778 ( .a(FE_OFN2020_n_4778), .o(FE_OFN2022_n_4778) );
in01s02 FE_OFC202_n_9228 ( .a(n_9228), .o(FE_OFN202_n_9228) );
in01s04 FE_OFC203_n_9228 ( .a(FE_OFN202_n_9228), .o(FE_OFN203_n_9228) );
in01f02 FE_OFC204_n_9140 ( .a(n_9140), .o(FE_OFN204_n_9140) );
in01f04 FE_OFC2051_n_6965 ( .a(n_6965), .o(FE_OFN2051_n_6965) );
in01f06 FE_OFC2052_n_6965 ( .a(FE_OFN2051_n_6965), .o(FE_OFN2052_n_6965) );
in01f80 FE_OFC2053_n_8831 ( .a(n_8831), .o(FE_OFN2053_n_8831) );
in01f80 FE_OFC2054_n_8831 ( .a(FE_OFN2053_n_8831), .o(FE_OFN2054_n_8831) );
in01f80 FE_OFC2055_n_8831 ( .a(FE_OFN2053_n_8831), .o(FE_OFN2055_n_8831) );
in01f02 FE_OFC2056_n_2117 ( .a(n_2117), .o(FE_OFN2056_n_2117) );
in01f04 FE_OFC2057_n_2117 ( .a(FE_OFN2056_n_2117), .o(FE_OFN2057_n_2117) );
in01f10 FE_OFC2058_n_13447 ( .a(n_13447), .o(FE_OFN2058_n_13447) );
in01f20 FE_OFC2059_n_13447 ( .a(FE_OFN2058_n_13447), .o(FE_OFN2059_n_13447) );
in01f06 FE_OFC205_n_9140 ( .a(FE_OFN204_n_9140), .o(FE_OFN205_n_9140) );
in01m02 FE_OFC2060_g66087_p ( .a(g66087_p), .o(FE_OFN2060_g66087_p) );
in01m06 FE_OFC2061_g66087_p ( .a(FE_OFN2060_g66087_p), .o(FE_OFN2061_g66087_p) );
in01f20 FE_OFC2062_n_6391 ( .a(FE_OFN1223_n_6391), .o(FE_OFN2062_n_6391) );
in01f10 FE_OFC2063_n_6391 ( .a(FE_OFN2062_n_6391), .o(FE_OFN2063_n_6391) );
in01f10 FE_OFC2064_n_6391 ( .a(FE_OFN2062_n_6391), .o(FE_OFN2064_n_6391) );
in01f10 FE_OFC2069_n_15978 ( .a(FE_OFN1000_n_15978), .o(FE_OFN2069_n_15978) );
in01m04 FE_OFC206_n_9865 ( .a(n_9865), .o(FE_OFN206_n_9865) );
in01f08 FE_OFC2070_n_15978 ( .a(FE_OFN2069_n_15978), .o(FE_OFN2070_n_15978) );
in01f08 FE_OFC2071_n_15978 ( .a(FE_OFN1001_n_15978), .o(FE_OFN2071_n_15978) );
in01f10 FE_OFC2072_n_15978 ( .a(FE_OFN2071_n_15978), .o(FE_OFN2072_n_15978) );
in01f02 FE_OFC2073_n_2723 ( .a(n_2723), .o(FE_OFN2073_n_2723) );
in01f04 FE_OFC2074_n_2723 ( .a(FE_OFN2073_n_2723), .o(FE_OFN2074_n_2723) );
in01f10 FE_OFC2075_FE_OCPUNCON1952_FE_OFN697_n_16760 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(FE_OFN2075_FE_OCPUNCON1952_FE_OFN697_n_16760) );
in01f20 FE_OFC2076_FE_OCPUNCON1952_FE_OFN697_n_16760 ( .a(FE_OFN2075_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760) );
in01f40 FE_OFC2077_n_8069 ( .a(n_8069), .o(FE_OFN2077_n_8069) );
in01f20 FE_OFC2079_n_8069 ( .a(FE_OFN2077_n_8069), .o(FE_OFN2079_n_8069) );
in01m08 FE_OFC207_n_9865 ( .a(FE_OFN206_n_9865), .o(FE_OFN207_n_9865) );
in01f02 FE_OFC2080_n_8176 ( .a(n_8176), .o(FE_OFN2080_n_8176) );
in01f08 FE_OFC2081_n_8176 ( .a(FE_OFN2080_n_8176), .o(FE_OFN2081_n_8176) );
in01f06 FE_OFC2082_n_8407 ( .a(n_8407), .o(FE_OFN2082_n_8407) );
in01f06 FE_OFC2083_n_8407 ( .a(FE_OFN2082_n_8407), .o(FE_OFN2083_n_8407) );
in01f03 FE_OFC2084_n_8407 ( .a(FE_OFN2082_n_8407), .o(FE_OFN2084_n_8407) );
in01f02 FE_OFC2085_n_8448 ( .a(n_8448), .o(FE_OFN2085_n_8448) );
in01f02 FE_OFC2086_n_8448 ( .a(FE_OFN2085_n_8448), .o(FE_OFN2086_n_8448) );
in01f02 FE_OFC2088_n_13124 ( .a(FE_OFN2132_n_13124), .o(FE_OFN2088_n_13124) );
in01m02 FE_OFC208_n_9126 ( .a(n_9126), .o(FE_OFN208_n_9126) );
in01f20 FE_OFC2092_n_2301 ( .a(n_2301), .o(FE_OFN2092_n_2301) );
in01f20 FE_OFC2093_n_2301 ( .a(FE_OFN2092_n_2301), .o(FE_OFN2093_n_2301) );
in01f04 FE_OFC2094_n_2520 ( .a(n_2520), .o(FE_OFN2094_n_2520) );
in01m06 FE_OFC2095_n_2520 ( .a(FE_OFN2094_n_2520), .o(FE_OFN2095_n_2520) );
in01m04 FE_OFC2096_n_2520 ( .a(FE_OFN2094_n_2520), .o(FE_OFN2096_n_2520) );
in01f02 FE_OFC2099_n_3281 ( .a(n_3281), .o(FE_OFN2099_n_3281) );
in01m06 FE_OFC209_n_9126 ( .a(FE_OFN208_n_9126), .o(FE_OFN209_n_9126) );
in01f04 FE_OFC2100_n_3281 ( .a(FE_OFN2099_n_3281), .o(FE_OFN2100_n_3281) );
in01f02 FE_OFC2101_n_2834 ( .a(n_2834), .o(FE_OFN2101_n_2834) );
in01f02 FE_OFC2102_n_2834 ( .a(FE_OFN2101_n_2834), .o(FE_OFN2102_n_2834) );
in01f10 FE_OFC2103_g64577_p ( .a(FE_OFN1106_g64577_p), .o(FE_OFN2103_g64577_p) );
in01f08 FE_OFC2104_g64577_p ( .a(FE_OFN2103_g64577_p), .o(FE_OFN2104_g64577_p) );
in01f10 FE_OFC2105_g64577_p ( .a(FE_OFN2103_g64577_p), .o(FE_OFN2105_g64577_p) );
in01f10 FE_OFC2106_g64577_p ( .a(FE_OFN2103_g64577_p), .o(FE_OFN2106_g64577_p) );
in01f10 FE_OFC2107_n_2047 ( .a(FE_OFN1003_n_2047), .o(FE_OFN2107_n_2047) );
in01f10 FE_OFC2108_n_2047 ( .a(FE_OFN2107_n_2047), .o(FE_OFN2108_n_2047) );
in01f08 FE_OFC2109_n_2047 ( .a(FE_OFN2107_n_2047), .o(FE_OFN2109_n_2047) );
in01f10 FE_OFC210_n_9858 ( .a(n_9858), .o(FE_OFN210_n_9858) );
in01f06 FE_OFC2110_n_2248 ( .a(FE_OFN945_n_2248), .o(FE_OFN2110_n_2248) );
in01f08 FE_OFC2111_n_2248 ( .a(FE_OFN2110_n_2248), .o(FE_OFN2111_n_2248) );
in01m10 FE_OFC2112_n_2053 ( .a(FE_OFN1016_n_2053), .o(FE_OFN2112_n_2053) );
in01m10 FE_OFC2113_n_2053 ( .a(FE_OFN2112_n_2053), .o(FE_OFN2113_n_2053) );
in01f08 FE_OFC2114_wishbone_slave_unit_pci_initiator_if_data_source ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source) );
in01m03 FE_OFC2115_wishbone_slave_unit_pci_initiator_if_data_source ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source) );
in01m10 FE_OFC2116_wishbone_slave_unit_pci_initiator_if_data_source ( .a(FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source) );
in01m06 FE_OFC2118_wishbone_slave_unit_pci_initiator_if_data_source ( .a(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source) );
in01s02 FE_OFC2119_wishbone_slave_unit_pci_initiator_if_data_source ( .a(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source) );
in01f10 FE_OFC211_n_9858 ( .a(FE_OFN210_n_9858), .o(FE_OFN211_n_9858) );
in01f10 FE_OFC2121_n_2687 ( .a(FE_OFN1790_n_2687), .o(FE_OFN2121_n_2687) );
in01f08 FE_OFC2123_n_16497 ( .a(n_16497), .o(FE_OFN2123_n_16497) );
in01f08 FE_OFC2124_n_16497 ( .a(n_16497), .o(FE_OFN2124_n_16497) );
in01f08 FE_OFC2125_n_16497 ( .a(FE_OFN2124_n_16497), .o(FE_OFN2125_n_16497) );
in01f08 FE_OFC2126_n_16497 ( .a(FE_OFN2123_n_16497), .o(FE_OFN2126_n_16497) );
in01f08 FE_OFC2127_n_16497 ( .a(FE_OFN2124_n_16497), .o(FE_OFN2127_n_16497) );
in01f10 FE_OFC2128_n_16497 ( .a(FE_OFN2123_n_16497), .o(FE_OFN2128_n_16497) );
in01f08 FE_OFC2129_n_16720 ( .a(FE_OFN1060_n_16720), .o(FE_OFN2129_n_16720) );
in01s02 FE_OFC212_n_9124 ( .a(n_9124), .o(FE_OFN212_n_9124) );
in01f08 FE_OFC2130_n_10588 ( .a(FE_OFN1451_n_10588), .o(FE_OFN2130_n_10588) );
in01f08 FE_OFC2131_n_10588 ( .a(FE_OFN1451_n_10588), .o(FE_OFN2131_n_10588) );
in01f01 FE_OFC2132_n_13124 ( .a(FE_OFN1304_n_13124), .o(FE_OFN2132_n_13124) );
in01f10 FE_OFC2133_n_13124 ( .a(FE_OFN1304_n_13124), .o(FE_OFN2133_n_13124) );
in01f10 FE_OFC2134_n_13124 ( .a(FE_OFN2133_n_13124), .o(FE_OFN2134_n_13124) );
in01f08 FE_OFC2135_n_13124 ( .a(FE_OFN2133_n_13124), .o(FE_OFN2135_n_13124) );
in01f08 FE_OFC2136_n_13124 ( .a(FE_OFN2133_n_13124), .o(FE_OFN2136_n_13124) );
in01f10 FE_OFC2137_n_15534 ( .a(FE_OFN1481_n_15534), .o(FE_OFN2137_n_15534) );
in01f08 FE_OFC2139_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2139_n_16992) );
in01s04 FE_OFC213_n_9124 ( .a(FE_OFN212_n_9124), .o(FE_OFN213_n_9124) );
in01f01 FE_OFC2140_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2140_n_16992) );
in01f01 FE_OFC2141_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2141_n_16992) );
in01f10 FE_OFC2142_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2142_n_16992) );
in01f01 FE_OFC2143_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2143_n_16992) );
in01f01 FE_OFC2144_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2144_n_16992) );
in01f01 FE_OFC2145_n_16992 ( .a(FE_OFN1486_n_16992), .o(FE_OFN2145_n_16992) );
in01f06 FE_OFC2146_n_9320 ( .a(FE_OFN1488_n_9320), .o(FE_OFN2146_n_9320) );
in01f08 FE_OFC2147_n_10595 ( .a(FE_OFN1540_n_10595), .o(FE_OFN2147_n_10595) );
in01f01 FE_OFC2148_n_10595 ( .a(FE_OFN1540_n_10595), .o(FE_OFN2148_n_10595) );
in01f08 FE_OFC2149_n_10595 ( .a(FE_OFN1541_n_10595), .o(FE_OFN2149_n_10595) );
in01s02 FE_OFC214_n_9856 ( .a(n_9856), .o(FE_OFN214_n_9856) );
in01f08 FE_OFC2150_n_10595 ( .a(FE_OFN1541_n_10595), .o(FE_OFN2150_n_10595) );
in01f20 FE_OFC2151_n_16439 ( .a(FE_OFN1337_n_16439), .o(FE_OFN2151_n_16439) );
in01f06 FE_OFC2152_n_16439 ( .a(FE_OFN1337_n_16439), .o(FE_OFN2152_n_16439) );
in01f20 FE_OFC2153_n_16439 ( .a(FE_OFN2151_n_16439), .o(FE_OFN2153_n_16439) );
in01f10 FE_OFC2154_n_16439 ( .a(FE_OFN1337_n_16439), .o(FE_OFN2154_n_16439) );
in01f10 FE_OFC2155_n_16439 ( .a(FE_OFN2151_n_16439), .o(FE_OFN2155_n_16439) );
in01f08 FE_OFC2156_n_16439 ( .a(FE_OFN2152_n_16439), .o(FE_OFN2156_n_16439) );
in01f10 FE_OFC2157_n_16439 ( .a(FE_OFN2154_n_16439), .o(FE_OFN2157_n_16439) );
in01f10 FE_OFC2158_n_16439 ( .a(FE_OFN2154_n_16439), .o(FE_OFN2158_n_16439) );
in01f10 FE_OFC2159_n_16301 ( .a(n_16301), .o(FE_OFN2159_n_16301) );
in01s06 FE_OFC215_n_9856 ( .a(FE_OFN214_n_9856), .o(FE_OFN215_n_9856) );
in01f08 FE_OFC2160_n_16301 ( .a(n_16301), .o(FE_OFN2160_n_16301) );
in01f04 FE_OFC2161_n_16301 ( .a(n_16301), .o(FE_OFN2161_n_16301) );
in01f10 FE_OFC2162_n_16301 ( .a(FE_OFN2159_n_16301), .o(FE_OFN2162_n_16301) );
in01f08 FE_OFC2163_n_16301 ( .a(FE_OFN2161_n_16301), .o(FE_OFN2163_n_16301) );
in01f10 FE_OFC2164_n_16301 ( .a(FE_OFN2159_n_16301), .o(FE_OFN2164_n_16301) );
in01f10 FE_OFC2165_n_16301 ( .a(FE_OFN2160_n_16301), .o(FE_OFN2165_n_16301) );
in01f20 FE_OFC2166_n_8567 ( .a(FE_OFN1372_n_8567), .o(FE_OFN2166_n_8567) );
in01f10 FE_OFC2167_n_8567 ( .a(FE_OFN2166_n_8567), .o(FE_OFN2167_n_8567) );
in01f10 FE_OFC2168_n_8567 ( .a(FE_OFN2166_n_8567), .o(FE_OFN2168_n_8567) );
in01f10 FE_OFC2169_n_8567 ( .a(FE_OFN2166_n_8567), .o(FE_OFN2169_n_8567) );
in01s02 FE_OFC216_n_9889 ( .a(n_9889), .o(FE_OFN216_n_9889) );
in01f10 FE_OFC2170_n_8567 ( .a(FE_OFN2166_n_8567), .o(FE_OFN2170_n_8567) );
in01f20 FE_OFC2171_n_8567 ( .a(FE_OFN1373_n_8567), .o(FE_OFN2171_n_8567) );
in01f10 FE_OFC2172_n_8567 ( .a(FE_OFN1373_n_8567), .o(FE_OFN2172_n_8567) );
in01f10 FE_OFC2173_n_8567 ( .a(FE_OFN2171_n_8567), .o(FE_OFN2173_n_8567) );
in01f10 FE_OFC2174_n_8567 ( .a(FE_OFN2171_n_8567), .o(FE_OFN2174_n_8567) );
in01f10 FE_OFC2175_n_8567 ( .a(FE_OFN2172_n_8567), .o(FE_OFN2175_n_8567) );
in01f40 FE_OFC2176_n_8567 ( .a(FE_OFN1378_n_8567), .o(FE_OFN2176_n_8567) );
in01f20 FE_OFC2177_n_8567 ( .a(FE_OFN2176_n_8567), .o(FE_OFN2177_n_8567) );
in01f08 FE_OFC2178_n_8567 ( .a(FE_OFN2176_n_8567), .o(FE_OFN2178_n_8567) );
in01f20 FE_OFC2179_n_8567 ( .a(FE_OFN2176_n_8567), .o(FE_OFN2179_n_8567) );
in01s06 FE_OFC217_n_9889 ( .a(FE_OFN216_n_9889), .o(FE_OFN217_n_9889) );
in01f20 FE_OFC2180_n_8567 ( .a(FE_OFN2176_n_8567), .o(FE_OFN2180_n_8567) );
in01f10 FE_OFC2181_n_8567 ( .a(FE_OFN1394_n_8567), .o(FE_OFN2181_n_8567) );
in01f10 FE_OFC2182_n_8567 ( .a(FE_OFN2181_n_8567), .o(FE_OFN2182_n_8567) );
in01f10 FE_OFC2183_n_8567 ( .a(FE_OFN1394_n_8567), .o(FE_OFN2183_n_8567) );
in01f20 FE_OFC2184_n_8567 ( .a(FE_OFN2183_n_8567), .o(FE_OFN2184_n_8567) );
in01f10 FE_OFC2185_n_8567 ( .a(FE_OFN2181_n_8567), .o(FE_OFN2185_n_8567) );
in01f20 FE_OFC2186_n_8567 ( .a(FE_OFN1410_n_8567), .o(FE_OFN2186_n_8567) );
in01f10 FE_OFC2187_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2187_n_8567) );
in01f10 FE_OFC2188_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2188_n_8567) );
in01f06 FE_OFC2189_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2189_n_8567) );
in01m02 FE_OFC218_n_9853 ( .a(n_9853), .o(FE_OFN218_n_9853) );
in01f08 FE_OFC2190_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2190_n_8567) );
in01f10 FE_OFC2191_n_8567 ( .a(FE_OFN2186_n_8567), .o(FE_OFN2191_n_8567) );
in01f08 FE_OFC2192_n_16779 ( .a(FE_OFN1430_n_16779), .o(FE_OFN2192_n_16779) );
in01f06 FE_OFC2193_n_9163 ( .a(FE_OFN1447_n_9163), .o(FE_OFN2193_n_9163) );
in01f08 FE_OFC2194_n_9163 ( .a(FE_OFN1447_n_9163), .o(FE_OFN2194_n_9163) );
in01f02 FE_OFC2195_n_9163 ( .a(FE_OFN1447_n_9163), .o(FE_OFN2195_n_9163) );
in01f01 FE_OFC2196_n_9163 ( .a(FE_OFN1447_n_9163), .o(FE_OFN2196_n_9163) );
in01f10 FE_OFC2197_n_10256 ( .a(n_10256), .o(FE_OFN2197_n_10256) );
in01f20 FE_OFC2198_n_10256 ( .a(FE_OFN2197_n_10256), .o(FE_OFN2198_n_10256) );
in01f10 FE_OFC2199_n_10256 ( .a(n_10256), .o(FE_OFN2199_n_10256) );
in01s06 FE_OFC219_n_9853 ( .a(FE_OFN218_n_9853), .o(FE_OFN219_n_9853) );
in01f02 FE_OFC21_n_9372 ( .a(FE_OFN1434_n_9372), .o(FE_OFN21_n_9372) );
in01f20 FE_OFC2200_n_10256 ( .a(FE_OFN2199_n_10256), .o(FE_OFN2200_n_10256) );
in01f04 FE_OFC2201_n_12042 ( .a(n_15969), .o(FE_OFN2201_n_12042) );
in01f03 FE_OFC2202_n_12042 ( .a(n_15969), .o(FE_OFN2202_n_12042) );
in01f08 FE_OFC2203_n_12042 ( .a(FE_OFN2201_n_12042), .o(FE_OFN2203_n_12042) );
in01f01 FE_OFC2204_n_12028 ( .a(FE_OFN1576_n_12028), .o(FE_OFN2204_n_12028) );
in01f08 FE_OFC2205_n_10538 ( .a(FE_OFN1514_n_10538), .o(FE_OFN2205_n_10538) );
in01f04 FE_OFC2206_n_10892 ( .a(FE_OFN1520_n_10892), .o(FE_OFN2206_n_10892) );
in01f04 FE_OFC2207_n_10892 ( .a(FE_OFN1520_n_10892), .o(FE_OFN2207_n_10892) );
in01f08 FE_OFC2208_n_11795 ( .a(FE_OFN1459_n_11795), .o(FE_OFN2208_n_11795) );
in01f08 FE_OFC2209_n_11027 ( .a(FE_OCP_RBN2274_n_10268), .o(FE_OFN2209_n_11027) );
in01s02 FE_OFC220_n_9846 ( .a(n_9846), .o(FE_OFN220_n_9846) );
in01f06 FE_OFC2210_n_11027 ( .a(FE_OCP_RBN2274_n_10268), .o(FE_OFN2210_n_11027) );
in01f08 FE_OFC2211_n_8407 ( .a(FE_OFN2083_n_8407), .o(FE_OFN2211_n_8407) );
in01f10 FE_OFC2212_n_8407 ( .a(FE_OFN2211_n_8407), .o(FE_OFN2212_n_8407) );
in01f01 FE_OFC2213_n_15366 ( .a(FE_OFN995_n_15366), .o(FE_OFN2213_n_15366) );
in01f20 FE_OFC2214_n_15366 ( .a(FE_OFN995_n_15366), .o(FE_OFN2214_n_15366) );
in01f04 FE_OFC2215_n_15366 ( .a(FE_OFN2213_n_15366), .o(FE_OFN2215_n_15366) );
in01f08 FE_OFC2216_n_10143 ( .a(FE_OFN1531_n_10143), .o(FE_OFN2216_n_10143) );
in01s06 FE_OFC221_n_9846 ( .a(FE_OFN220_n_9846), .o(FE_OFN221_n_9846) );
in01m02 FE_OFC222_n_9844 ( .a(n_9844), .o(FE_OFN222_n_9844) );
in01m06 FE_OFC223_n_9844 ( .a(FE_OFN222_n_9844), .o(FE_OFN223_n_9844) );
in01f10 FE_OFC2240_g52675_p ( .a(FE_OFN1470_g52675_p), .o(FE_OFN2240_g52675_p) );
in01f04 FE_OFC2241_g52675_p ( .a(FE_OFN2240_g52675_p), .o(FE_OFN2241_g52675_p) );
in01f08 FE_OFC2242_g52675_p ( .a(FE_OFN2240_g52675_p), .o(FE_OFN2242_g52675_p) );
in01f20 FE_OFC2243_g52675_p ( .a(FE_OFN2240_g52675_p), .o(FE_OFN2243_g52675_p) );
in01f02 FE_OFC2244_n_4792 ( .a(n_4792), .o(FE_OFN2244_n_4792) );
in01f02 FE_OFC2245_n_4792 ( .a(FE_OFN2244_n_4792), .o(FE_OFN2245_n_4792) );
in01f02 FE_OFC2246_n_2113 ( .a(n_2113), .o(FE_OFN2246_n_2113) );
in01f02 FE_OFC2247_n_2113 ( .a(FE_OFN2246_n_2113), .o(FE_OFN2247_n_2113) );
in01f02 FE_OFC2248_n_1790 ( .a(n_1790), .o(FE_OFN2248_n_1790) );
in01f04 FE_OFC2249_n_1790 ( .a(FE_OFN2248_n_1790), .o(FE_OFN2249_n_1790) );
in01f10 FE_OFC224_n_9122 ( .a(n_9122), .o(FE_OFN224_n_9122) );
in01f02 FE_OFC2250_n_2101 ( .a(n_2101), .o(FE_OFN2250_n_2101) );
in01f02 FE_OFC2251_n_2101 ( .a(FE_OFN2250_n_2101), .o(FE_OFN2251_n_2101) );
in01m04 FE_OFC2252_n_9687 ( .a(FE_OFN602_n_9687), .o(FE_OFN2252_n_9687) );
in01s04 FE_OFC2253_n_9687 ( .a(FE_OFN2252_n_9687), .o(FE_OFN2253_n_9687) );
in01s01 FE_OFC2254_n_9687 ( .a(FE_OFN2252_n_9687), .o(FE_OFN2254_n_9687) );
in01f04 FE_OFC2255_n_8060 ( .a(n_8060), .o(FE_OFN2255_n_8060) );
in01f02 FE_OFC2256_n_8060 ( .a(FE_OFN2255_n_8060), .o(FE_OFN2256_n_8060) );
in01f04 FE_OFC2257_n_8060 ( .a(FE_OFN2255_n_8060), .o(FE_OFN2257_n_8060) );
in01f08 FE_OFC2258_n_8060 ( .a(FE_OFN2255_n_8060), .o(FE_OFN2258_n_8060) );
in01f02 FE_OFC2259_n_2775 ( .a(n_2775), .o(FE_OFN2259_n_2775) );
in01f20 FE_OFC225_n_9122 ( .a(FE_OFN224_n_9122), .o(FE_OFN225_n_9122) );
in01f02 FE_OFC2260_n_2775 ( .a(FE_OFN2259_n_2775), .o(FE_OFN2260_n_2775) );
in01s02 FE_OFC226_n_9841 ( .a(n_9841), .o(FE_OFN226_n_9841) );
in01s06 FE_OFC227_n_9841 ( .a(FE_OFN226_n_9841), .o(FE_OFN227_n_9841) );
in01m02 FE_OFC228_n_9120 ( .a(n_9120), .o(FE_OFN228_n_9120) );
in01m06 FE_OFC229_n_9120 ( .a(FE_OFN228_n_9120), .o(FE_OFN229_n_9120) );
in01f02 FE_OFC230_n_9839 ( .a(n_9839), .o(FE_OFN230_n_9839) );
in01m08 FE_OFC231_n_9839 ( .a(FE_OFN230_n_9839), .o(FE_OFN231_n_9839) );
in01m06 FE_OFC232_n_9876 ( .a(n_9876), .o(FE_OFN232_n_9876) );
in01s10 FE_OFC233_n_9876 ( .a(FE_OFN232_n_9876), .o(FE_OFN233_n_9876) );
in01f02 FE_OFC234_n_9834 ( .a(n_9834), .o(FE_OFN234_n_9834) );
in01f06 FE_OFC235_n_9834 ( .a(FE_OFN234_n_9834), .o(FE_OFN235_n_9834) );
in01f02 FE_OFC236_n_9118 ( .a(n_9118), .o(FE_OFN236_n_9118) );
in01f06 FE_OFC237_n_9118 ( .a(FE_OFN236_n_9118), .o(FE_OFN237_n_9118) );
in01f20 FE_OFC238_n_9832 ( .a(n_9832), .o(FE_OFN238_n_9832) );
in01f20 FE_OFC239_n_9832 ( .a(FE_OFN238_n_9832), .o(FE_OFN239_n_9832) );
in01m02 FE_OFC240_n_9830 ( .a(n_9830), .o(FE_OFN240_n_9830) );
in01m06 FE_OFC241_n_9830 ( .a(FE_OFN240_n_9830), .o(FE_OFN241_n_9830) );
in01s04 FE_OFC242_n_9116 ( .a(n_9116), .o(FE_OFN242_n_9116) );
in01s08 FE_OFC243_n_9116 ( .a(FE_OFN242_n_9116), .o(FE_OFN243_n_9116) );
in01s02 FE_OFC244_n_9114 ( .a(n_9114), .o(FE_OFN244_n_9114) );
in01s04 FE_OFC245_n_9114 ( .a(FE_OFN244_n_9114), .o(FE_OFN245_n_9114) );
in01f02 FE_OFC246_n_9112 ( .a(n_9112), .o(FE_OFN246_n_9112) );
in01f06 FE_OFC247_n_9112 ( .a(FE_OFN246_n_9112), .o(FE_OFN247_n_9112) );
in01m02 FE_OFC248_n_9789 ( .a(n_9789), .o(FE_OFN248_n_9789) );
in01m06 FE_OFC250_n_9789 ( .a(FE_OFN248_n_9789), .o(FE_OFN250_n_9789) );
in01f06 FE_OFC251_n_9868 ( .a(n_9868), .o(FE_OFN251_n_9868) );
in01m10 FE_OFC252_n_9868 ( .a(FE_OFN251_n_9868), .o(FE_OFN252_n_9868) );
in01s04 FE_OFC253_n_9825 ( .a(n_9825), .o(FE_OFN253_n_9825) );
in01s08 FE_OFC254_n_9825 ( .a(FE_OFN253_n_9825), .o(FE_OFN254_n_9825) );
in01s02 FE_OFC255_n_8969 ( .a(n_8969), .o(FE_OFN255_n_8969) );
in01s04 FE_OFC256_n_8969 ( .a(FE_OFN255_n_8969), .o(FE_OFN256_n_8969) );
in01f02 FE_OFC257_n_9862 ( .a(n_9862), .o(FE_OFN257_n_9862) );
in01f06 FE_OFC258_n_9862 ( .a(FE_OFN257_n_9862), .o(FE_OFN258_n_9862) );
in01m02 FE_OFC259_n_9860 ( .a(n_9860), .o(FE_OFN259_n_9860) );
in01m06 FE_OFC260_n_9860 ( .a(FE_OFN259_n_9860), .o(FE_OFN260_n_9860) );
in01f20 FE_OFC261_n_9851 ( .a(n_9851), .o(FE_OFN261_n_9851) );
in01f20 FE_OFC262_n_9851 ( .a(FE_OFN261_n_9851), .o(FE_OFN262_n_9851) );
in01m04 FE_OFC263_n_9849 ( .a(n_9849), .o(FE_OFN263_n_9849) );
in01m08 FE_OFC264_n_9849 ( .a(FE_OFN263_n_9849), .o(FE_OFN264_n_9849) );
in01m06 FE_OFC265_n_9884 ( .a(n_9884), .o(FE_OFN265_n_9884) );
in01s10 FE_OFC266_n_9884 ( .a(FE_OFN265_n_9884), .o(FE_OFN266_n_9884) );
in01m02 FE_OFC267_n_9880 ( .a(n_9880), .o(FE_OFN267_n_9880) );
in01m06 FE_OFC268_n_9880 ( .a(FE_OFN267_n_9880), .o(FE_OFN268_n_9880) );
in01m02 FE_OFC269_n_9836 ( .a(n_9836), .o(FE_OFN269_n_9836) );
in01s08 FE_OFC270_n_9836 ( .a(FE_OFN269_n_9836), .o(FE_OFN270_n_9836) );
in01f02 FE_OFC271_n_9828 ( .a(n_9828), .o(FE_OFN271_n_9828) );
in01f08 FE_OFC272_n_9828 ( .a(FE_OFN271_n_9828), .o(FE_OFN272_n_9828) );
in01f40 FE_OFC275_n_9941 ( .a(n_9941), .o(FE_OFN275_n_9941) );
in01f40 FE_OFC276_n_9941 ( .a(FE_OFN275_n_9941), .o(FE_OFN276_n_9941) );
in01m02 FE_OFC2_n_4778 ( .a(FE_OFN1_n_4778), .o(FE_OFN2_n_4778) );
in01m02 FE_OFC334_g66081_p ( .a(g66081_p), .o(FE_OFN334_g66081_p) );
in01m06 FE_OFC335_g66081_p ( .a(FE_OFN334_g66081_p), .o(FE_OFN335_g66081_p) );
in01m02 FE_OFC336_g66089_p ( .a(g66089_p), .o(FE_OFN336_g66089_p) );
in01m06 FE_OFC337_g66089_p ( .a(FE_OFN336_g66089_p), .o(FE_OFN337_g66089_p) );
in01f01 FE_OFC365_n_4093 ( .a(FE_OFN1245_n_4093), .o(FE_OFN365_n_4093) );
in01f02 FE_OFC369_n_4092 ( .a(FE_OFN1237_n_4092), .o(FE_OFN369_n_4092) );
in01f02 FE_OFC3_n_4778 ( .a(FE_OFN1_n_4778), .o(FE_OFN3_n_4778) );
in01f08 FE_OFC514_n_9697 ( .a(n_9697), .o(FE_OFN514_n_9697) );
in01f10 FE_OFC515_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN515_n_9697) );
in01s06 FE_OFC516_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN516_n_9697) );
in01f03 FE_OFC517_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN517_n_9697) );
in01s02 FE_OFC518_n_9697 ( .a(FE_OFN514_n_9697), .o(TIMEBOOST_net_21135) );
in01s02 FE_OFC519_n_9697 ( .a(FE_OFN514_n_9697), .o(FE_OFN519_n_9697) );
in01s04 FE_OFC523_n_9428 ( .a(FE_OFN1646_n_9428), .o(FE_OFN523_n_9428) );
in01f20 FE_OFC524_n_9899 ( .a(n_9899), .o(FE_OFN524_n_9899) );
in01s06 FE_OFC525_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN525_n_9899) );
in01s06 FE_OFC526_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN526_n_9899) );
in01f40 FE_OFC527_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN527_n_9899) );
in01s02 FE_OFC528_n_9899 ( .a(FE_OFN524_n_9899), .o(TIMEBOOST_net_21131) );
in01m06 FE_OFC529_n_9899 ( .a(FE_OFN524_n_9899), .o(FE_OFN529_n_9899) );
in01f10 FE_OFC530_n_9823 ( .a(n_9823), .o(FE_OFN530_n_9823) );
in01f01 FE_OFC531_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN531_n_9823) );
in01s02 FE_OFC532_n_9823 ( .a(FE_OFN530_n_9823), .o(TIMEBOOST_net_20140) );
in01s08 FE_OFC533_n_9823 ( .a(FE_OFN530_n_9823), .o(TIMEBOOST_net_21133) );
in01m01 FE_OFC534_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN534_n_9823) );
in01f20 FE_OFC535_n_9823 ( .a(FE_OFN530_n_9823), .o(FE_OFN535_n_9823) );
in01f10 FE_OFC537_n_9690 ( .a(n_9690), .o(FE_OFN537_n_9690) );
in01f01 FE_OFC539_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN539_n_9690) );
in01m01 FE_OFC540_n_9690 ( .a(FE_OFN537_n_9690), .o(TIMEBOOST_net_21225) );
in01f10 FE_OFC541_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN541_n_9690) );
in01m01 FE_OFC542_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN542_n_9690) );
in01m01 FE_OFC543_n_9690 ( .a(FE_OFN537_n_9690), .o(FE_OFN543_n_9690) );
in01s04 FE_OFC548_n_9477 ( .a(FE_OFN1664_n_9477), .o(FE_OFN548_n_9477) );
in01m01 FE_OFC549_n_9864 ( .a(n_9864), .o(FE_OFN549_n_9864) );
in01f06 FE_OFC550_n_9864 ( .a(n_9864), .o(FE_OFN550_n_9864) );
in01s02 FE_OFC551_n_9864 ( .a(FE_OFN549_n_9864), .o(FE_OFN551_n_9864) );
in01s01 FE_OFC552_n_9864 ( .a(FE_OFN549_n_9864), .o(FE_OFN552_n_9864) );
in01s02 FE_OFC553_n_9864 ( .a(FE_OFN550_n_9864), .o(FE_OFN553_n_9864) );
in01s06 FE_OFC554_n_9864 ( .a(FE_OFN550_n_9864), .o(TIMEBOOST_net_20138) );
in01f10 FE_OFC555_n_9864 ( .a(FE_OFN550_n_9864), .o(FE_OFN555_n_9864) );
in01m01 FE_OFC556_n_9864 ( .a(FE_OFN550_n_9864), .o(FE_OFN556_n_9864) );
in01f01 FE_OFC557_n_9895 ( .a(n_9895), .o(FE_OFN557_n_9895) );
in01f02 FE_OFC558_n_9895 ( .a(n_9895), .o(FE_OFN558_n_9895) );
in01m01 FE_OFC559_n_9895 ( .a(FE_OFN557_n_9895), .o(FE_OFN559_n_9895) );
in01m03 FE_OFC560_n_9895 ( .a(FE_OFN557_n_9895), .o(FE_OFN560_n_9895) );
in01f02 FE_OFC561_n_9895 ( .a(FE_OFN558_n_9895), .o(FE_OFN561_n_9895) );
in01f06 FE_OFC562_n_9895 ( .a(FE_OFN558_n_9895), .o(FE_OFN562_n_9895) );
in01f02 FE_OFC563_n_9895 ( .a(FE_OFN558_n_9895), .o(FE_OFN563_n_9895) );
in01m02 FE_OFC564_n_9895 ( .a(FE_OFN558_n_9895), .o(FE_OFN564_n_9895) );
in01f03 FE_OFC568_n_9528 ( .a(FE_OFN1683_n_9528), .o(FE_OFN568_n_9528) );
in01f04 FE_OFC569_n_9528 ( .a(FE_OFN1683_n_9528), .o(FE_OFN569_n_9528) );
in01f08 FE_OFC572_n_9502 ( .a(FE_OFN1652_n_9502), .o(FE_OFN572_n_9502) );
in01f04 FE_OFC573_n_9902 ( .a(n_9902), .o(FE_OFN573_n_9902) );
in01f04 FE_OFC574_n_9902 ( .a(FE_OFN573_n_9902), .o(FE_OFN574_n_9902) );
in01f04 FE_OFC575_n_9902 ( .a(FE_OFN573_n_9902), .o(FE_OFN575_n_9902) );
in01f04 FE_OFC576_n_9902 ( .a(FE_OFN573_n_9902), .o(FE_OFN576_n_9902) );
in01f06 FE_OFC577_n_9902 ( .a(FE_OFN573_n_9902), .o(FE_OFN577_n_9902) );
in01f06 FE_OFC579_n_9531 ( .a(FE_OFN1629_n_9531), .o(FE_OFN579_n_9531) );
in01f08 FE_OFC580_n_9531 ( .a(FE_OFN1629_n_9531), .o(FE_OFN580_n_9531) );
in01m06 FE_OFC582_n_9692 ( .a(n_9692), .o(FE_OFN582_n_9692) );
in01f10 FE_OFC583_n_9692 ( .a(n_9692), .o(FE_OFN583_n_9692) );
in01f02 FE_OFC584_n_9692 ( .a(FE_OFN582_n_9692), .o(FE_OFN584_n_9692) );
in01f10 FE_OFC585_n_9692 ( .a(FE_OFN583_n_9692), .o(FE_OFN585_n_9692) );
in01m04 FE_OFC587_n_9692 ( .a(FE_OFN582_n_9692), .o(FE_OFN587_n_9692) );
in01f02 FE_OFC588_n_9692 ( .a(FE_OFN582_n_9692), .o(FE_OFN588_n_9692) );
in01m02 FE_OFC589_n_9692 ( .a(FE_OFN582_n_9692), .o(FE_OFN589_n_9692) );
in01f02 FE_OFC590_n_9694 ( .a(n_9694), .o(FE_OFN590_n_9694) );
in01m01 FE_OFC591_n_9694 ( .a(n_9694), .o(FE_OFN591_n_9694) );
in01m03 FE_OFC592_n_9694 ( .a(FE_OFN590_n_9694), .o(FE_OFN592_n_9694) );
in01s04 FE_OFC593_n_9694 ( .a(FE_OFN591_n_9694), .o(FE_OFN593_n_9694) );
in01m04 FE_OFC595_n_9694 ( .a(FE_OFN590_n_9694), .o(FE_OFN595_n_9694) );
in01m03 FE_OFC596_n_9694 ( .a(FE_OFN590_n_9694), .o(FE_OFN596_n_9694) );
in01m02 FE_OFC597_n_9694 ( .a(FE_OFN590_n_9694), .o(TIMEBOOST_net_13969) );
in01f02 FE_OFC598_n_9687 ( .a(n_9687), .o(FE_OFN598_n_9687) );
in01f01 FE_OFC599_n_9687 ( .a(n_9687), .o(FE_OFN599_n_9687) );
in01m02 FE_OFC600_n_9687 ( .a(FE_OFN598_n_9687), .o(FE_OFN600_n_9687) );
in01m06 FE_OFC601_n_9687 ( .a(FE_OFN598_n_9687), .o(FE_OFN601_n_9687) );
in01m04 FE_OFC602_n_9687 ( .a(FE_OFN598_n_9687), .o(FE_OFN602_n_9687) );
in01s04 FE_OFC603_n_9687 ( .a(FE_OFN599_n_9687), .o(FE_OFN603_n_9687) );
in01f10 FE_OFC605_n_9904 ( .a(n_9904), .o(FE_OFN605_n_9904) );
in01s02 FE_OFC606_n_9904 ( .a(FE_OFN605_n_9904), .o(TIMEBOOST_net_21223) );
in01f10 FE_OFC607_n_9904 ( .a(FE_OFN605_n_9904), .o(FE_OFN607_n_9904) );
in01s01 FE_OFC608_n_9904 ( .a(FE_OFN605_n_9904), .o(FE_OFN608_n_9904) );
in01f20 FE_OFC611_n_4501 ( .a(n_4501), .o(FE_OFN611_n_4501) );
in01m10 FE_OFC612_n_4501 ( .a(FE_OFN611_n_4501), .o(FE_OFN612_n_4501) );
in01m10 FE_OFC613_n_4501 ( .a(FE_OFN611_n_4501), .o(FE_OFN613_n_4501) );
in01f08 FE_OFC614_n_4501 ( .a(FE_OFN611_n_4501), .o(FE_OFN614_n_4501) );
in01m20 FE_OFC615_n_4501 ( .a(FE_OFN611_n_4501), .o(FE_OFN615_n_4501) );
in01f10 FE_OFC618_n_4490 ( .a(FE_OFN1661_n_4490), .o(FE_OFN618_n_4490) );
in01f04 FE_OFC619_n_4490 ( .a(FE_OFN1661_n_4490), .o(FE_OFN619_n_4490) );
in01m10 FE_OFC620_n_4490 ( .a(FE_OFN1661_n_4490), .o(FE_OFN620_n_4490) );
in01f20 FE_OFC621_n_4409 ( .a(n_4409), .o(FE_OFN621_n_4409) );
in01m10 FE_OFC622_n_4409 ( .a(FE_OFN621_n_4409), .o(FE_OFN622_n_4409) );
in01f08 FE_OFC623_n_4409 ( .a(FE_OFN621_n_4409), .o(FE_OFN623_n_4409) );
in01m10 FE_OFC624_n_4409 ( .a(FE_OFN621_n_4409), .o(FE_OFN624_n_4409) );
in01m20 FE_OFC625_n_4409 ( .a(FE_OFN621_n_4409), .o(FE_OFN625_n_4409) );
in01f20 FE_OFC627_n_4454 ( .a(n_4454), .o(FE_OFN627_n_4454) );
in01m02 FE_OFC628_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN628_n_4454) );
in01m03 FE_OFC629_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN629_n_4454) );
in01m03 FE_OFC630_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN630_n_4454) );
in01f08 FE_OFC631_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN631_n_4454) );
in01m10 FE_OFC632_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN632_n_4454) );
in01m08 FE_OFC633_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN633_n_4454) );
in01m10 FE_OFC634_n_4454 ( .a(FE_OFN627_n_4454), .o(FE_OFN634_n_4454) );
in01f20 FE_OFC636_n_4669 ( .a(FE_OFN1682_n_4669), .o(FE_OFN636_n_4669) );
in01m02 FE_OFC638_n_4669 ( .a(FE_OFN1682_n_4669), .o(FE_OFN638_n_4669) );
in01m20 FE_OFC639_n_4669 ( .a(FE_OFN1682_n_4669), .o(FE_OFN639_n_4669) );
in01m20 FE_OFC640_n_4669 ( .a(FE_OFN1681_n_4669), .o(FE_OFN640_n_4669) );
in01f20 FE_OFC641_n_4677 ( .a(n_4677), .o(FE_OFN641_n_4677) );
in01m10 FE_OFC642_n_4677 ( .a(FE_OFN641_n_4677), .o(FE_OFN642_n_4677) );
in01f10 FE_OFC643_n_4677 ( .a(FE_OFN641_n_4677), .o(FE_OFN643_n_4677) );
in01m20 FE_OFC644_n_4677 ( .a(FE_OFN641_n_4677), .o(FE_OFN644_n_4677) );
in01f20 FE_OFC645_n_4497 ( .a(n_4497), .o(FE_OFN645_n_4497) );
in01m10 FE_OFC646_n_4497 ( .a(FE_OFN645_n_4497), .o(FE_OFN646_n_4497) );
in01m10 FE_OFC647_n_4497 ( .a(FE_OFN645_n_4497), .o(FE_OFN647_n_4497) );
in01f10 FE_OFC648_n_4497 ( .a(FE_OFN645_n_4497), .o(FE_OFN648_n_4497) );
in01m20 FE_OFC649_n_4497 ( .a(FE_OFN645_n_4497), .o(FE_OFN649_n_4497) );
in01f10 FE_OFC650_n_4508 ( .a(n_4508), .o(FE_OFN650_n_4508) );
in01f08 FE_OFC651_n_4508 ( .a(FE_OFN650_n_4508), .o(FE_OFN651_n_4508) );
in01m10 FE_OFC652_n_4508 ( .a(FE_OFN650_n_4508), .o(FE_OFN652_n_4508) );
in01m10 FE_OFC653_n_4508 ( .a(FE_OFN650_n_4508), .o(FE_OFN653_n_4508) );
in01f08 FE_OFC654_n_4508 ( .a(FE_OFN650_n_4508), .o(FE_OFN654_n_4508) );
in01f20 FE_OFC658_n_4392 ( .a(n_4392), .o(FE_OFN658_n_4392) );
in01f10 FE_OFC659_n_4392 ( .a(FE_OFN658_n_4392), .o(FE_OFN659_n_4392) );
in01m10 FE_OFC660_n_4392 ( .a(FE_OFN658_n_4392), .o(FE_OFN660_n_4392) );
in01m20 FE_OFC661_n_4392 ( .a(FE_OFN658_n_4392), .o(FE_OFN661_n_4392) );
in01m10 FE_OFC662_n_4392 ( .a(FE_OFN658_n_4392), .o(FE_OFN662_n_4392) );
in01f10 FE_OFC663_n_4495 ( .a(n_4495), .o(FE_OFN663_n_4495) );
in01f06 FE_OFC664_n_4495 ( .a(FE_OFN663_n_4495), .o(FE_OFN664_n_4495) );
in01m08 FE_OFC665_n_4495 ( .a(FE_OFN663_n_4495), .o(FE_OFN665_n_4495) );
in01m10 FE_OFC666_n_4495 ( .a(FE_OFN663_n_4495), .o(FE_OFN666_n_4495) );
in01m10 FE_OFC667_n_4495 ( .a(FE_OFN663_n_4495), .o(FE_OFN667_n_4495) );
in01m20 FE_OFC668_n_4505 ( .a(n_4505), .o(FE_OFN668_n_4505) );
in01m10 FE_OFC669_n_4505 ( .a(FE_OFN668_n_4505), .o(FE_OFN669_n_4505) );
in01m20 FE_OFC670_n_4505 ( .a(FE_OFN668_n_4505), .o(FE_OFN670_n_4505) );
in01m06 FE_OFC671_n_4505 ( .a(FE_OFN668_n_4505), .o(FE_OFN671_n_4505) );
in01m20 FE_OFC672_n_4505 ( .a(FE_OFN668_n_4505), .o(FE_OFN672_n_4505) );
in01f01 FE_OFC678_n_4460 ( .a(FE_OFN1636_n_4460), .o(FE_OFN678_n_4460) );
in01m08 FE_OFC679_n_4460 ( .a(FE_OFN1636_n_4460), .o(FE_OFN679_n_4460) );
in01f10 FE_OFC681_n_4460 ( .a(FE_OFN1636_n_4460), .o(FE_OFN681_n_4460) );
in01f20 FE_OFC682_n_4460 ( .a(FE_OFN1636_n_4460), .o(FE_OFN682_n_4460) );
in01f20 FE_OFC683_n_4417 ( .a(n_4417), .o(FE_OFN683_n_4417) );
in01m08 FE_OFC684_n_4417 ( .a(FE_OFN683_n_4417), .o(FE_OFN684_n_4417) );
in01m08 FE_OFC685_n_4417 ( .a(FE_OFN683_n_4417), .o(FE_OFN685_n_4417) );
in01f20 FE_OFC686_n_4417 ( .a(FE_OFN683_n_4417), .o(FE_OFN686_n_4417) );
in01m10 FE_OFC687_n_4417 ( .a(FE_OFN683_n_4417), .o(FE_OFN687_n_4417) );
in01m10 FE_OFC689_n_4438 ( .a(FE_OFN1622_n_4438), .o(FE_OFN689_n_4438) );
in01f06 FE_OFC697_n_16760 ( .a(FE_OFN1026_n_16760), .o(FE_OFN697_n_16760) );
in01f04 FE_OFC698_n_7845 ( .a(n_7845), .o(FE_OFN698_n_7845) );
in01f04 FE_OFC699_n_7845 ( .a(FE_OFN698_n_7845), .o(FE_OFN699_n_7845) );
in01f04 FE_OFC700_n_7845 ( .a(FE_OFN698_n_7845), .o(FE_OFN700_n_7845) );
in01f03 FE_OFC701_n_7845 ( .a(FE_OFN698_n_7845), .o(FE_OFN701_n_7845) );
in01f04 FE_OFC702_n_7845 ( .a(FE_OFN698_n_7845), .o(FE_OFN702_n_7845) );
in01f01 FE_OFC703_n_8069 ( .a(n_8069), .o(FE_OFN703_n_8069) );
in01f04 FE_OFC704_n_8069 ( .a(FE_OFN703_n_8069), .o(FE_OFN704_n_8069) );
in01f08 FE_OFC705_n_8119 ( .a(n_8119), .o(FE_OFN705_n_8119) );
in01f08 FE_OFC706_n_8119 ( .a(FE_OFN705_n_8119), .o(FE_OFN706_n_8119) );
in01f08 FE_OFC707_n_8119 ( .a(FE_OFN705_n_8119), .o(FE_OFN707_n_8119) );
in01f08 FE_OFC708_n_8232 ( .a(n_8232), .o(FE_OFN708_n_8232) );
in01f10 FE_OFC709_n_8232 ( .a(FE_OFN708_n_8232), .o(FE_OFN709_n_8232) );
in01f08 FE_OFC710_n_8232 ( .a(FE_OFN708_n_8232), .o(FE_OFN710_n_8232) );
in01f06 FE_OFC711_n_8140 ( .a(n_8140), .o(FE_OFN711_n_8140) );
in01f08 FE_OFC712_n_8140 ( .a(FE_OFN711_n_8140), .o(FE_OFN712_n_8140) );
in01f06 FE_OFC713_n_8140 ( .a(FE_OFN711_n_8140), .o(FE_OFN713_n_8140) );
in01f08 FE_OFC714_n_8140 ( .a(FE_OFN711_n_8140), .o(FE_OFN714_n_8140) );
in01f04 FE_OFC715_n_8176 ( .a(n_8176), .o(FE_OFN715_n_8176) );
in01f08 FE_OFC716_n_8176 ( .a(FE_OFN715_n_8176), .o(FE_OFN716_n_8176) );
in01f06 FE_OFC717_n_8176 ( .a(FE_OFN715_n_8176), .o(FE_OFN717_n_8176) );
in01f10 FE_OFC718_n_8060 ( .a(FE_OFN2258_n_8060), .o(FE_OFN718_n_8060) );
in01f10 FE_OFC719_n_8060 ( .a(FE_OFN718_n_8060), .o(FE_OFN719_n_8060) );
in01m10 FE_OFC720_n_8060 ( .a(FE_OFN718_n_8060), .o(FE_OFN720_n_8060) );
in01f08 FE_OFC732_n_7498 ( .a(FE_OFN1156_n_7498), .o(FE_OFN732_n_7498) );
in01m04 FE_OFC775_n_15366 ( .a(FE_OFN2215_n_15366), .o(FE_OFN775_n_15366) );
in01m08 FE_OFC776_n_15366 ( .a(FE_OFN2215_n_15366), .o(FE_OFN776_n_15366) );
in01f02 FE_OFC777_n_4152 ( .a(n_4152), .o(FE_OFN777_n_4152) );
in01f06 FE_OFC778_n_4152 ( .a(FE_OFN777_n_4152), .o(FE_OFN778_n_4152) );
in01f02 FE_OFC779_n_2746 ( .a(n_2746), .o(FE_OFN779_n_2746) );
in01f02 FE_OFC780_n_2746 ( .a(FE_OFN779_n_2746), .o(FE_OFN780_n_2746) );
in01m01 FE_OFC781_n_2746 ( .a(FE_OFN779_n_2746), .o(FE_OFN781_n_2746) );
in01f08 FE_OFC782_n_2678 ( .a(n_2678), .o(FE_OFN782_n_2678) );
in01f02 FE_OFC783_n_2678 ( .a(n_2678), .o(FE_OFN783_n_2678) );
in01f08 FE_OFC784_n_2678 ( .a(FE_OFN782_n_2678), .o(FE_OFN784_n_2678) );
in01f08 FE_OFC785_n_2678 ( .a(FE_OFN782_n_2678), .o(FE_OFN785_n_2678) );
in01f06 FE_OFC786_n_2678 ( .a(FE_OFN782_n_2678), .o(FE_OFN786_n_2678) );
in01f04 FE_OFC787_n_2678 ( .a(FE_OFN783_n_2678), .o(FE_OFN787_n_2678) );
in01f04 FE_OFC789_n_2678 ( .a(FE_OFN782_n_2678), .o(FE_OFN789_n_2678) );
in01f01 FE_OFC792_n_2547 ( .a(n_2547), .o(FE_OFN792_n_2547) );
in01f02 FE_OFC793_n_2547 ( .a(FE_OFN792_n_2547), .o(FE_OFN793_n_2547) );
in01m02 FE_OFC794_n_2520 ( .a(n_2520), .o(FE_OFN794_n_2520) );
in01m06 FE_OFC795_n_2520 ( .a(FE_OFN794_n_2520), .o(FE_OFN795_n_2520) );
in01f08 FE_OFC877_g64577_p ( .a(FE_OFN1099_g64577_p), .o(FE_OFN877_g64577_p) );
in01f06 FE_OFC881_g64577_p ( .a(FE_OFN1086_g64577_p), .o(FE_OFN881_g64577_p) );
in01f10 FE_OFC882_g64577_p ( .a(FE_OFN1098_g64577_p), .o(FE_OFN882_g64577_p) );
in01m04 FE_OFC8_n_11877 ( .a(FE_OFN1020_n_11877), .o(FE_OFN8_n_11877) );
in01f02 FE_OFC900_n_4736 ( .a(n_4736), .o(FE_OFN900_n_4736) );
in01f10 FE_OFC901_n_4736 ( .a(n_4736), .o(FE_OFN901_n_4736) );
in01m01 FE_OFC902_n_4736 ( .a(FE_OFN900_n_4736), .o(FE_OFN902_n_4736) );
in01f06 FE_OFC903_n_4736 ( .a(FE_OFN900_n_4736), .o(FE_OFN903_n_4736) );
in01f08 FE_OFC904_n_4736 ( .a(FE_OFN901_n_4736), .o(FE_OFN904_n_4736) );
in01f10 FE_OFC905_n_4736 ( .a(FE_OFN901_n_4736), .o(FE_OFN905_n_4736) );
in01f10 FE_OFC906_n_4736 ( .a(FE_OFN901_n_4736), .o(FE_OFN906_n_4736) );
in01f06 FE_OFC908_n_4734 ( .a(FE_OFN1007_n_4734), .o(FE_OFN908_n_4734) );
in01f10 FE_OFC912_n_4727 ( .a(FE_OFN1052_n_4727), .o(FE_OFN912_n_4727) );
in01f20 FE_OFC915_n_4725 ( .a(n_4725), .o(FE_OFN915_n_4725) );
in01f08 FE_OFC916_n_4725 ( .a(FE_OFN915_n_4725), .o(FE_OFN916_n_4725) );
in01f10 FE_OFC917_n_4725 ( .a(FE_OFN915_n_4725), .o(FE_OFN917_n_4725) );
in01f20 FE_OFC918_n_4725 ( .a(FE_OFN915_n_4725), .o(FE_OFN918_n_4725) );
in01f20 FE_OFC923_n_4740 ( .a(FE_OFN1072_n_4740), .o(FE_OFN923_n_4740) );
in01f20 FE_OFC926_n_4730 ( .a(n_4730), .o(FE_OFN926_n_4730) );
in01f08 FE_OFC927_n_4730 ( .a(FE_OFN926_n_4730), .o(FE_OFN927_n_4730) );
in01f20 FE_OFC928_n_4730 ( .a(FE_OFN926_n_4730), .o(FE_OFN928_n_4730) );
in01m08 FE_OFC929_n_4730 ( .a(FE_OFN926_n_4730), .o(FE_OFN929_n_4730) );
in01f08 FE_OFC930_n_4730 ( .a(FE_OFN926_n_4730), .o(FE_OFN930_n_4730) );
in01f03 FE_OFC934_n_2292 ( .a(n_2292), .o(FE_OFN934_n_2292) );
in01f03 FE_OFC935_n_2292 ( .a(FE_OFN934_n_2292), .o(FE_OFN935_n_2292) );
in01f04 FE_OFC936_n_2292 ( .a(FE_OFN934_n_2292), .o(FE_OFN936_n_2292) );
in01f04 FE_OFC937_n_2292 ( .a(FE_OFN934_n_2292), .o(FE_OFN937_n_2292) );
in01f04 FE_OFC938_n_2292 ( .a(FE_OFN934_n_2292), .o(FE_OFN938_n_2292) );
in01m02 FE_OFC941_n_2047 ( .a(FE_OFN1002_n_2047), .o(FE_OFN941_n_2047) );
in01m06 FE_OFC944_n_2248 ( .a(n_2248), .o(FE_OFN944_n_2248) );
in01f06 FE_OFC945_n_2248 ( .a(FE_OFN944_n_2248), .o(FE_OFN945_n_2248) );
in01f02 FE_OFC946_n_2248 ( .a(FE_OFN944_n_2248), .o(FE_OFN946_n_2248) );
in01f08 FE_OFC947_n_2248 ( .a(FE_OFN2111_n_2248), .o(FE_OFN947_n_2248) );
in01f10 FE_OFC948_n_2248 ( .a(FE_OFN947_n_2248), .o(FE_OFN948_n_2248) );
in01f04 FE_OFC949_n_2055 ( .a(n_2055), .o(FE_OFN949_n_2055) );
in01f03 FE_OFC950_n_2055 ( .a(FE_OFN949_n_2055), .o(FE_OFN950_n_2055) );
in01m04 FE_OFC951_n_2055 ( .a(FE_OFN949_n_2055), .o(FE_OFN951_n_2055) );
in01f06 FE_OFC952_n_2055 ( .a(FE_OFN949_n_2055), .o(FE_OFN952_n_2055) );
in01m06 FE_OFC953_n_2055 ( .a(FE_OFN949_n_2055), .o(FE_OFN953_n_2055) );
in01f10 FE_OFC954_n_1699 ( .a(FE_OFN1783_n_1699), .o(FE_OFN954_n_1699) );
in01m08 FE_OFC955_n_1699 ( .a(FE_OFN954_n_1699), .o(FE_OFN955_n_1699) );
in01f10 FE_OFC956_n_1699 ( .a(FE_OFN954_n_1699), .o(FE_OFN956_n_1699) );
in01f08 FE_OFC957_n_2299 ( .a(n_2299), .o(FE_OFN957_n_2299) );
in01f06 FE_OFC958_n_2299 ( .a(FE_OFN957_n_2299), .o(FE_OFN958_n_2299) );
in01f08 FE_OFC959_n_2299 ( .a(FE_OFN957_n_2299), .o(FE_OFN959_n_2299) );
in01f02 FE_OFC966_n_2233 ( .a(n_2233), .o(FE_OFN966_n_2233) );
in01f02 FE_OFC967_n_2233 ( .a(FE_OFN966_n_2233), .o(FE_OFN967_n_2233) );
in01f20 FE_OFC968_n_13784 ( .a(FE_OFN1946_n_13784), .o(FE_OFN968_n_13784) );
in01f40 FE_OFC969_n_13784 ( .a(FE_OFN968_n_13784), .o(FE_OFN969_n_13784) );
in01f02 FE_OFC982_n_2700 ( .a(n_2700), .o(FE_OFN982_n_2700) );
in01f02 FE_OFC983_n_2700 ( .a(FE_OFN982_n_2700), .o(FE_OFN983_n_2700) );
in01f02 FE_OFC984_n_2697 ( .a(n_2697), .o(FE_OFN984_n_2697) );
in01f02 FE_OFC985_n_2697 ( .a(FE_OFN984_n_2697), .o(FE_OFN985_n_2697) );
in01f02 FE_OFC986_n_2696 ( .a(n_2696), .o(FE_OFN986_n_2696) );
in01f02 FE_OFC987_n_2696 ( .a(FE_OFN986_n_2696), .o(FE_OFN987_n_2696) );
in01f08 FE_OFC988_n_574 ( .a(n_574), .o(FE_OFN988_n_574) );
in01f10 FE_OFC989_n_574 ( .a(FE_OFN988_n_574), .o(FE_OFN989_n_574) );
in01f04 FE_OFC991_n_2373 ( .a(n_2373), .o(FE_OFN991_n_2373) );
in01f06 FE_OFC992_n_2373 ( .a(FE_OFN991_n_2373), .o(FE_OFN992_n_2373) );
in01f10 FE_OFC994_n_15366 ( .a(FE_OFN993_n_15366), .o(FE_OFN994_n_15366) );
in01f20 FE_OFC995_n_15366 ( .a(FE_OFN994_n_15366), .o(FE_OFN995_n_15366) );
in01f10 FE_OFC996_n_15366 ( .a(FE_OFN993_n_15366), .o(FE_OFN996_n_15366) );
in01f08 FE_OFC999_n_15978 ( .a(FE_OFN997_n_15978), .o(FE_OFN999_n_15978) );
in01f02 FE_OFC9_n_11877 ( .a(FE_OFN1020_n_11877), .o(FE_OFN9_n_11877) );
in01f20 FE_RC_0_0 ( .a(pci_target_unit_wishbone_master_first_data_is_burst_reg), .o(FE_RN_0_0) );
in01f20 FE_RC_1000_0 ( .a(n_3078), .o(FE_RN_695_0) );
oa12f08 FE_RC_1002_0 ( .a(FE_RN_694_0), .b(FE_RN_695_0), .c(FE_RN_693_0), .o(FE_RN_697_0) );
na02f10 FE_RC_1003_0 ( .a(n_2835), .b(n_419), .o(FE_RN_698_0) );
oa12f06 FE_RC_1004_0 ( .a(FE_RN_698_0), .b(n_2835), .c(n_419), .o(FE_RN_699_0) );
no02f06 FE_RC_1005_0 ( .a(FE_RN_697_0), .b(FE_RN_699_0), .o(FE_RN_700_0) );
na02f04 FE_RC_1006_0 ( .a(FE_RN_691_0), .b(FE_RN_700_0), .o(FE_RN_701_0) );
no02f02 FE_RC_1007_0 ( .a(FE_RN_684_0), .b(FE_RN_701_0), .o(FE_RN_702_0) );
na02f04 TIMEBOOST_cell_63204 ( .a(wbm_adr_o_15_), .b(g62067_sb), .o(TIMEBOOST_net_20549) );
na04f04 TIMEBOOST_cell_24167 ( .a(n_9744), .b(g57182_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q), .d(FE_OFN1408_n_8567), .o(n_11572) );
na04f04 TIMEBOOST_cell_67602 ( .a(g65019_da), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q), .c(TIMEBOOST_net_330), .d(g62575_sb), .o(n_6402) );
na02m06 TIMEBOOST_cell_69060 ( .a(FE_OFN612_n_4501), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q), .o(TIMEBOOST_net_21738) );
na03f01 TIMEBOOST_cell_69028 ( .a(n_3777), .b(FE_OFN625_n_4409), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_21722) );
in01f10 FE_RC_1014_0 ( .a(n_15998), .o(n_15746) );
in01f02 FE_RC_1015_0 ( .a(n_15998), .o(FE_RN_708_0) );
na02f03 FE_RC_1016_0 ( .a(FE_RN_708_0), .b(n_15924), .o(n_15754) );
in01f03 FE_RC_1017_0 ( .a(n_15924), .o(FE_RN_709_0) );
na02s02 TIMEBOOST_cell_51402 ( .a(TIMEBOOST_net_15918), .b(TIMEBOOST_net_11174), .o(TIMEBOOST_net_9349) );
na04f02 FE_RC_1019_0 ( .a(n_11097), .b(n_11788), .c(n_11095), .d(n_11096), .o(n_12545) );
in01f40 FE_RC_101_0 ( .a(wishbone_slave_unit_fifos_outGreyCount_2_), .o(FE_RN_57_0) );
in01f01 FE_RC_1020_0 ( .a(n_7822), .o(FE_RN_710_0) );
in01f02 FE_RC_1021_0 ( .a(n_12981), .o(FE_RN_711_0) );
na03s02 TIMEBOOST_cell_73345 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q), .b(FE_OFN606_n_9904), .c(g58060_sb), .o(TIMEBOOST_net_21000) );
na03f02 TIMEBOOST_cell_72621 ( .a(TIMEBOOST_net_16897), .b(FE_OFN1013_n_4734), .c(g64159_sb), .o(TIMEBOOST_net_13051) );
in01f02 FE_RC_1026_0 ( .a(n_9274), .o(FE_RN_713_0) );
in01f02 FE_RC_1027_0 ( .a(n_17043), .o(FE_RN_714_0) );
no02f02 FE_RC_1028_0 ( .a(FE_RN_714_0), .b(FE_RN_713_0), .o(FE_RN_715_0) );
na02s01 TIMEBOOST_cell_18141 ( .a(pci_target_unit_del_sync_be_out_reg_2__Q), .b(FE_OFN786_n_2678), .o(TIMEBOOST_net_5434) );
in01f40 FE_RC_102_0 ( .a(wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_), .o(FE_RN_58_0) );
ao22f02 FE_RC_1031_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q), .b(FE_OCP_RBN1968_FE_OFN1532_n_10143), .c(n_10185), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q), .o(n_10599) );
ao22f02 FE_RC_1032_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q), .b(FE_OFN2149_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q), .d(FE_OFN1522_n_10892), .o(n_10728) );
in01f02 FE_RC_1033_0 ( .a(FE_RN_716_0), .o(n_16317) );
na02f02 FE_RC_1034_0 ( .a(n_16313), .b(n_16445), .o(FE_RN_716_0) );
na04f04 FE_RC_1035_0 ( .a(n_12310), .b(n_12036), .c(n_12037), .d(n_12038), .o(n_12818) );
in01s01 FE_RC_1037_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q), .o(FE_RN_717_0) );
na02m04 TIMEBOOST_cell_53257 ( .a(n_9775), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q), .o(TIMEBOOST_net_16846) );
na02f02 TIMEBOOST_cell_69853 ( .a(TIMEBOOST_net_22134), .b(FE_OFN2129_n_16720), .o(TIMEBOOST_net_13222) );
in01m08 FE_RC_1041_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__531), .o(FE_RN_720_0) );
ao22f01 FE_RC_1043_0 ( .a(FE_RN_720_0), .b(FE_OFN1581_n_12306), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q), .d(FE_OFN1759_n_10780), .o(n_12721) );
in01m10 FE_RC_1044_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q), .o(FE_RN_722_0) );
in01f01 FE_RC_1045_0 ( .a(FE_OFN1559_n_12042), .o(FE_RN_723_0) );
na02s01 TIMEBOOST_cell_64074 ( .a(wishbone_slave_unit_fifos_outGreyCount_2_), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(TIMEBOOST_net_21023) );
in01s01 FE_RC_1048_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q), .o(FE_RN_725_0) );
in01f02 FE_RC_1049_0 ( .a(FE_OFN1556_n_12042), .o(FE_RN_726_0) );
na03f02 TIMEBOOST_cell_33523 ( .a(TIMEBOOST_net_8787), .b(FE_OFN1163_n_5615), .c(g62075_sb), .o(n_5636) );
na03m02 TIMEBOOST_cell_69100 ( .a(FE_OFN652_n_4508), .b(g65342_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q), .o(TIMEBOOST_net_21758) );
na02m02 TIMEBOOST_cell_44441 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q), .b(FE_OFN577_n_9902), .o(TIMEBOOST_net_13115) );
in01s01 FE_RC_1052_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q), .o(FE_RN_728_0) );
in01f01 FE_RC_1053_0 ( .a(FE_OFN1556_n_12042), .o(FE_RN_729_0) );
na03m02 TIMEBOOST_cell_68826 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q), .b(g65096_sb), .c(g65096_db), .o(TIMEBOOST_net_21621) );
in01s01 TIMEBOOST_cell_63591 ( .a(TIMEBOOST_net_20771), .o(TIMEBOOST_net_20770) );
na03f02 FE_RC_1056_0 ( .a(n_14535), .b(n_14407), .c(n_14497), .o(n_14579) );
na03f02 FE_RC_1057_0 ( .a(n_14549), .b(n_14253), .c(n_14440), .o(n_14594) );
in01f40 FE_RC_105_0 ( .a(wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_), .o(FE_RN_60_0) );
ao22f02 FE_RC_1060_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN1511_n_15587), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q), .d(FE_OFN1725_n_16891), .o(n_16845) );
ao22f02 FE_RC_1061_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q), .b(FE_OCP_RBN1969_FE_OFN1532_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q), .d(n_10195), .o(n_10078) );
in01f40 FE_RC_1062_0 ( .a(parchk_pci_ad_out_in_1174), .o(FE_RN_731_0) );
in01f40 FE_RC_1063_0 ( .a(parchk_pci_ad_out_in_1173), .o(FE_RN_732_0) );
in01f04 FE_RC_1066_0 ( .a(n_13415), .o(FE_RN_734_0) );
in01f02 FE_RC_1067_0 ( .a(n_7312), .o(FE_RN_735_0) );
na03f02 TIMEBOOST_cell_70054 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN707_n_8119), .c(n_2210), .o(TIMEBOOST_net_22235) );
na03f02 TIMEBOOST_cell_34952 ( .a(TIMEBOOST_net_9455), .b(FE_OFN1414_n_8567), .c(g57088_sb), .o(n_11653) );
in01f40 FE_RC_106_0 ( .a(wishbone_slave_unit_fifos_outGreyCount_1_), .o(FE_RN_61_0) );
in01f02 FE_RC_1070_0 ( .a(n_3070), .o(FE_RN_737_0) );
in01f02 FE_RC_1071_0 ( .a(n_3292), .o(FE_RN_738_0) );
no02f02 FE_RC_1072_0 ( .a(FE_RN_737_0), .b(FE_RN_738_0), .o(FE_RN_739_0) );
na02m02 TIMEBOOST_cell_69385 ( .a(TIMEBOOST_net_21900), .b(g64757_sb), .o(TIMEBOOST_net_12685) );
in01m02 FE_RC_1074_0 ( .a(n_2284), .o(FE_RN_740_0) );
in01m02 FE_RC_1075_0 ( .a(n_2137), .o(FE_RN_741_0) );
na04f02 FE_RC_1078_0 ( .a(n_11062), .b(n_11061), .c(n_11777), .d(n_11060), .o(n_12535) );
na04f02 FE_RC_1079_0 ( .a(n_11056), .b(n_11053), .c(n_11055), .d(n_11054), .o(n_12533) );
na03f04 TIMEBOOST_cell_71338 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_515), .c(n_2809), .o(TIMEBOOST_net_22877) );
na04f02 FE_RC_1080_0 ( .a(n_11140), .b(n_11136), .c(n_11139), .d(n_11137), .o(n_12554) );
na04f02 FE_RC_1081_0 ( .a(n_11039), .b(n_11773), .c(n_11040), .d(n_11041), .o(n_12530) );
na02f02 TIMEBOOST_cell_30711 ( .a(n_9019), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q), .o(TIMEBOOST_net_9460) );
in01f02 FE_RC_1083_0 ( .a(n_10688), .o(FE_RN_743_0) );
in01f02 FE_RC_1084_0 ( .a(FE_RN_179_0), .o(FE_RN_744_0) );
no02f02 FE_RC_1085_0 ( .a(FE_RN_744_0), .b(FE_RN_743_0), .o(FE_RN_745_0) );
na02f02 FE_RC_1086_0 ( .a(FE_RN_745_0), .b(n_12579), .o(n_12841) );
ao22f02 FE_RC_1087_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q), .b(FE_OFN1511_n_15587), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q), .d(FE_OFN1725_n_16891), .o(n_16985) );
in01f02 FE_RC_1088_0 ( .a(n_10851), .o(FE_RN_746_0) );
in01f02 FE_RC_1089_0 ( .a(FE_RN_465_0), .o(FE_RN_747_0) );
no02f02 FE_RC_1090_0 ( .a(FE_RN_746_0), .b(FE_RN_747_0), .o(FE_RN_748_0) );
na02f02 FE_RC_1091_0 ( .a(n_12559), .b(FE_RN_748_0), .o(n_12821) );
na02s01 g65784_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q), .b(FE_OFN941_n_2047), .o(g65784_db) );
in01s01 FE_RC_1093_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q), .o(FE_RN_749_0) );
in01f01 FE_RC_1094_0 ( .a(FE_OFN1720_n_16891), .o(FE_RN_750_0) );
no02f02 FE_RC_1095_0 ( .a(FE_RN_749_0), .b(FE_RN_750_0), .o(FE_RN_751_0) );
no02f02 FE_RC_1096_0 ( .a(n_15592), .b(FE_RN_751_0), .o(n_15593) );
ao22f02 FE_RC_1097_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q), .b(FE_OFN2147_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q), .d(FE_OFN1523_n_10892), .o(n_10596) );
na03f02 FE_RC_1098_0 ( .a(n_16260), .b(n_16255), .c(n_16258), .o(n_16261) );
ao22f02 FE_RC_1099_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q), .b(FE_OCP_RBN1968_FE_OFN1532_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q), .d(n_10185), .o(n_10188) );
in01f40 FE_RC_109_0 ( .a(wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_), .o(FE_RN_63_0) );
in01f02 FE_RC_10_0 ( .a(n_16021), .o(FE_RN_6_0) );
ao22f02 FE_RC_1100_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN1511_n_15587), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q), .d(FE_OFN1725_n_16891), .o(n_9982) );
ao22f02 FE_RC_1101_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q), .b(FE_OCP_RBN1968_FE_OFN1532_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q), .d(n_10185), .o(n_10026) );
in01s01 TIMEBOOST_cell_45941 ( .a(wbu_sel_in_314), .o(TIMEBOOST_net_13902) );
ao22f02 FE_RC_1103_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q), .b(FE_OFN2147_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q), .d(FE_OFN1523_n_10892), .o(n_10173) );
ao22f02 FE_RC_1104_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q), .b(FE_OFN2147_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q), .d(FE_OFN1523_n_10892), .o(n_10877) );
ao22f02 FE_RC_1105_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q), .d(FE_OFN1547_n_10566), .o(n_9979) );
in01f08 FE_RC_1106_0 ( .a(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(FE_RN_752_0) );
in01f08 FE_RC_1107_0 ( .a(n_15859), .o(FE_RN_753_0) );
na02f10 FE_RC_1108_0 ( .a(FE_RN_752_0), .b(FE_RN_753_0), .o(FE_OFN997_n_15978) );
no02f02 FE_RC_1109_0 ( .a(n_15859), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(TIMEBOOST_net_5257) );
in01f40 FE_RC_110_0 ( .a(wishbone_slave_unit_fifos_outGreyCount_0_), .o(FE_RN_64_0) );
in01f20 FE_RC_1110_0 ( .a(wishbone_slave_unit_pci_initiator_if_err_recovery), .o(FE_RN_754_0) );
no03f20 FE_RC_1111_0 ( .a(FE_RN_754_0), .b(n_15859), .c(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_15979) );
no02m10 FE_RC_1112_0 ( .a(wbu_pciif_devsel_reg_in), .b(n_16763), .o(n_15798) );
na02f08 FE_RC_1114_0 ( .a(g75418_da), .b(g75418_db), .o(n_16974) );
in01f04 FE_RC_1115_0 ( .a(g75418_db), .o(FE_RN_755_0) );
in01f06 FE_RC_1116_0 ( .a(g75418_da), .o(FE_RN_756_0) );
no02f10 FE_RC_1117_0 ( .a(FE_RN_756_0), .b(FE_RN_755_0), .o(n_16205) );
in01f08 FE_RC_1118_0 ( .a(n_16966), .o(n_16967) );
na02s02 TIMEBOOST_cell_49474 ( .a(TIMEBOOST_net_14954), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9499) );
na02f02 TIMEBOOST_cell_51328 ( .a(TIMEBOOST_net_15881), .b(g62500_sb), .o(n_6582) );
in01f02 FE_RC_1123_0 ( .a(n_16974), .o(FE_RN_758_0) );
na02f02 FE_RC_1124_0 ( .a(FE_OCP_RBN2016_n_16970), .b(n_16967), .o(FE_RN_759_0) );
no02f08 FE_RC_1125_0 ( .a(FE_RN_759_0), .b(FE_RN_758_0), .o(n_13901) );
na02m08 TIMEBOOST_cell_48227 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q), .b(FE_OFN1626_n_4438), .o(TIMEBOOST_net_14331) );
in01f20 FE_RC_1130_0 ( .a(n_16516), .o(FE_RN_764_0) );
na04f02 FE_RC_1135_0 ( .a(n_13930), .b(n_14499), .c(n_14536), .d(n_13849), .o(n_14580) );
na03f02 TIMEBOOST_cell_34882 ( .a(TIMEBOOST_net_9330), .b(FE_OFN1387_n_8567), .c(g57189_sb), .o(n_11564) );
in01f02 FE_RC_1138_0 ( .a(n_13854), .o(FE_RN_767_0) );
in01s01 FE_RC_1139_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q), .o(FE_RN_768_0) );
in01f08 FE_RC_113_0 ( .a(n_15401), .o(FE_RN_66_0) );
in01f02 FE_RC_1140_0 ( .a(FE_OCP_RBN1996_n_13971), .o(FE_RN_769_0) );
na03f02 TIMEBOOST_cell_34975 ( .a(TIMEBOOST_net_9566), .b(FE_OFN1370_n_8567), .c(g57564_sb), .o(n_10297) );
na03f10 TIMEBOOST_cell_64289 ( .a(n_16499), .b(n_16501), .c(n_16516), .o(n_16503) );
na04f02 FE_RC_1143_0 ( .a(n_11781), .b(n_11071), .c(n_11070), .d(n_11069), .o(n_12538) );
ao22f02 FE_RC_1144_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN1462_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q), .d(FE_OFN1457_n_11138), .o(n_17017) );
ao22f02 FE_RC_1145_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q), .b(FE_OCP_RBN2010_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q), .d(FE_OFN1465_n_10789), .o(n_11093) );
na04f03 FE_RC_1146_0 ( .a(n_12959), .b(n_12897), .c(n_12896), .d(n_12789), .o(n_13135) );
na03f20 FE_RC_1149_0 ( .a(n_16434), .b(n_16462), .c(n_16265), .o(n_16499) );
in01f08 FE_RC_114_0 ( .a(n_16798), .o(FE_RN_67_0) );
in01f20 FE_RC_1153_0 ( .a(n_16264), .o(n_15823) );
no02f40 FE_RC_1155_0 ( .a(FE_OCP_RBN2270_g75061_p), .b(n_16264), .o(FE_RN_772_0) );
na02f20 FE_RC_1156_0 ( .a(n_16599), .b(FE_RN_772_0), .o(n_16980) );
in01f02 FE_RC_1157_0 ( .a(n_16154), .o(FE_RN_773_0) );
in01f02 FE_RC_1158_0 ( .a(n_16153), .o(FE_RN_774_0) );
no02f04 FE_RC_1159_0 ( .a(FE_RN_774_0), .b(FE_RN_773_0), .o(FE_RN_775_0) );
na02f06 FE_RC_1160_0 ( .a(FE_RN_775_0), .b(n_16980), .o(n_16156) );
in01f06 FE_RC_1161_0 ( .a(FE_RN_776_0), .o(n_3421) );
na02f08 FE_RC_1162_0 ( .a(FE_OCP_RBN2238_g74749_p), .b(n_3310), .o(FE_RN_776_0) );
in01f01 FE_RC_1166_0 ( .a(n_16966), .o(FE_RN_778_0) );
no02f04 FE_RC_1167_0 ( .a(FE_RN_778_0), .b(FE_OCP_RBN2279_n_16974), .o(FE_RN_779_0) );
na02f08 FE_RC_1168_0 ( .a(FE_RN_779_0), .b(FE_OCP_RBN2017_n_16970), .o(FE_OFN1772_n_13800) );
na02f04 FE_RC_1169_0 ( .a(FE_OCP_RBN2019_n_16970), .b(n_16966), .o(FE_RN_780_0) );
na03f02 TIMEBOOST_cell_68718 ( .a(TIMEBOOST_net_20217), .b(FE_OFN916_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q), .o(TIMEBOOST_net_21567) );
no02f10 FE_RC_1170_0 ( .a(FE_RN_780_0), .b(FE_OCP_RBN2278_n_16974), .o(FE_OFN1774_n_13800) );
in01f08 FE_RC_117_0 ( .a(pci_target_unit_pci_target_sm_rd_from_fifo), .o(FE_RN_69_0) );
in01f08 FE_RC_118_0 ( .a(pci_target_unit_pci_target_sm_same_read_reg), .o(FE_RN_70_0) );
in01f02 FE_RC_1194_0 ( .a(FE_RN_8_0), .o(FE_RN_795_0) );
no02f02 FE_RC_1195_0 ( .a(n_15919), .b(FE_RN_795_0), .o(n_15917) );
in01f04 FE_RC_1196_0 ( .a(n_16075), .o(n_16076) );
in01f02 FE_RC_1197_0 ( .a(n_16075), .o(FE_RN_796_0) );
na02f04 FE_RC_1198_0 ( .a(FE_RN_796_0), .b(n_16444), .o(n_15581) );
in01f40 FE_RC_1199_0 ( .a(parchk_pci_ad_out_in), .o(FE_RN_797_0) );
no02f10 FE_RC_119_0 ( .a(FE_RN_69_0), .b(FE_RN_70_0), .o(FE_RN_71_0) );
in01f02 FE_RC_11_0 ( .a(n_16914), .o(FE_RN_7_0) );
in01f40 FE_RC_1200_0 ( .a(parchk_pci_ad_out_in_1168), .o(FE_RN_798_0) );
na03f02 TIMEBOOST_cell_66225 ( .a(TIMEBOOST_net_13237), .b(FE_OFN1244_n_4092), .c(g62514_sb), .o(n_6550) );
na02f02 TIMEBOOST_cell_39380 ( .a(TIMEBOOST_net_7255), .b(FE_OFN1092_g64577_p), .o(TIMEBOOST_net_11302) );
in01s01 FE_RC_1203_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q), .o(FE_RN_800_0) );
no02f04 FE_RC_1204_0 ( .a(FE_OCPN1856_FE_OFN1774_n_13800), .b(FE_RN_800_0), .o(FE_RN_801_0) );
in01f02 FE_RC_1205_0 ( .a(FE_RN_802_0), .o(g53187_p) );
ao12f02 FE_RC_1206_0 ( .a(FE_RN_801_0), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q), .c(FE_OFN1771_n_14054), .o(FE_RN_802_0) );
na03m02 TIMEBOOST_cell_72517 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(g64199_sb), .c(g64199_db), .o(n_3970) );
na04f04 TIMEBOOST_cell_67626 ( .a(n_3786), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q), .c(FE_OFN1261_n_4143), .d(g62536_sb), .o(n_6498) );
na02f01 TIMEBOOST_cell_53380 ( .a(TIMEBOOST_net_16907), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_14523) );
na02s02 TIMEBOOST_cell_48822 ( .a(TIMEBOOST_net_14628), .b(g58169_sb), .o(TIMEBOOST_net_12791) );
in01f02 FE_RC_1211_0 ( .a(n_14963), .o(FE_RN_805_0) );
in01s01 FE_RC_1212_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q), .o(FE_RN_806_0) );
in01f02 FE_RC_1213_0 ( .a(FE_OCP_RBN1985_FE_OFN1591_n_13741), .o(FE_RN_807_0) );
na03f02 TIMEBOOST_cell_73346 ( .a(n_3815), .b(g63139_sb), .c(TIMEBOOST_net_6490), .o(n_4970) );
na02m01 TIMEBOOST_cell_62830 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q), .o(TIMEBOOST_net_20362) );
na03f02 TIMEBOOST_cell_34811 ( .a(TIMEBOOST_net_9391), .b(FE_OFN1388_n_8567), .c(g57576_sb), .o(n_11175) );
na02s01 TIMEBOOST_cell_49078 ( .a(TIMEBOOST_net_14756), .b(g65892_sb), .o(n_2592) );
na04f03 FE_RC_1219_0 ( .a(n_13050), .b(n_12886), .c(n_12887), .d(n_12786), .o(n_13133) );
in01m10 FE_RC_121_0 ( .a(n_2629), .o(FE_RN_72_0) );
ao22f02 FE_RC_1220_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q), .b(FE_OFN1727_n_9975), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q), .d(FE_OCP_RBN2005_FE_RN_459_0), .o(n_9303) );
ao22f02 FE_RC_1221_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q), .b(FE_OFN2149_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q), .d(FE_OFN1522_n_10892), .o(n_17046) );
ao22f02 FE_RC_1222_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q), .b(FE_OFN2147_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q), .d(FE_OFN1523_n_10892), .o(n_10054) );
ao22f02 FE_RC_1223_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q), .b(FE_OFN2149_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q), .d(FE_OFN1522_n_10892), .o(n_10930) );
ao22f02 FE_RC_1224_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q), .b(FE_OFN1536_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q), .d(n_10141), .o(n_17045) );
na02f01 TIMEBOOST_cell_47758 ( .a(TIMEBOOST_net_14096), .b(FE_OFN903_n_4736), .o(TIMEBOOST_net_10318) );
ao22f10 FE_RC_1226_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_), .c(n_16175), .d(FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .o(n_16433) );
na02f08 FE_RC_1227_0 ( .a(FE_OCP_RBN1955_n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .o(FE_RN_809_0) );
in01f02 FE_RC_1229_0 ( .a(n_13856), .o(FE_RN_810_0) );
in01f08 FE_RC_122_0 ( .a(n_2623), .o(FE_RN_73_0) );
in01s01 FE_RC_1230_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q), .o(FE_RN_811_0) );
in01f02 FE_RC_1231_0 ( .a(FE_OCP_RBN1995_n_13971), .o(FE_RN_812_0) );
na02f01 TIMEBOOST_cell_18751 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_5739) );
na03f02 TIMEBOOST_cell_34954 ( .a(TIMEBOOST_net_9456), .b(FE_OFN1399_n_8567), .c(g57348_sb), .o(n_11402) );
in01f02 FE_RC_1234_0 ( .a(n_13990), .o(FE_RN_814_0) );
in01f02 FE_RC_1235_0 ( .a(n_13991), .o(FE_RN_815_0) );
no02f02 FE_RC_1236_0 ( .a(FE_RN_814_0), .b(FE_RN_815_0), .o(n_14283) );
in01f02 FE_RC_1237_0 ( .a(n_14197), .o(FE_RN_816_0) );
in01s01 FE_RC_1238_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q), .o(FE_RN_817_0) );
in01f02 FE_RC_1239_0 ( .a(FE_OFN1769_n_14054), .o(FE_RN_818_0) );
na03f02 TIMEBOOST_cell_34836 ( .a(TIMEBOOST_net_9426), .b(FE_OFN1386_n_8567), .c(g57358_sb), .o(n_11390) );
na03f02 TIMEBOOST_cell_73563 ( .a(TIMEBOOST_net_17082), .b(FE_OFN2063_n_6391), .c(g62550_sb), .o(n_6465) );
na02m02 g52458_u1 ( .a(wbs_adr_i_12_), .b(g52458_sb), .o(g52458_da) );
na02s02 TIMEBOOST_cell_49524 ( .a(TIMEBOOST_net_14979), .b(FE_OFN272_n_9828), .o(n_9410) );
na02f20 FE_RC_1243_0 ( .a(n_16501), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in_86), .o(FE_RN_820_0) );
in01f20 FE_RC_1244_0 ( .a(pci_target_unit_wishbone_master_burst_chopped_delayed), .o(FE_RN_821_0) );
no03f20 FE_RC_1245_0 ( .a(FE_RN_764_0), .b(FE_RN_820_0), .c(FE_RN_821_0), .o(FE_RN_822_0) );
na02f10 FE_RC_1246_0 ( .a(n_16499), .b(FE_RN_822_0), .o(n_16513) );
in01f02 FE_RC_1250_0 ( .a(FE_RN_824_0), .o(n_14054) );
na03f03 FE_RC_1251_0 ( .a(n_16974), .b(n_16966), .c(n_16970), .o(FE_RN_824_0) );
na02f02 TIMEBOOST_cell_30911 ( .a(n_9013), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q), .o(TIMEBOOST_net_9560) );
in01s01 TIMEBOOST_cell_67742 ( .a(TIMEBOOST_net_21168), .o(TIMEBOOST_net_21169) );
na03f02 TIMEBOOST_cell_34977 ( .a(TIMEBOOST_net_9555), .b(FE_OFN1421_n_8567), .c(g57220_sb), .o(n_11535) );
in01f02 FE_RC_1256_0 ( .a(n_13847), .o(FE_RN_827_0) );
in01s01 FE_RC_1257_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q), .o(FE_RN_828_0) );
in01s02 FE_RC_1258_0 ( .a(FE_OCP_RBN1996_n_13971), .o(FE_RN_829_0) );
na03f02 TIMEBOOST_cell_34961 ( .a(TIMEBOOST_net_9464), .b(FE_OFN1411_n_8567), .c(g57372_sb), .o(n_11377) );
na03f02 TIMEBOOST_cell_34956 ( .a(TIMEBOOST_net_9458), .b(FE_OFN1400_n_8567), .c(g57477_sb), .o(n_11260) );
in01f02 FE_RC_1261_0 ( .a(n_14099), .o(FE_RN_831_0) );
in01m10 FE_RC_1262_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q), .o(FE_RN_832_0) );
in01f02 FE_RC_1263_0 ( .a(FE_OCPN2218_n_13997), .o(FE_RN_833_0) );
na03f08 TIMEBOOST_cell_23953 ( .a(n_7321), .b(n_4875), .c(n_17030), .o(n_15188) );
in01f02 FE_RC_1266_0 ( .a(n_14507), .o(FE_RN_835_0) );
na04f02 FE_RC_1267_0 ( .a(n_16170), .b(n_13937), .c(n_13938), .d(FE_RN_835_0), .o(n_16173) );
na03f10 FE_RC_1268_0 ( .a(n_16392), .b(n_16391), .c(n_16393), .o(n_16394) );
na03f02 TIMEBOOST_cell_73585 ( .a(n_3357), .b(FE_OFN1700_n_5751), .c(TIMEBOOST_net_15708), .o(n_14847) );
na04f02 FE_RC_1270_0 ( .a(n_11101), .b(n_11099), .c(n_11102), .d(n_11100), .o(n_12546) );
na04f04 FE_RC_1271_0 ( .a(n_11819), .b(n_12248), .c(n_12246), .d(n_11960), .o(n_12814) );
ao22f02 FE_RC_1273_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q), .b(FE_OFN2137_n_15534), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q), .d(FE_OFN2144_n_16992), .o(n_16984) );
ao22f02 FE_RC_1274_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q), .b(FE_OFN2149_n_10595), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q), .d(FE_OFN1522_n_10892), .o(n_10524) );
ao22f02 FE_RC_1275_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q), .b(FE_OFN2216_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q), .d(n_11728), .o(n_11733) );
ao22f02 FE_RC_1276_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q), .d(FE_OFN1547_n_10566), .o(n_9311) );
ao22f02 FE_RC_1277_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q), .b(FE_OFN1535_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q), .d(n_11728), .o(n_10947) );
ao22f02 FE_RC_1278_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q), .b(FE_OFN1493_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q), .d(FE_OFN1546_n_10566), .o(n_10903) );
ao22f02 FE_RC_1279_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q), .b(FE_OFN1478_n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q), .d(FE_OFN2193_n_9163), .o(n_11118) );
na03f02 FE_RC_1280_0 ( .a(n_13051), .b(FE_RN_113_0), .c(n_12787), .o(n_13134) );
ao22f02 FE_RC_1281_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q), .b(FE_OFN2131_n_10588), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q), .d(FE_OFN1528_n_10853), .o(n_10533) );
ao22f02 FE_RC_1282_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q), .b(FE_OFN1508_n_15587), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q), .d(FE_OFN1720_n_16891), .o(n_9988) );
ao22f02 FE_RC_1283_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q), .b(FE_OFN2216_n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q), .d(n_11728), .o(n_11726) );
ao22f02 FE_RC_1284_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q), .b(FE_OFN1727_n_9975), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q), .d(FE_OCP_RBN1932_FE_OFN1515_n_10538), .o(n_17044) );
ao22f02 FE_RC_1285_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q), .b(FE_OFN1493_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q), .d(FE_OFN1546_n_10566), .o(n_10702) );
ao22f02 FE_RC_1286_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q), .b(n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q), .d(FE_OFN2194_n_9163), .o(n_11091) );
ao22f02 FE_RC_1287_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q), .b(FE_OCP_RBN2010_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q), .d(FE_OFN1465_n_10789), .o(n_11059) );
ao22f02 FE_RC_1288_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q), .b(FE_OFN1479_n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q), .d(FE_OFN2194_n_9163), .o(n_11073) );
in01f02 FE_RC_1289_0 ( .a(n_16358), .o(FE_RN_836_0) );
in01f08 FE_RC_1291_0 ( .a(FE_RN_0_0), .o(FE_RN_837_0) );
in01f03 FE_RC_1293_0 ( .a(n_16513), .o(FE_RN_839_0) );
na02s01 TIMEBOOST_cell_48038 ( .a(TIMEBOOST_net_14236), .b(g58155_db), .o(TIMEBOOST_net_9509) );
na02m04 TIMEBOOST_cell_38212 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q), .b(g65339_sb), .o(TIMEBOOST_net_10718) );
na03f02 TIMEBOOST_cell_34791 ( .a(TIMEBOOST_net_9544), .b(FE_OFN1391_n_8567), .c(g57527_sb), .o(n_11214) );
na03f02 TIMEBOOST_cell_34710 ( .a(TIMEBOOST_net_8560), .b(FE_OFN2136_n_13124), .c(g54364_sb), .o(n_13078) );
in01f02 FE_RC_1299_0 ( .a(n_14111), .o(FE_RN_843_0) );
no02f04 FE_RC_12_0 ( .a(FE_RN_7_0), .b(FE_RN_6_0), .o(FE_RN_8_0) );
in01m10 FE_RC_1300_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q), .o(FE_RN_844_0) );
in01f02 FE_RC_1301_0 ( .a(FE_OFN1602_n_13995), .o(FE_RN_845_0) );
na03f02 FE_RC_1304_0 ( .a(FE_RN_847_0), .b(n_14515), .c(n_14433), .o(n_14591) );
ao22f02 FE_RC_1305_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q), .d(FE_OFN1547_n_10566), .o(n_10023) );
ao22f02 FE_RC_1306_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q), .b(FE_OFN1489_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q), .d(FE_OFN1548_n_10566), .o(n_9287) );
ao22f02 FE_RC_1307_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q), .d(FE_OFN1547_n_10566), .o(n_9297) );
ao22f02 FE_RC_1308_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q), .b(FE_OCP_RBN2011_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q), .d(FE_OFN1467_n_10789), .o(n_10791) );
na03f10 FE_RC_1309_0 ( .a(FE_OFN996_n_15366), .b(n_16049), .c(n_16046), .o(n_16310) );
na03m02 TIMEBOOST_cell_73201 ( .a(TIMEBOOST_net_16333), .b(TIMEBOOST_net_12902), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q), .o(TIMEBOOST_net_22317) );
ao22f02 FE_RC_1310_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q), .b(FE_OFN2146_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q), .d(FE_OFN1547_n_10566), .o(n_9319) );
ao22f02 FE_RC_1311_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q), .b(FE_OCP_RBN2009_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q), .d(FE_OFN1466_n_10789), .o(n_11137) );
na04f04 FE_RC_1312_0 ( .a(n_12052), .b(n_12053), .c(n_12055), .d(n_12054), .o(n_12819) );
in01f02 FE_RC_1335_0 ( .a(n_16403), .o(FE_RN_862_0) );
in01f02 FE_RC_1336_0 ( .a(n_16406), .o(FE_RN_863_0) );
na03f02 FE_RC_1338_0 ( .a(n_13059), .b(FE_RN_107_0), .c(n_12799), .o(n_13141) );
in01f04 FE_RC_1364_0 ( .a(n_16547), .o(FE_RN_880_0) );
in01f04 FE_RC_1365_0 ( .a(n_16550), .o(FE_RN_881_0) );
no02f08 FE_RC_1366_0 ( .a(FE_RN_880_0), .b(FE_RN_881_0), .o(n_16552) );
na04f02 FE_RC_1367_0 ( .a(n_13065), .b(n_12932), .c(n_12931), .d(n_12801), .o(n_13142) );
na04f03 FE_RC_1368_0 ( .a(n_13049), .b(n_12884), .c(n_12883), .d(n_12785), .o(n_13132) );
na03f02 FE_RC_1369_0 ( .a(n_13120), .b(n_12928), .c(FE_RN_236_0), .o(n_13323) );
in01s01 TIMEBOOST_cell_45939 ( .a(TIMEBOOST_net_13900), .o(TIMEBOOST_net_5291) );
na02s01 TIMEBOOST_cell_44443 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q), .b(FE_OFN542_n_9690), .o(TIMEBOOST_net_13116) );
no02f08 FE_RC_1372_0 ( .a(n_3448), .b(n_3320), .o(FE_RN_882_0) );
na02s02 TIMEBOOST_cell_54174 ( .a(TIMEBOOST_net_17304), .b(g57925_sb), .o(TIMEBOOST_net_14951) );
no02f20 FE_RC_1375_0 ( .a(FE_RN_428_0), .b(FE_RN_430_0), .o(FE_OFN1026_n_16760) );
ao22f02 FE_RC_1377_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q), .b(FE_OFN1493_n_9320), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q), .d(FE_OFN1546_n_10566), .o(n_10741) );
ao22f02 FE_RC_1378_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q), .b(FE_OFN2130_n_10588), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q), .d(FE_OFN1530_n_10853), .o(n_10951) );
na03f02 TIMEBOOST_cell_72937 ( .a(pci_target_unit_del_sync_addr_in_221), .b(g65248_sb), .c(TIMEBOOST_net_7147), .o(n_2634) );
in01f20 FE_RC_137_0 ( .a(configuration_sync_command_bit1), .o(FE_RN_81_0) );
no02f10 FE_RC_1383_0 ( .a(n_16433), .b(FE_OCP_RBN2271_g75061_p), .o(n_16434) );
na02f08 FE_RC_1384_0 ( .a(FE_RN_809_0), .b(g75413_db), .o(n_16966) );
na02f02 FE_RC_1385_0 ( .a(FE_RN_809_0), .b(g75413_db), .o(n_14939) );
na02f02 TIMEBOOST_cell_54712 ( .a(TIMEBOOST_net_17573), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_15371) );
na02f02 FE_RC_1388_0 ( .a(n_13891), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q), .o(FE_RN_887_0) );
in01s01 FE_RC_1389_0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q), .o(FE_RN_888_0) );
in01m20 FE_RC_138_0 ( .a(conf_pci_init_complete_out), .o(FE_RN_82_0) );
oa12f02 FE_RC_1390_0 ( .a(FE_RN_887_0), .b(FE_RN_888_0), .c(FE_OCP_RBN1964_FE_OFN1591_n_13741), .o(g53206_p) );
na02f02 TIMEBOOST_cell_68839 ( .a(TIMEBOOST_net_21627), .b(g64995_sb), .o(TIMEBOOST_net_20962) );
na02m08 TIMEBOOST_cell_69690 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q), .b(FE_OFN1680_n_4655), .o(TIMEBOOST_net_22053) );
no02f02 FE_RC_1393_0 ( .a(FE_RN_890_0), .b(n_14268), .o(n_14556) );
ao22f02 FE_RC_1394_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q), .b(FE_OFN1478_n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q), .d(FE_OFN2193_n_9163), .o(n_11104) );
ao22f02 FE_RC_1395_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q), .b(n_15566), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q), .d(n_15558), .o(n_9328) );
ao22f02 FE_RC_1396_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q), .b(n_15566), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q), .d(FE_OFN1499_n_15558), .o(n_10002) );
ao22f02 FE_RC_1397_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q), .b(FE_OFN2137_n_15534), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q), .d(FE_OCPN1873_FE_OFN474_n_16992), .o(n_10755) );
ao22f04 FE_RC_1398_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q), .b(FE_OFN1485_n_15534), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q), .d(FE_OCPN1888_FE_OFN473_n_16992), .o(n_10758) );
ao22f02 FE_RC_1399_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q), .b(FE_OFN1433_n_16779), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q), .d(FE_OFN1445_n_11125), .o(n_11051) );
no02f10 FE_RC_139_0 ( .a(FE_RN_81_0), .b(FE_RN_82_0), .o(FE_RN_83_0) );
ao22f02 FE_RC_1400_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q), .b(FE_OFN1432_n_16779), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q), .d(FE_OFN1445_n_11125), .o(n_11113) );
ao22f02 FE_RC_1401_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q), .b(FE_OFN2208_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q), .d(FE_OFN1455_n_11138), .o(n_11777) );
ao22f02 FE_RC_1402_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q), .b(FE_OFN1462_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q), .d(FE_OFN1457_n_11138), .o(n_11107) );
na04f04 TIMEBOOST_cell_24235 ( .a(n_9547), .b(g57388_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q), .d(FE_OFN1424_n_8567), .o(n_11355) );
na02s02 TIMEBOOST_cell_50057 ( .a(g58417_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q), .o(TIMEBOOST_net_15246) );
na04s02 TIMEBOOST_cell_46578 ( .a(TIMEBOOST_net_10786), .b(g65834_sb), .c(g61899_sb), .d(g61899_db), .o(n_8027) );
na03f02 TIMEBOOST_cell_34958 ( .a(TIMEBOOST_net_9527), .b(FE_OFN1382_n_8567), .c(g57578_sb), .o(n_10292) );
no02f02 FE_RC_1407_0 ( .a(n_14505), .b(FE_RN_893_0), .o(n_14539) );
na04f02 FE_RC_1408_0 ( .a(n_14275), .b(n_13980), .c(n_13859), .d(n_14560), .o(n_14605) );
na02s01 TIMEBOOST_cell_47515 ( .a(parchk_pci_ad_reg_in_1223), .b(g67049_db), .o(TIMEBOOST_net_13975) );
ao22f02 FE_RC_1410_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q), .b(FE_OFN1460_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q), .d(FE_OFN1456_n_11138), .o(n_11058) );
na03f02 FE_RC_1411_0 ( .a(FE_RN_863_0), .b(n_13067), .c(FE_RN_862_0), .o(n_13408) );
ao22f02 FE_RC_1412_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN1731_n_9975), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q), .d(FE_OCP_RBN2006_FE_RN_459_0), .o(n_10530) );
ao22f02 FE_RC_1413_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q), .b(n_15566), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q), .d(FE_OFN1501_n_15558), .o(n_9265) );
ao22f02 FE_RC_1414_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q), .b(FE_OCPN1884_n_15566), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q), .d(FE_OFN1498_n_15558), .o(n_10179) );
ao22f02 FE_RC_1415_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q), .b(FE_OFN2208_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q), .d(FE_OFN1455_n_11138), .o(n_11048) );
ao22f02 FE_RC_1416_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q), .b(FE_OCP_RBN2009_n_16698), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q), .d(FE_OFN1466_n_10789), .o(n_11106) );
ao22f02 FE_RC_1417_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q), .b(FE_OFN1484_n_15534), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q), .d(n_16992), .o(n_16834) );
ao22f02 FE_RC_1418_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN1462_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q), .d(FE_OFN1457_n_11138), .o(n_11139) );
ao22f02 FE_RC_1419_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q), .b(FE_OFN2208_n_11795), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q), .d(FE_OFN1455_n_11138), .o(n_11796) );
in01f02 FE_RC_1420_0 ( .a(n_15917), .o(FE_RN_894_0) );
no02f06 FE_RC_1421_0 ( .a(FE_RN_894_0), .b(FE_RN_390_0), .o(FE_RN_895_0) );
na03f02 TIMEBOOST_cell_73132 ( .a(TIMEBOOST_net_22142), .b(g64230_sb), .c(FE_OFN2104_g64577_p), .o(TIMEBOOST_net_22509) );
in01f06 FE_RC_1423_0 ( .a(n_16523), .o(FE_RN_896_0) );
oa22f08 FE_RC_1424_0 ( .a(n_16523), .b(FE_RN_493_0), .c(FE_RN_896_0), .d(FE_RN_491_0), .o(n_16075) );
in01f08 FE_RC_1425_0 ( .a(FE_RN_15_0), .o(FE_RN_897_0) );
in01f06 FE_RC_1426_0 ( .a(FE_RN_899_0), .o(FE_RN_898_0) );
no02f10 FE_RC_1427_0 ( .a(FE_RN_897_0), .b(FE_RN_898_0), .o(n_14971) );
na02f08 FE_RC_1428_0 ( .a(n_15915), .b(n_16524), .o(FE_RN_899_0) );
in01f04 FE_RC_1429_0 ( .a(FE_RN_15_0), .o(FE_RN_900_0) );
in01f10 FE_RC_1430_0 ( .a(n_135), .o(FE_RN_901_0) );
no02f08 FE_RC_1431_0 ( .a(FE_RN_900_0), .b(FE_RN_901_0), .o(FE_RN_902_0) );
na02f08 FE_RC_1432_0 ( .a(FE_RN_899_0), .b(FE_RN_902_0), .o(n_16564) );
ao22f02 FE_RC_1433_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q), .b(n_10143), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q), .d(n_11728), .o(n_10931) );
na02f02 FE_RC_1436_0 ( .a(wbm_dat_o_22_), .b(n_14800), .o(FE_RN_904_0) );
in01s01 FE_RC_1437_0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71), .o(FE_RN_905_0) );
oa12f02 FE_RC_1438_0 ( .a(FE_RN_904_0), .b(FE_RN_905_0), .c(n_14725), .o(FE_RN_906_0) );
in01f02 FE_RC_1439_0 ( .a(FE_RN_907_0), .o(n_16304) );
ao22f02 FE_RC_1440_0 ( .a(n_16300), .b(FE_RN_906_0), .c(wbm_dat_o_22_), .d(FE_OFN2164_n_16301), .o(FE_RN_907_0) );
na02f01 TIMEBOOST_cell_70324 ( .a(TIMEBOOST_net_8808), .b(FE_OFN1095_g64577_p), .o(TIMEBOOST_net_22370) );
in01f02 FE_RC_1443_0 ( .a(n_12753), .o(FE_RN_909_0) );
in01f02 FE_RC_1444_0 ( .a(FE_RN_908_0), .o(FE_RN_910_0) );
in01f02 FE_RC_1447_0 ( .a(n_16022), .o(FE_RN_911_0) );
no02f02 FE_RC_1448_0 ( .a(n_15919), .b(FE_RN_911_0), .o(n_15914) );
in01f04 FE_RC_1449_0 ( .a(FE_RN_912_0), .o(n_16313) );
na02f06 FE_RC_1450_0 ( .a(n_16547), .b(n_16554), .o(FE_RN_912_0) );
in01f02 FE_RC_1451_0 ( .a(n_12257), .o(FE_RN_913_0) );
in01f02 FE_RC_1452_0 ( .a(n_11975), .o(FE_RN_914_0) );
no02f02 FE_RC_1453_0 ( .a(FE_RN_913_0), .b(FE_RN_914_0), .o(n_16411) );
in01f02 FE_RC_1454_0 ( .a(n_12031), .o(FE_RN_915_0) );
no02f02 FE_RC_1455_0 ( .a(FE_RN_25_0), .b(FE_RN_915_0), .o(FE_RN_26_0) );
in01f02 FE_RC_1456_0 ( .a(n_15935), .o(FE_RN_916_0) );
in01f02 FE_RC_1457_0 ( .a(n_15937), .o(FE_RN_917_0) );
ao22f02 FE_RC_1459_0 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q), .b(FE_OFN1479_n_16637), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q), .d(FE_OFN2195_n_9163), .o(n_11077) );
na03m02 TIMEBOOST_cell_73202 ( .a(TIMEBOOST_net_14598), .b(g65843_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q), .o(TIMEBOOST_net_22327) );
na04f04 FE_RC_1461_0 ( .a(n_15940), .b(FE_RN_917_0), .c(FE_RN_916_0), .d(n_15941), .o(n_15942) );
na04f04 FE_RC_1462_0 ( .a(n_11914), .b(n_11915), .c(n_11913), .d(n_11912), .o(n_12810) );
na03f02 FE_RC_148_0 ( .a(n_14557), .b(n_14456), .c(n_14269), .o(n_14602) );
in01f02 FE_RC_149_0 ( .a(n_10650), .o(FE_RN_87_0) );
in01f02 FE_RC_150_0 ( .a(n_10647), .o(FE_RN_88_0) );
no02f02 FE_RC_151_0 ( .a(FE_RN_87_0), .b(FE_RN_88_0), .o(FE_RN_89_0) );
in01f02 FE_RC_153_0 ( .a(n_10179), .o(FE_RN_90_0) );
in01f02 FE_RC_154_0 ( .a(n_10754), .o(FE_RN_91_0) );
no02f02 FE_RC_155_0 ( .a(FE_RN_90_0), .b(FE_RN_91_0), .o(FE_RN_92_0) );
na03f02 TIMEBOOST_cell_34857 ( .a(TIMEBOOST_net_9322), .b(FE_OFN1391_n_8567), .c(g57201_sb), .o(n_10445) );
in01f02 FE_RC_157_0 ( .a(n_10750), .o(FE_RN_93_0) );
in01f02 FE_RC_158_0 ( .a(n_10747), .o(FE_RN_94_0) );
no02f02 FE_RC_159_0 ( .a(FE_RN_93_0), .b(FE_RN_94_0), .o(FE_RN_95_0) );
in01f08 FE_RC_15_0 ( .a(n_16159), .o(FE_RN_9_0) );
na03f02 FE_RC_160_0 ( .a(n_12585), .b(n_10744), .c(FE_RN_95_0), .o(n_12847) );
in01f02 FE_RC_161_0 ( .a(n_10774), .o(FE_RN_96_0) );
in01f02 FE_RC_162_0 ( .a(n_10771), .o(FE_RN_97_0) );
no02f02 FE_RC_163_0 ( .a(FE_RN_96_0), .b(FE_RN_97_0), .o(FE_RN_98_0) );
in01f10 TIMEBOOST_cell_17842 ( .a(TIMEBOOST_net_5253), .o(TIMEBOOST_net_5252) );
in01f02 FE_RC_165_0 ( .a(n_10544), .o(FE_RN_99_0) );
in01f02 FE_RC_166_0 ( .a(n_10541), .o(FE_RN_100_0) );
no02f02 FE_RC_167_0 ( .a(FE_RN_99_0), .b(FE_RN_100_0), .o(FE_RN_101_0) );
in01s01 TIMEBOOST_cell_63590 ( .a(TIMEBOOST_net_20770), .o(TIMEBOOST_net_20719) );
in01f04 FE_RC_169_0 ( .a(parchk_pci_cbe_reg_in_1236), .o(FE_RN_102_0) );
in01f08 FE_RC_170_0 ( .a(n_2071), .o(FE_RN_103_0) );
na03s04 TIMEBOOST_cell_72675 ( .a(TIMEBOOST_net_14266), .b(FE_OFN955_n_1699), .c(g65793_sb), .o(n_1593) );
na02f02 TIMEBOOST_cell_70709 ( .a(TIMEBOOST_net_22562), .b(g63084_sb), .o(n_5086) );
in01f02 FE_RC_173_0 ( .a(n_12922), .o(FE_RN_105_0) );
in01f02 FE_RC_174_0 ( .a(n_12923), .o(FE_RN_106_0) );
no02f02 FE_RC_175_0 ( .a(FE_RN_106_0), .b(FE_RN_105_0), .o(FE_RN_107_0) );
in01f02 FE_RC_178_0 ( .a(n_12949), .o(FE_RN_108_0) );
in01f02 FE_RC_179_0 ( .a(n_12950), .o(FE_RN_109_0) );
na03f02 TIMEBOOST_cell_66309 ( .a(TIMEBOOST_net_17055), .b(n_6232), .c(g62926_sb), .o(n_6029) );
no02f02 FE_RC_180_0 ( .a(FE_RN_109_0), .b(FE_RN_108_0), .o(FE_RN_110_0) );
na03f02 FE_RC_181_0 ( .a(FE_RN_110_0), .b(n_12809), .c(n_12964), .o(n_13144) );
in01f02 FE_RC_182_0 ( .a(n_12889), .o(FE_RN_111_0) );
in01f02 FE_RC_183_0 ( .a(n_12890), .o(FE_RN_112_0) );
no02f02 FE_RC_184_0 ( .a(FE_RN_112_0), .b(FE_RN_111_0), .o(FE_RN_113_0) );
in01f02 FE_RC_186_0 ( .a(n_12913), .o(FE_RN_114_0) );
in01f02 FE_RC_187_0 ( .a(n_12912), .o(FE_RN_115_0) );
no02f02 FE_RC_188_0 ( .a(FE_RN_115_0), .b(FE_RN_114_0), .o(FE_RN_116_0) );
na03f02 FE_RC_189_0 ( .a(n_12795), .b(FE_RN_116_0), .c(n_13118), .o(n_13320) );
in01s01 FE_RC_196_0 ( .a(n_16635), .o(FE_RN_120_0) );
in01s01 FE_RC_197_0 ( .a(n_1963), .o(FE_RN_121_0) );
no02s01 FE_RC_198_0 ( .a(FE_RN_121_0), .b(FE_RN_120_0), .o(FE_RN_122_0) );
na04f04 TIMEBOOST_cell_73188 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q), .c(FE_OFN1670_n_9477), .d(g58366_sb), .o(n_9013) );
in01f02 FE_RC_201_0 ( .a(n_13672), .o(FE_RN_124_0) );
na02s02 TIMEBOOST_cell_48011 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_14223) );
in01s01 TIMEBOOST_cell_45962 ( .a(TIMEBOOST_net_13922), .o(TIMEBOOST_net_13923) );
in01f02 FE_RC_205_0 ( .a(n_13651), .o(FE_RN_127_0) );
in01f02 FE_RC_209_0 ( .a(n_13661), .o(FE_RN_130_0) );
na03f04 TIMEBOOST_cell_70382 ( .a(n_2995), .b(n_4743), .c(n_2329), .o(TIMEBOOST_net_22399) );
in01s01 TIMEBOOST_cell_17889 ( .a(TIMEBOOST_net_5300), .o(wbs_dat_i_2_) );
na04f04 FE_RC_217_0 ( .a(n_14961), .b(n_14142), .c(n_14144), .d(n_14960), .o(n_16222) );
in01f02 FE_RC_218_0 ( .a(n_11733), .o(FE_RN_135_0) );
in01f02 FE_RC_219_0 ( .a(n_10908), .o(FE_RN_136_0) );
no02f02 FE_RC_220_0 ( .a(FE_RN_135_0), .b(FE_RN_136_0), .o(FE_RN_137_0) );
in01f02 FE_RC_222_0 ( .a(n_10699), .o(FE_RN_138_0) );
in01f02 FE_RC_223_0 ( .a(n_10702), .o(FE_RN_139_0) );
no02f02 FE_RC_224_0 ( .a(FE_RN_138_0), .b(FE_RN_139_0), .o(FE_RN_140_0) );
na03f02 TIMEBOOST_cell_65701 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q), .b(g65915_sb), .c(g65915_db), .o(n_3178) );
in01f02 FE_RC_227_0 ( .a(n_11719), .o(FE_RN_141_0) );
in01f02 FE_RC_228_0 ( .a(n_10866), .o(FE_RN_142_0) );
no02f02 FE_RC_229_0 ( .a(FE_RN_141_0), .b(FE_RN_142_0), .o(FE_RN_143_0) );
in01m02 TIMEBOOST_cell_45964 ( .a(TIMEBOOST_net_13924), .o(TIMEBOOST_net_13925) );
in01f02 FE_RC_231_0 ( .a(n_10608), .o(FE_RN_144_0) );
in01f02 FE_RC_232_0 ( .a(n_11735), .o(FE_RN_145_0) );
no02f02 FE_RC_233_0 ( .a(FE_RN_144_0), .b(FE_RN_145_0), .o(FE_RN_146_0) );
na02m02 TIMEBOOST_cell_68278 ( .a(TIMEBOOST_net_21143), .b(g65707_sb), .o(TIMEBOOST_net_21347) );
in01f06 FE_RC_238_0 ( .a(FE_OCPN1850_n_15998), .o(FE_RN_147_0) );
in01f10 FE_RC_239_0 ( .a(FE_OCPN1852_n_16538), .o(FE_RN_148_0) );
na02f20 FE_RC_240_0 ( .a(FE_RN_148_0), .b(FE_RN_147_0), .o(FE_RN_149_0) );
in01f08 FE_RC_242_0 ( .a(n_1399), .o(FE_RN_150_0) );
in01f06 FE_RC_243_0 ( .a(n_2227), .o(FE_RN_151_0) );
na03f02 TIMEBOOST_cell_64882 ( .a(TIMEBOOST_net_16585), .b(FE_OFN785_n_2678), .c(g65250_sb), .o(n_2632) );
in01f04 FE_RC_246_0 ( .a(n_2250), .o(FE_RN_153_0) );
in01f03 FE_RC_247_0 ( .a(n_3466), .o(FE_RN_154_0) );
na02m02 TIMEBOOST_cell_68319 ( .a(TIMEBOOST_net_21367), .b(g64896_db), .o(n_3697) );
na03f02 TIMEBOOST_cell_33524 ( .a(TIMEBOOST_net_8791), .b(FE_OFN1168_n_5592), .c(g62100_sb), .o(n_5603) );
na02f04 TIMEBOOST_cell_40503 ( .a(TIMEBOOST_net_11863), .b(n_7821), .o(FE_RN_176_0) );
in01f02 FE_RC_251_0 ( .a(n_16160), .o(FE_RN_156_0) );
no02f04 FE_RC_253_0 ( .a(FE_RN_156_0), .b(FE_RN_9_0), .o(FE_RN_158_0) );
in01f04 FE_RC_255_0 ( .a(n_4874), .o(FE_RN_159_0) );
in01f02 FE_RC_256_0 ( .a(n_3432), .o(FE_RN_160_0) );
na03f02 TIMEBOOST_cell_73809 ( .a(TIMEBOOST_net_16547), .b(FE_OFN1775_n_13800), .c(FE_OFN1768_n_14054), .o(g53262_p) );
na02f02 TIMEBOOST_cell_72088 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q), .b(g64341_sb), .o(TIMEBOOST_net_23252) );
na03f06 FE_RC_25_0 ( .a(n_16967), .b(n_16974), .c(n_16970), .o(n_13674) );
in01s01 TIMEBOOST_cell_63558 ( .a(TIMEBOOST_net_20738), .o(wbs_adr_i_7_) );
na02m10 TIMEBOOST_cell_28011 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q), .o(TIMEBOOST_net_8110) );
in01f02 FE_RC_282_0 ( .a(FE_RN_176_0), .o(n_13577) );
na03f02 FE_RC_285_0 ( .a(n_14565), .b(n_14473), .c(n_14292), .o(n_14610) );
na03f02 FE_RC_286_0 ( .a(n_14273), .b(n_14460), .c(n_14559), .o(n_14604) );
in01f02 FE_RC_287_0 ( .a(n_10951), .o(FE_RN_177_0) );
in01f02 FE_RC_288_0 ( .a(n_10691), .o(FE_RN_178_0) );
no02f04 FE_RC_289_0 ( .a(FE_RN_178_0), .b(FE_RN_177_0), .o(FE_RN_179_0) );
in01f02 FE_RC_291_0 ( .a(n_10875), .o(FE_RN_180_0) );
in01f02 FE_RC_292_0 ( .a(n_10873), .o(FE_RN_181_0) );
no02f02 FE_RC_293_0 ( .a(FE_RN_180_0), .b(FE_RN_181_0), .o(FE_RN_182_0) );
in01f02 FE_RC_295_0 ( .a(n_10579), .o(FE_RN_183_0) );
in01f02 FE_RC_296_0 ( .a(n_11726), .o(FE_RN_184_0) );
no02f02 FE_RC_297_0 ( .a(FE_RN_183_0), .b(FE_RN_184_0), .o(FE_RN_185_0) );
na03f02 TIMEBOOST_cell_68028 ( .a(TIMEBOOST_net_17540), .b(FE_OFN1268_n_4095), .c(g62505_sb), .o(n_6569) );
in01f02 FE_RC_299_0 ( .a(n_10891), .o(FE_RN_186_0) );
in01f02 FE_RC_300_0 ( .a(n_10576), .o(FE_RN_187_0) );
no02f02 FE_RC_301_0 ( .a(FE_RN_186_0), .b(FE_RN_187_0), .o(FE_RN_188_0) );
in01f02 FE_RC_303_0 ( .a(n_10109), .o(FE_RN_189_0) );
in01f02 FE_RC_304_0 ( .a(n_10685), .o(FE_RN_190_0) );
no02f02 FE_RC_305_0 ( .a(FE_RN_189_0), .b(FE_RN_190_0), .o(FE_RN_191_0) );
na03m02 TIMEBOOST_cell_65885 ( .a(n_3904), .b(g63056_sb), .c(g63056_db), .o(n_5138) );
in01f02 FE_RC_307_0 ( .a(n_10147), .o(FE_RN_192_0) );
in01f02 FE_RC_308_0 ( .a(n_10970), .o(FE_RN_193_0) );
no02f02 FE_RC_309_0 ( .a(FE_RN_192_0), .b(FE_RN_193_0), .o(FE_RN_194_0) );
na03f06 TIMEBOOST_cell_72427 ( .a(n_1515), .b(wishbone_slave_unit_pcim_sm_rdy_in), .c(n_2245), .o(n_6965) );
in01f02 FE_RC_311_0 ( .a(n_10041), .o(FE_RN_195_0) );
in01f02 FE_RC_312_0 ( .a(n_10038), .o(FE_RN_196_0) );
no02f02 FE_RC_313_0 ( .a(FE_RN_195_0), .b(FE_RN_196_0), .o(FE_RN_197_0) );
na02m02 TIMEBOOST_cell_63992 ( .a(n_424), .b(n_4912), .o(TIMEBOOST_net_20982) );
in01s01 FE_RC_315_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q), .o(FE_RN_198_0) );
in01f01 FE_RC_316_0 ( .a(FE_OFN1453_n_10588), .o(FE_RN_199_0) );
no02f02 FE_RC_317_0 ( .a(FE_RN_198_0), .b(FE_RN_199_0), .o(FE_RN_200_0) );
no02f02 FE_RC_318_0 ( .a(n_15590), .b(FE_RN_200_0), .o(n_15591) );
in01f02 FE_RC_319_0 ( .a(n_12914), .o(FE_RN_201_0) );
in01f02 FE_RC_320_0 ( .a(n_12915), .o(FE_RN_202_0) );
no02f02 FE_RC_321_0 ( .a(FE_RN_201_0), .b(FE_RN_202_0), .o(FE_RN_203_0) );
na04f04 FE_RC_324_0 ( .a(n_11992), .b(n_12393), .c(n_12122), .d(n_12276), .o(n_12920) );
na02m04 TIMEBOOST_cell_53359 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q), .b(TIMEBOOST_net_12409), .o(TIMEBOOST_net_16897) );
na03f02 TIMEBOOST_cell_65689 ( .a(TIMEBOOST_net_20389), .b(FE_OFN2128_n_16497), .c(g54310_sb), .o(n_13020) );
na02s02 TIMEBOOST_cell_48920 ( .a(TIMEBOOST_net_14677), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_10880) );
na04f04 FE_RC_328_0 ( .a(n_10524), .b(n_10521), .c(n_9950), .d(n_9953), .o(n_12128) );
ao22f02 FE_RC_329_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q), .b(FE_OFN1731_n_9975), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q), .d(FE_OCP_RBN2005_FE_RN_459_0), .o(n_9332) );
na03f80 FE_RC_32_0 ( .a(n_16910), .b(n_326), .c(n_15204), .o(n_15317) );
na02s01 TIMEBOOST_cell_50017 ( .a(FE_OFN529_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q), .o(TIMEBOOST_net_15226) );
in01f40 FE_RC_335_0 ( .a(pci_target_unit_wishbone_master_read_bound), .o(FE_RN_207_0) );
in01f20 FE_RC_336_0 ( .a(n_16275), .o(FE_RN_208_0) );
no02f20 FE_RC_337_0 ( .a(FE_RN_207_0), .b(FE_RN_208_0), .o(FE_RN_209_0) );
na02m02 TIMEBOOST_cell_52295 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q), .b(g64272_sb), .o(TIMEBOOST_net_16365) );
na02f02 TIMEBOOST_cell_40851 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_12037), .o(n_12626) );
in01f02 FE_RC_341_0 ( .a(n_13667), .o(FE_RN_211_0) );
na03m04 TIMEBOOST_cell_72754 ( .a(TIMEBOOST_net_21577), .b(g65084_sb), .c(TIMEBOOST_net_21831), .o(TIMEBOOST_net_17416) );
na03f02 TIMEBOOST_cell_34960 ( .a(TIMEBOOST_net_9463), .b(FE_OFN1370_n_8567), .c(g57072_sb), .o(n_10497) );
na02f40 TIMEBOOST_cell_45004 ( .a(TIMEBOOST_net_13396), .b(n_15442), .o(n_16438) );
in01f02 FE_RC_345_0 ( .a(n_13571), .o(FE_RN_214_0) );
in01f02 FE_RC_346_0 ( .a(FE_RN_215_0), .o(n_13768) );
na02f04 FE_RC_347_0 ( .a(FE_RN_214_0), .b(FE_RN_213_0), .o(FE_RN_215_0) );
na02f40 FE_RC_348_0 ( .a(n_16492), .b(n_16494), .o(FE_RN_216_0) );
in01f10 FE_RC_349_0 ( .a(n_16490), .o(FE_RN_217_0) );
in01f08 FE_RC_34_0 ( .a(n_15645), .o(FE_RN_15_0) );
in01f10 FE_RC_350_0 ( .a(FE_RN_218_0), .o(n_16495) );
no02f20 FE_RC_351_0 ( .a(FE_RN_216_0), .b(FE_RN_217_0), .o(FE_RN_218_0) );
in01f02 FE_RC_353_0 ( .a(n_10075), .o(FE_RN_219_0) );
in01f02 FE_RC_354_0 ( .a(n_10659), .o(FE_RN_220_0) );
no02f02 FE_RC_355_0 ( .a(FE_RN_219_0), .b(FE_RN_220_0), .o(FE_RN_221_0) );
na04f02 TIMEBOOST_cell_73185 ( .a(g62028_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q), .c(FE_OFN699_n_7845), .d(TIMEBOOST_net_22352), .o(n_7840) );
in01f20 FE_RC_358_0 ( .a(pci_target_unit_pcit_if_strd_bc_in_717), .o(FE_RN_222_0) );
in01f20 FE_RC_359_0 ( .a(pci_target_unit_pcit_if_strd_bc_in_718), .o(FE_RN_223_0) );
no02f20 FE_RC_360_0 ( .a(FE_RN_222_0), .b(FE_RN_223_0), .o(FE_RN_224_0) );
na02f20 FE_RC_361_0 ( .a(FE_RN_224_0), .b(n_1219), .o(n_1507) );
na02m03 TIMEBOOST_cell_68083 ( .a(TIMEBOOST_net_21249), .b(g67069_db), .o(n_1647) );
in01f02 FE_RC_364_0 ( .a(n_10901), .o(FE_RN_225_0) );
in01f02 FE_RC_365_0 ( .a(n_10902), .o(FE_RN_226_0) );
no02f02 FE_RC_366_0 ( .a(FE_RN_225_0), .b(FE_RN_226_0), .o(FE_RN_227_0) );
na02m04 TIMEBOOST_cell_69389 ( .a(TIMEBOOST_net_21902), .b(g64860_sb), .o(TIMEBOOST_net_12691) );
in01f02 FE_RC_368_0 ( .a(n_10569), .o(FE_RN_228_0) );
in01f02 FE_RC_369_0 ( .a(n_11723), .o(FE_RN_229_0) );
no02f02 FE_RC_370_0 ( .a(FE_RN_228_0), .b(FE_RN_229_0), .o(FE_RN_230_0) );
in01s01 TIMEBOOST_cell_73833 ( .a(TIMEBOOST_net_23397), .o(TIMEBOOST_net_23398) );
na03m04 TIMEBOOST_cell_72494 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q), .b(n_3741), .c(TIMEBOOST_net_21682), .o(TIMEBOOST_net_17071) );
na04f04 TIMEBOOST_cell_73115 ( .a(n_1563), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q), .c(FE_OFN716_n_8176), .d(g61937_sb), .o(n_7949) );
na02s01 TIMEBOOST_cell_47754 ( .a(TIMEBOOST_net_14094), .b(FE_OFN606_n_9904), .o(TIMEBOOST_net_10316) );
in01f02 FE_RC_375_0 ( .a(n_9979), .o(FE_RN_231_0) );
in01f02 FE_RC_376_0 ( .a(n_10877), .o(FE_RN_232_0) );
no02f02 FE_RC_377_0 ( .a(FE_RN_232_0), .b(FE_RN_231_0), .o(FE_RN_233_0) );
na03m04 TIMEBOOST_cell_70326 ( .a(g65845_db), .b(TIMEBOOST_net_16328), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_22371) );
na03f02 FE_RC_379_0 ( .a(n_16227), .b(n_16228), .c(n_16230), .o(n_16231) );
na03f02 FE_RC_380_0 ( .a(n_16625), .b(n_14446), .c(n_16624), .o(n_14597) );
na03f02 FE_RC_381_0 ( .a(n_16239), .b(n_16237), .c(n_16234), .o(n_16240) );
na03f02 FE_RC_382_0 ( .a(n_14402), .b(n_14494), .c(n_14534), .o(n_14578) );
na03f02 FE_RC_383_0 ( .a(n_14547), .b(n_14435), .c(n_14250), .o(n_14592) );
na03f02 FE_RC_384_0 ( .a(n_14541), .b(n_14421), .c(n_14420), .o(n_14585) );
na03f02 FE_RC_385_0 ( .a(n_14563), .b(n_14286), .c(n_14468), .o(n_14608) );
na03f02 FE_RC_386_0 ( .a(n_14545), .b(n_14431), .c(n_14513), .o(n_14590) );
na03f02 FE_RC_387_0 ( .a(n_16251), .b(n_16253), .c(n_16248), .o(n_16254) );
na03f02 FE_RC_389_0 ( .a(n_14261), .b(n_16623), .c(n_16622), .o(n_14598) );
na04f02 FE_RC_390_0 ( .a(n_12962), .b(n_12939), .c(n_12940), .d(n_12805), .o(n_13143) );
na03f02 FE_RC_391_0 ( .a(n_12960), .b(n_13034), .c(n_12677), .o(n_13319) );
in01f02 FE_RC_392_0 ( .a(n_12721), .o(FE_RN_234_0) );
in01f02 FE_RC_393_0 ( .a(n_12929), .o(FE_RN_235_0) );
no02f02 FE_RC_394_0 ( .a(FE_RN_235_0), .b(FE_RN_234_0), .o(FE_RN_236_0) );
na04f02 FE_RC_396_0 ( .a(n_13054), .b(n_12903), .c(n_12791), .d(n_12902), .o(n_13137) );
na04f03 FE_RC_397_0 ( .a(n_13055), .b(n_12906), .c(n_12907), .d(n_12792), .o(n_13138) );
in01s01 FE_RC_401_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q), .o(FE_RN_237_0) );
in01f02 FE_RC_402_0 ( .a(FE_OFN1565_n_12502), .o(FE_RN_238_0) );
na02f02 TIMEBOOST_cell_26566 ( .a(TIMEBOOST_net_7387), .b(FE_OCPN1909_n_16497), .o(TIMEBOOST_net_387) );
na03f02 TIMEBOOST_cell_72419 ( .a(n_4939), .b(FE_OFN276_n_9941), .c(TIMEBOOST_net_21317), .o(TIMEBOOST_net_20666) );
in01s01 FE_RC_405_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q), .o(FE_RN_240_0) );
in01f02 FE_RC_406_0 ( .a(FE_OFN1563_n_12502), .o(FE_RN_241_0) );
na04m02 TIMEBOOST_cell_67851 ( .a(n_3749), .b(FE_OFN1640_n_4671), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q), .d(g65415_sb), .o(TIMEBOOST_net_7597) );
na03f02 TIMEBOOST_cell_66816 ( .a(TIMEBOOST_net_16840), .b(FE_OFN1345_n_8567), .c(g57489_sb), .o(n_11247) );
in01s01 FE_RC_409_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q), .o(FE_RN_243_0) );
in01f04 FE_RC_410_0 ( .a(FE_OFN1563_n_12502), .o(FE_RN_244_0) );
na03f02 TIMEBOOST_cell_72938 ( .a(pci_target_unit_del_sync_addr_in_229), .b(g65218_sb), .c(TIMEBOOST_net_7152), .o(n_2669) );
na03s02 TIMEBOOST_cell_73654 ( .a(FE_OFN532_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q), .c(TIMEBOOST_net_22921), .o(TIMEBOOST_net_14937) );
in01s01 FE_RC_413_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q), .o(FE_RN_246_0) );
in01f01 FE_RC_414_0 ( .a(FE_OFN1563_n_12502), .o(FE_RN_247_0) );
na02m02 TIMEBOOST_cell_68466 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q), .b(n_3764), .o(TIMEBOOST_net_21441) );
in01f10 TIMEBOOST_cell_17841 ( .a(TIMEBOOST_net_5252), .o(n_13721) );
na04f04 FE_RC_418_0 ( .a(n_11961), .b(n_12117), .c(n_11962), .d(n_12379), .o(n_12904) );
in01f02 FE_RC_41_0 ( .a(n_12881), .o(FE_RN_18_0) );
in01f02 FE_RC_422_0 ( .a(n_11991), .o(FE_RN_249_0) );
in01f02 FE_RC_423_0 ( .a(n_11990), .o(FE_RN_250_0) );
no02f02 FE_RC_424_0 ( .a(FE_RN_250_0), .b(FE_RN_249_0), .o(FE_RN_251_0) );
na02f02 FE_RC_425_0 ( .a(FE_RN_29_0), .b(FE_RN_251_0), .o(n_12816) );
in01f02 FE_RC_42_0 ( .a(n_12880), .o(FE_RN_19_0) );
in01f03 FE_RC_437_0 ( .a(FE_RN_259_0), .o(n_13410) );
na02f03 FE_RC_438_0 ( .a(n_13122), .b(n_16299), .o(FE_RN_259_0) );
in01f10 FE_RC_439_0 ( .a(pci_target_unit_pci_target_sm_wr_to_fifo), .o(FE_RN_260_0) );
no02f02 FE_RC_43_0 ( .a(FE_RN_18_0), .b(FE_RN_19_0), .o(FE_RN_20_0) );
in01f01 FE_RC_440_0 ( .a(n_978), .o(FE_RN_261_0) );
no02f02 FE_RC_441_0 ( .a(FE_RN_260_0), .b(FE_RN_261_0), .o(FE_RN_262_0) );
in01f01 FE_RC_442_0 ( .a(n_653), .o(FE_RN_263_0) );
no02f02 FE_RC_443_0 ( .a(FE_RN_263_0), .b(pci_target_unit_pci_target_sm_state_transfere_reg), .o(FE_RN_264_0) );
na03m02 TIMEBOOST_cell_72739 ( .a(TIMEBOOST_net_21572), .b(g64344_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q), .o(TIMEBOOST_net_22412) );
in01s01 TIMEBOOST_cell_63589 ( .a(TIMEBOOST_net_20769), .o(TIMEBOOST_net_20768) );
na03f02 TIMEBOOST_cell_34884 ( .a(TIMEBOOST_net_9325), .b(FE_OFN1381_n_8567), .c(g57311_sb), .o(n_10402) );
no02f02 FE_RC_448_0 ( .a(n_1724), .b(pci_target_unit_pci_target_sm_cnf_progress), .o(FE_RN_269_0) );
in01f02 FE_RC_449_0 ( .a(n_2031), .o(FE_RN_270_0) );
na03f02 FE_RC_44_0 ( .a(FE_RN_20_0), .b(n_12957), .c(n_12632), .o(n_13131) );
in01f10 FE_RC_450_0 ( .a(pci_target_unit_pci_target_sm_state_backoff_reg_reg_Q), .o(FE_RN_271_0) );
na02s02 TIMEBOOST_cell_31398 ( .a(TIMEBOOST_net_9803), .b(FE_OFN704_n_8069), .o(n_8100) );
oa12f06 FE_RC_453_0 ( .a(FE_RN_267_0), .b(FE_RN_268_0), .c(FE_RN_273_0), .o(n_8566) );
in01f40 FE_RC_454_0 ( .a(n_2078), .o(FE_RN_274_0) );
na02f40 FE_RC_455_0 ( .a(FE_RN_274_0), .b(n_525), .o(n_16287) );
in01s01 FE_RC_456_0 ( .a(parchk_pci_cbe_out_in_1204), .o(FE_RN_275_0) );
in01f03 FE_RC_457_0 ( .a(n_4702), .o(FE_RN_276_0) );
ao22f04 FE_RC_458_0 ( .a(FE_RN_275_0), .b(FE_RN_276_0), .c(parchk_pci_cbe_out_in_1204), .d(n_4702), .o(n_4703) );
in01m01 FE_RC_460_0 ( .a(n_532), .o(FE_RN_278_0) );
na02f04 FE_RC_461_0 ( .a(n_1196), .b(FE_RN_278_0), .o(FE_RN_279_0) );
na02f06 FE_RC_462_0 ( .a(FE_RN_279_0), .b(n_15292), .o(FE_RN_280_0) );
in01f04 FE_RC_463_0 ( .a(n_15607), .o(FE_RN_281_0) );
na02f02 TIMEBOOST_cell_70637 ( .a(TIMEBOOST_net_22526), .b(g62731_sb), .o(n_5517) );
in01s01 TIMEBOOST_cell_45903 ( .a(TIMEBOOST_net_13915), .o(TIMEBOOST_net_13864) );
in01s01 FE_RC_467_0 ( .a(parchk_pci_cbe_out_in), .o(FE_RN_284_0) );
in01f02 FE_RC_468_0 ( .a(n_4703), .o(FE_RN_285_0) );
na02m02 TIMEBOOST_cell_44481 ( .a(n_3361), .b(n_2092), .o(TIMEBOOST_net_13135) );
na04f20 FE_RC_481_0 ( .a(n_653), .b(pci_target_unit_pci_target_sm_same_read_reg), .c(n_1724), .d(pci_target_unit_pci_target_sm_rd_from_fifo), .o(FE_RN_294_0) );
no02f10 FE_RC_482_0 ( .a(FE_RN_294_0), .b(n_1435), .o(n_15401) );
no02f80 FE_RC_483_0 ( .a(wbm_ack_i), .b(FE_RN_295_0), .o(n_1445) );
na02f80 FE_RC_484_0 ( .a(n_705), .b(wbm_err_i), .o(FE_RN_295_0) );
na04f02 FE_RC_490_0 ( .a(n_11092), .b(n_11093), .c(n_11094), .d(n_11091), .o(n_12544) );
na04f02 FE_RC_491_0 ( .a(n_11130), .b(n_11792), .c(n_10791), .d(n_11791), .o(n_12771) );
na03f80 TIMEBOOST_cell_7 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_), .b(FE_RN_552_0), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_), .o(n_16462) );
in01f20 FE_RC_493_0 ( .a(FE_RN_299_0), .o(n_15981) );
na02f02 TIMEBOOST_cell_30587 ( .a(n_9440), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q), .o(TIMEBOOST_net_9398) );
na02f06 FE_RC_497_0 ( .a(n_16511), .b(n_16268), .o(n_14967) );
na02s02 TIMEBOOST_cell_43812 ( .a(TIMEBOOST_net_12800), .b(g58232_sb), .o(TIMEBOOST_net_10825) );
na04f02 TIMEBOOST_cell_73347 ( .a(TIMEBOOST_net_11133), .b(g65680_sb), .c(g63435_sb), .d(TIMEBOOST_net_5504), .o(n_4625) );
na02f02 FE_RC_49_0 ( .a(FE_RN_23_0), .b(n_13061), .o(n_13321) );
in01f10 FE_RC_501_0 ( .a(pciu_bar0_in_378), .o(FE_RN_303_0) );
in01f20 FE_RC_502_0 ( .a(n_396), .o(FE_RN_304_0) );
ao22f10 FE_RC_503_0 ( .a(FE_RN_303_0), .b(FE_RN_304_0), .c(pciu_bar0_in_378), .d(n_396), .o(FE_RN_305_0) );
na04m02 TIMEBOOST_cell_67850 ( .a(n_3752), .b(FE_OFN640_n_4669), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q), .d(g65393_sb), .o(n_3523) );
no02f20 FE_RC_505_0 ( .a(pciu_bar0_in_379), .b(parchk_pci_ad_reg_in_1235), .o(FE_RN_307_0) );
ao12f06 FE_RC_506_0 ( .a(FE_RN_307_0), .b(pciu_bar0_in_379), .c(parchk_pci_ad_reg_in_1235), .o(FE_RN_308_0) );
no02f20 FE_RC_507_0 ( .a(pciu_bar0_in_376), .b(parchk_pci_ad_reg_in_1232), .o(FE_RN_309_0) );
ao12f08 FE_RC_508_0 ( .a(FE_RN_309_0), .b(pciu_bar0_in_376), .c(parchk_pci_ad_reg_in_1232), .o(FE_RN_310_0) );
no02f20 FE_RC_509_0 ( .a(pciu_bar0_in_377), .b(parchk_pci_ad_reg_in_1233), .o(FE_RN_311_0) );
ao12f10 FE_RC_510_0 ( .a(FE_RN_311_0), .b(pciu_bar0_in_377), .c(parchk_pci_ad_reg_in_1233), .o(FE_RN_312_0) );
no02f06 FE_RC_511_0 ( .a(FE_RN_310_0), .b(FE_RN_312_0), .o(FE_RN_313_0) );
no02f20 FE_RC_512_0 ( .a(pciu_bar0_in), .b(parchk_pci_ad_reg_in_1216), .o(FE_RN_314_0) );
ao12f08 FE_RC_513_0 ( .a(FE_RN_314_0), .b(pciu_bar0_in), .c(parchk_pci_ad_reg_in_1216), .o(FE_RN_315_0) );
no02f40 FE_RC_514_0 ( .a(pciu_bar0_in_362), .b(parchk_pci_ad_reg_in_1218), .o(FE_RN_316_0) );
ao12f10 FE_RC_515_0 ( .a(FE_RN_316_0), .b(pciu_bar0_in_362), .c(parchk_pci_ad_reg_in_1218), .o(FE_RN_317_0) );
na02f40 FE_RC_516_0 ( .a(pciu_bar0_in_363), .b(parchk_pci_ad_reg_in_1219), .o(FE_RN_318_0) );
oa12f10 FE_RC_517_0 ( .a(FE_RN_318_0), .b(pciu_bar0_in_363), .c(parchk_pci_ad_reg_in_1219), .o(FE_RN_319_0) );
na02f40 FE_RC_518_0 ( .a(pciu_bar0_in_361), .b(parchk_pci_ad_reg_in_1217), .o(FE_RN_320_0) );
oa12f10 FE_RC_519_0 ( .a(FE_RN_320_0), .b(pciu_bar0_in_361), .c(parchk_pci_ad_reg_in_1217), .o(FE_RN_321_0) );
in01f02 FE_RC_51_0 ( .a(n_12032), .o(FE_RN_25_0) );
na02f10 FE_RC_520_0 ( .a(FE_RN_319_0), .b(FE_RN_321_0), .o(FE_RN_322_0) );
na02f40 FE_RC_522_0 ( .a(pciu_bar0_in_367), .b(parchk_pci_ad_reg_in_1223), .o(FE_RN_324_0) );
oa12f10 FE_RC_523_0 ( .a(FE_RN_324_0), .b(pciu_bar0_in_367), .c(parchk_pci_ad_reg_in_1223), .o(FE_RN_325_0) );
na02f40 FE_RC_524_0 ( .a(pciu_bar0_in_364), .b(parchk_pci_ad_reg_in_1220), .o(FE_RN_326_0) );
oa12f10 FE_RC_525_0 ( .a(FE_RN_326_0), .b(pciu_bar0_in_364), .c(parchk_pci_ad_reg_in_1220), .o(FE_RN_327_0) );
na02f08 FE_RC_526_0 ( .a(FE_RN_325_0), .b(FE_RN_327_0), .o(FE_RN_328_0) );
no02f10 FE_RC_527_0 ( .a(pciu_bar0_in_365), .b(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(FE_RN_329_0) );
ao12f06 FE_RC_528_0 ( .a(FE_RN_329_0), .b(pciu_bar0_in_365), .c(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(FE_RN_330_0) );
no02f10 FE_RC_529_0 ( .a(pciu_bar0_in_366), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(FE_RN_331_0) );
ao12f06 FE_RC_530_0 ( .a(FE_RN_331_0), .b(pciu_bar0_in_366), .c(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(FE_RN_332_0) );
na02f20 FE_RC_532_0 ( .a(pciu_bar0_in_368), .b(parchk_pci_ad_reg_in_1224), .o(FE_RN_334_0) );
oa12f10 FE_RC_533_0 ( .a(FE_RN_334_0), .b(pciu_bar0_in_368), .c(parchk_pci_ad_reg_in_1224), .o(FE_RN_335_0) );
na02f20 FE_RC_534_0 ( .a(parchk_pci_ad_reg_in_1225), .b(pciu_bar0_in_369), .o(FE_RN_336_0) );
oa12f10 FE_RC_535_0 ( .a(FE_RN_336_0), .b(pciu_bar0_in_369), .c(parchk_pci_ad_reg_in_1225), .o(FE_RN_337_0) );
na02f08 FE_RC_536_0 ( .a(FE_RN_335_0), .b(FE_RN_337_0), .o(FE_RN_338_0) );
na02f20 FE_RC_537_0 ( .a(pciu_bar0_in_373), .b(parchk_pci_ad_reg_in_1229), .o(FE_RN_339_0) );
oa12f10 FE_RC_538_0 ( .a(FE_RN_339_0), .b(pciu_bar0_in_373), .c(parchk_pci_ad_reg_in_1229), .o(FE_RN_340_0) );
na02f40 FE_RC_539_0 ( .a(pciu_bar0_in_374), .b(parchk_pci_ad_reg_in_1230), .o(FE_RN_341_0) );
na03m02 TIMEBOOST_cell_73203 ( .a(TIMEBOOST_net_22080), .b(FE_OFN2256_n_8060), .c(g61901_sb), .o(n_8021) );
oa12f10 FE_RC_540_0 ( .a(FE_RN_341_0), .b(pciu_bar0_in_374), .c(parchk_pci_ad_reg_in_1230), .o(FE_RN_342_0) );
na02f08 FE_RC_541_0 ( .a(FE_RN_340_0), .b(FE_RN_342_0), .o(FE_RN_343_0) );
na02f40 FE_RC_542_0 ( .a(pciu_bar0_in_370), .b(parchk_pci_ad_reg_in_1226), .o(FE_RN_344_0) );
oa12f10 FE_RC_543_0 ( .a(FE_RN_344_0), .b(pciu_bar0_in_370), .c(parchk_pci_ad_reg_in_1226), .o(FE_RN_345_0) );
na02f20 FE_RC_544_0 ( .a(pciu_bar0_in_371), .b(parchk_pci_ad_reg_in_1227), .o(FE_RN_346_0) );
oa12f10 FE_RC_545_0 ( .a(FE_RN_346_0), .b(pciu_bar0_in_371), .c(parchk_pci_ad_reg_in_1227), .o(FE_RN_347_0) );
na02f08 FE_RC_546_0 ( .a(FE_RN_345_0), .b(FE_RN_347_0), .o(FE_RN_348_0) );
na02f20 FE_RC_547_0 ( .a(pciu_bar0_in_372), .b(parchk_pci_ad_reg_in_1228), .o(FE_RN_349_0) );
oa12f10 FE_RC_548_0 ( .a(FE_RN_349_0), .b(pciu_bar0_in_372), .c(parchk_pci_ad_reg_in_1228), .o(FE_RN_350_0) );
na02f20 FE_RC_549_0 ( .a(pciu_bar0_in_375), .b(parchk_pci_ad_reg_in_1231), .o(FE_RN_351_0) );
in01f02 FE_RC_54_0 ( .a(n_12275), .o(FE_RN_27_0) );
oa12f10 FE_RC_550_0 ( .a(FE_RN_351_0), .b(pciu_bar0_in_375), .c(parchk_pci_ad_reg_in_1231), .o(FE_RN_352_0) );
na02f08 FE_RC_551_0 ( .a(FE_RN_350_0), .b(FE_RN_352_0), .o(FE_RN_353_0) );
no02f02 FE_RC_554_0 ( .a(FE_RN_308_0), .b(FE_RN_355_0), .o(FE_RN_356_0) );
na02s01 TIMEBOOST_cell_29231 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q), .b(g64224_sb), .o(TIMEBOOST_net_8720) );
in01f10 FE_RC_557_0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_control_in), .o(FE_RN_357_0) );
na02f10 FE_RC_558_0 ( .a(FE_RN_357_0), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in_85), .o(FE_RN_358_0) );
in01f02 FE_RC_559_0 ( .a(n_16980), .o(FE_RN_359_0) );
in01f02 FE_RC_55_0 ( .a(n_12274), .o(FE_RN_28_0) );
no02f06 FE_RC_560_0 ( .a(FE_RN_359_0), .b(FE_RN_358_0), .o(FE_RN_360_0) );
in01f01 FE_RC_562_0 ( .a(n_13763), .o(FE_RN_361_0) );
in01f02 FE_RC_563_0 ( .a(n_13666), .o(FE_RN_362_0) );
na02m02 TIMEBOOST_cell_68129 ( .a(TIMEBOOST_net_21272), .b(g54171_sb), .o(TIMEBOOST_net_16140) );
in01f02 FE_RC_567_0 ( .a(n_13566), .o(FE_RN_365_0) );
in01f02 FE_RC_568_0 ( .a(FE_RN_366_0), .o(n_13761) );
na03f02 TIMEBOOST_cell_72523 ( .a(TIMEBOOST_net_21387), .b(g64207_sb), .c(FE_OFN2106_g64577_p), .o(TIMEBOOST_net_22468) );
no02f02 FE_RC_56_0 ( .a(FE_RN_28_0), .b(FE_RN_27_0), .o(FE_RN_29_0) );
na02s01 TIMEBOOST_cell_47753 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q), .o(TIMEBOOST_net_14094) );
in01f02 FE_RC_571_0 ( .a(n_13568), .o(FE_RN_368_0) );
in01f02 FE_RC_572_0 ( .a(FE_RN_369_0), .o(n_13764) );
in01f01 FE_RC_574_0 ( .a(n_7822), .o(FE_RN_370_0) );
in01f02 FE_RC_575_0 ( .a(n_13028), .o(FE_RN_371_0) );
na02f02 TIMEBOOST_cell_27784 ( .a(TIMEBOOST_net_7996), .b(n_14387), .o(n_14394) );
na03f02 TIMEBOOST_cell_34955 ( .a(TIMEBOOST_net_9457), .b(FE_OFN1422_n_8567), .c(g57443_sb), .o(n_11290) );
in01f01 FE_RC_578_0 ( .a(n_13354), .o(FE_RN_373_0) );
in01f02 FE_RC_579_0 ( .a(n_12982), .o(FE_RN_374_0) );
na04f02 TIMEBOOST_cell_73586 ( .a(TIMEBOOST_net_15048), .b(TIMEBOOST_net_7275), .c(TIMEBOOST_net_21012), .d(n_13921), .o(n_14628) );
na02f02 TIMEBOOST_cell_42931 ( .a(g65904_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q), .o(TIMEBOOST_net_12360) );
in01f02 FE_RC_582_0 ( .a(n_13354), .o(FE_RN_376_0) );
in01f02 FE_RC_583_0 ( .a(n_12984), .o(FE_RN_377_0) );
na02m01 TIMEBOOST_cell_62778 ( .a(n_4476), .b(n_0), .o(TIMEBOOST_net_20336) );
na03m02 TIMEBOOST_cell_72687 ( .a(g64970_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q), .c(TIMEBOOST_net_16269), .o(TIMEBOOST_net_17561) );
na03f02 TIMEBOOST_cell_67026 ( .a(FE_OFN1606_n_13997), .b(TIMEBOOST_net_13746), .c(FE_OFN1599_n_13995), .o(n_14457) );
in01f10 FE_RC_589_0 ( .a(FE_RN_381_0), .o(n_16791) );
na02f10 FE_RC_590_0 ( .a(n_15755), .b(n_16002), .o(FE_RN_381_0) );
in01f04 FE_RC_591_0 ( .a(n_16578), .o(FE_RN_382_0) );
no02f08 FE_RC_592_0 ( .a(FE_RN_382_0), .b(n_16573), .o(n_15453) );
na02f02 FE_RC_593_0 ( .a(parchk_pci_ad_out_in_1191), .b(FE_OFN1709_n_4868), .o(FE_RN_383_0) );
na02f02 FE_RC_594_0 ( .a(FE_RN_383_0), .b(n_14345), .o(n_14376) );
na03f06 FE_RC_597_0 ( .a(FE_OCP_RBN2016_n_16970), .b(n_14939), .c(n_16205), .o(n_13701) );
na02f01 TIMEBOOST_cell_18156 ( .a(TIMEBOOST_net_5441), .b(g65813_sb), .o(n_2570) );
in01f20 FE_RC_599_0 ( .a(FE_RN_384_0), .o(n_15919) );
na02f20 FE_RC_600_0 ( .a(n_16015), .b(n_16016), .o(FE_RN_384_0) );
in01f04 FE_RC_601_0 ( .a(FE_RN_385_0), .o(n_8800) );
no02f04 FE_RC_602_0 ( .a(n_16331), .b(n_9175), .o(FE_RN_385_0) );
no02f20 FE_RC_604_0 ( .a(n_16275), .b(configuration_sync_cache_lsize_to_wb_bits_reg_3__Q), .o(FE_RN_387_0) );
na02f10 FE_RC_605_0 ( .a(FE_RN_387_0), .b(FE_RN_386_0), .o(n_16280) );
in01f20 FE_RC_606_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(FE_RN_388_0) );
na02f10 FE_RC_607_0 ( .a(n_16576), .b(FE_RN_388_0), .o(FE_RN_389_0) );
oa12f10 FE_RC_608_0 ( .a(FE_RN_389_0), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .c(n_16576), .o(n_16577) );
in01f02 FE_RC_60_0 ( .a(n_10202), .o(FE_RN_30_0) );
na02f06 FE_RC_610_0 ( .a(n_15014), .b(n_15055), .o(FE_RN_390_0) );
no02f10 FE_RC_612_0 ( .a(n_12179), .b(n_15762), .o(FE_RN_392_0) );
in01f04 FE_RC_613_0 ( .a(n_15760), .o(FE_RN_393_0) );
in01f04 FE_RC_614_0 ( .a(n_15759), .o(FE_RN_394_0) );
no02f08 FE_RC_615_0 ( .a(FE_RN_393_0), .b(FE_RN_394_0), .o(FE_RN_395_0) );
ao12f08 FE_RC_616_0 ( .a(FE_RN_392_0), .b(FE_RN_395_0), .c(n_15758), .o(FE_OFN1503_n_15768) );
in01m20 FE_RC_617_0 ( .a(n_13784), .o(FE_RN_396_0) );
na02f01 FE_RC_618_0 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q), .b(FE_OFN2126_n_16497), .o(FE_RN_397_0) );
in01s01 FE_RC_619_0 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_773), .o(FE_RN_398_0) );
in01f02 FE_RC_61_0 ( .a(n_10205), .o(FE_RN_31_0) );
oa12f02 FE_RC_620_0 ( .a(FE_RN_397_0), .b(FE_RN_398_0), .c(FE_OFN2126_n_16497), .o(FE_RN_399_0) );
na02f02 FE_RC_621_0 ( .a(n_12595), .b(FE_RN_399_0), .o(FE_RN_400_0) );
in01f01 FE_RC_622_0 ( .a(n_3295), .o(FE_RN_401_0) );
ao22f01 FE_RC_623_0 ( .a(configuration_pci_err_cs_bit8), .b(n_3252), .c(configuration_sync_command_bit8), .d(n_3248), .o(FE_RN_402_0) );
ao22f01 FE_RC_624_0 ( .a(configuration_wb_err_addr_540), .b(n_15444), .c(n_2844), .d(n_16000), .o(FE_RN_403_0) );
na02s01 TIMEBOOST_cell_18211 ( .a(n_6986), .b(g60603_da), .o(TIMEBOOST_net_5469) );
ao22f01 FE_RC_626_0 ( .a(configuration_pci_err_addr_478), .b(FE_OFN1006_n_16288), .c(wbu_latency_tim_val_in), .d(FE_OFN1694_n_3368), .o(FE_RN_405_0) );
in01s01 FE_RC_627_0 ( .a(configuration_wb_err_data_578), .o(FE_RN_406_0) );
in01f01 FE_RC_628_0 ( .a(FE_OFN1068_n_15729), .o(FE_RN_407_0) );
no02f02 FE_RC_62_0 ( .a(FE_RN_30_0), .b(FE_RN_31_0), .o(FE_RN_32_0) );
in01f01 FE_RC_630_0 ( .a(FE_OCPN1845_n_16427), .o(FE_RN_409_0) );
oa22f02 FE_RC_631_0 ( .a(FE_RN_406_0), .b(FE_RN_407_0), .c(FE_RN_678_0), .d(FE_RN_409_0), .o(FE_RN_410_0) );
na02s03 TIMEBOOST_cell_68188 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q), .o(TIMEBOOST_net_21302) );
na02m02 TIMEBOOST_cell_68333 ( .a(TIMEBOOST_net_21374), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_17522) );
na03f02 TIMEBOOST_cell_66896 ( .a(FE_OFN1748_n_12004), .b(TIMEBOOST_net_13558), .c(n_11977), .o(n_12744) );
no02f02 FE_RC_637_0 ( .a(FE_RN_415_0), .b(FE_RN_410_0), .o(FE_RN_416_0) );
na02f02 FE_RC_638_0 ( .a(FE_RN_416_0), .b(FE_RN_405_0), .o(FE_RN_417_0) );
no02f02 FE_RC_639_0 ( .a(FE_RN_417_0), .b(FE_RN_404_0), .o(FE_RN_418_0) );
oa12f02 FE_RC_640_0 ( .a(FE_RN_400_0), .b(n_12595), .c(FE_RN_418_0), .o(FE_RN_419_0) );
ao22f01 FE_RC_641_0 ( .a(conf_wb_err_addr_in_949), .b(n_2115), .c(wishbone_slave_unit_pcim_sm_data_in_642), .d(FE_OFN1610_n_2122), .o(FE_RN_420_0) );
na02f08 FE_RC_642_0 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q), .b(FE_OCPN1913_FE_OFN1150_n_13249), .o(FE_RN_421_0) );
in01s01 FE_RC_643_0 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_391), .o(FE_RN_422_0) );
oa12f04 FE_RC_644_0 ( .a(FE_RN_421_0), .b(FE_RN_422_0), .c(FE_OCPN1913_FE_OFN1150_n_13249), .o(FE_RN_423_0) );
ao22f02 FE_RC_647_0 ( .a(FE_RN_396_0), .b(FE_RN_419_0), .c(n_13784), .d(FE_RN_425_0), .o(FE_RN_426_0) );
in01f02 FE_RC_648_0 ( .a(FE_RN_427_0), .o(n_14323) );
no02f02 FE_RC_649_0 ( .a(FE_RN_426_0), .b(FE_OFN1708_n_4868), .o(FE_RN_427_0) );
in01f02 FE_RC_64_0 ( .a(n_10738), .o(FE_RN_33_0) );
na02f40 FE_RC_650_0 ( .a(n_16462), .b(n_15823), .o(FE_RN_428_0) );
no02f20 FE_RC_651_0 ( .a(FE_OCP_RBN2270_g75061_p), .b(n_16262), .o(FE_RN_429_0) );
na02f20 FE_RC_652_0 ( .a(FE_RN_429_0), .b(n_15824), .o(FE_RN_430_0) );
in01s01 FE_RC_654_0 ( .a(n_7822), .o(FE_RN_431_0) );
ao22f02 FE_RC_655_0 ( .a(configuration_pci_err_data_520), .b(FE_OFN1063_n_15808), .c(n_14922), .d(FE_OCPN1900_n_16810), .o(FE_RN_432_0) );
ao22f02 FE_RC_656_0 ( .a(configuration_wb_err_data_589), .b(FE_OFN1069_n_15729), .c(n_15598), .d(FE_OCPN1845_n_16427), .o(FE_RN_433_0) );
na02f02 FE_RC_657_0 ( .a(FE_RN_432_0), .b(FE_RN_433_0), .o(FE_RN_434_0) );
na03s02 TIMEBOOST_cell_64651 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q), .b(FE_OFN542_n_9690), .c(TIMEBOOST_net_14670), .o(TIMEBOOST_net_12773) );
na02s01 TIMEBOOST_cell_37470 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(g65753_sb), .o(TIMEBOOST_net_10347) );
in01f02 FE_RC_65_0 ( .a(n_10160), .o(FE_RN_34_0) );
ao22f01 FE_RC_660_0 ( .a(configuration_wb_err_addr_551), .b(n_15445), .c(configuration_pci_err_addr_489), .d(FE_OFN1006_n_16288), .o(FE_RN_437_0) );
ao22f04 FE_RC_661_0 ( .a(pciu_am1_in_528), .b(FE_OCPN1903_FE_OFN1061_n_16720), .c(pciu_bar0_in_367), .d(FE_OCPN1898_n_3231), .o(FE_RN_438_0) );
no02f02 FE_RC_663_0 ( .a(FE_RN_439_0), .b(FE_RN_434_0), .o(FE_RN_440_0) );
na02f02 FE_RC_664_0 ( .a(FE_RN_440_0), .b(n_4880), .o(FE_RN_441_0) );
na02f01 FE_RC_665_0 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q), .b(FE_OFN2126_n_16497), .o(FE_RN_442_0) );
in01s01 FE_RC_666_0 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_784), .o(FE_RN_443_0) );
oa12f02 FE_RC_667_0 ( .a(FE_RN_442_0), .b(FE_RN_443_0), .c(FE_OFN2126_n_16497), .o(FE_RN_444_0) );
ao22f02 FE_RC_668_0 ( .a(FE_RN_431_0), .b(FE_RN_441_0), .c(n_7822), .d(FE_RN_444_0), .o(FE_RN_445_0) );
no02f02 FE_RC_669_0 ( .a(FE_RN_445_0), .b(n_13784), .o(FE_RN_446_0) );
no02f02 FE_RC_66_0 ( .a(FE_RN_33_0), .b(FE_RN_34_0), .o(FE_RN_35_0) );
ao22f01 FE_RC_670_0 ( .a(conf_wb_err_addr_in_960), .b(FE_OFN1620_n_1787), .c(wishbone_slave_unit_pcim_sm_data_in_653), .d(FE_OFN1611_n_2122), .o(FE_RN_447_0) );
na02f02 FE_RC_671_0 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q), .b(FE_OCPN1911_FE_OFN1152_n_13249), .o(FE_RN_448_0) );
in01s01 FE_RC_672_0 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_402), .o(FE_RN_449_0) );
oa12f02 FE_RC_673_0 ( .a(FE_RN_448_0), .b(FE_RN_449_0), .c(FE_OCPN1911_FE_OFN1152_n_13249), .o(FE_RN_450_0) );
in01s01 TIMEBOOST_cell_73863 ( .a(TIMEBOOST_net_23427), .o(TIMEBOOST_net_23428) );
na03m02 TIMEBOOST_cell_72866 ( .a(TIMEBOOST_net_21764), .b(g65068_sb), .c(TIMEBOOST_net_21928), .o(TIMEBOOST_net_17366) );
ao12f02 FE_RC_676_0 ( .a(FE_RN_446_0), .b(n_13781), .c(FE_RN_452_0), .o(FE_RN_453_0) );
in01f02 FE_RC_677_0 ( .a(FE_RN_454_0), .o(n_14351) );
no02f02 FE_RC_678_0 ( .a(FE_RN_453_0), .b(FE_OFN1706_n_4868), .o(FE_RN_454_0) );
na02m01 TIMEBOOST_cell_47721 ( .a(TIMEBOOST_net_10178), .b(FE_OFN945_n_2248), .o(TIMEBOOST_net_14078) );
in01f02 FE_RC_680_0 ( .a(n_13565), .o(FE_RN_456_0) );
in01f02 FE_RC_681_0 ( .a(FE_RN_457_0), .o(n_13760) );
na02f02 TIMEBOOST_cell_71005 ( .a(TIMEBOOST_net_22710), .b(g62430_sb), .o(n_6738) );
in01f06 FE_RC_683_0 ( .a(FE_RN_458_0), .o(n_10595) );
na02f06 FE_RC_684_0 ( .a(n_8867), .b(n_15453), .o(FE_RN_458_0) );
na02f08 FE_RC_686_0 ( .a(n_8863), .b(n_16579), .o(FE_RN_459_0) );
no02f40 FE_RC_688_0 ( .a(n_15371), .b(n_4853), .o(FE_RN_460_0) );
na02f80 FE_RC_689_0 ( .a(FE_RN_460_0), .b(n_4815), .o(n_16435) );
in01f10 FE_RC_68_0 ( .a(n_16307), .o(FE_RN_36_0) );
in01f02 FE_RC_693_0 ( .a(n_10855), .o(FE_RN_463_0) );
in01f02 FE_RC_694_0 ( .a(n_11715), .o(FE_RN_464_0) );
no02f04 FE_RC_695_0 ( .a(FE_RN_463_0), .b(FE_RN_464_0), .o(FE_RN_465_0) );
in01f02 FE_RC_697_0 ( .a(n_10230), .o(FE_RN_466_0) );
in01f02 FE_RC_698_0 ( .a(n_10768), .o(FE_RN_467_0) );
no02f02 FE_RC_699_0 ( .a(FE_RN_466_0), .b(FE_RN_467_0), .o(FE_RN_468_0) );
in01f06 FE_RC_69_0 ( .a(n_16309), .o(FE_RN_37_0) );
na02m02 TIMEBOOST_cell_39625 ( .a(TIMEBOOST_net_11424), .b(g63436_sb), .o(n_4623) );
in01f02 FE_RC_701_0 ( .a(n_10679), .o(FE_RN_469_0) );
in01f02 FE_RC_702_0 ( .a(n_10681), .o(FE_RN_470_0) );
no02f02 FE_RC_703_0 ( .a(FE_RN_469_0), .b(FE_RN_470_0), .o(FE_RN_471_0) );
na02f02 TIMEBOOST_cell_50931 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_409), .b(g54190_sb), .o(TIMEBOOST_net_15683) );
in01f02 FE_RC_705_0 ( .a(n_10637), .o(FE_RN_472_0) );
in01f02 FE_RC_706_0 ( .a(n_10060), .o(FE_RN_473_0) );
no02f02 FE_RC_707_0 ( .a(FE_RN_472_0), .b(FE_RN_473_0), .o(FE_RN_474_0) );
in01f02 FE_RC_709_0 ( .a(n_10905), .o(FE_RN_475_0) );
na03m02 TIMEBOOST_cell_72466 ( .a(TIMEBOOST_net_219), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q), .c(g64355_sb), .o(TIMEBOOST_net_13107) );
in01f02 FE_RC_710_0 ( .a(n_11732), .o(FE_RN_476_0) );
no02f02 FE_RC_711_0 ( .a(FE_RN_475_0), .b(FE_RN_476_0), .o(FE_RN_477_0) );
na03f02 FE_RC_712_0 ( .a(n_12569), .b(n_10904), .c(FE_RN_477_0), .o(n_12831) );
in01f02 FE_RC_713_0 ( .a(n_10981), .o(FE_RN_478_0) );
in01f02 FE_RC_714_0 ( .a(n_10758), .o(FE_RN_479_0) );
no02f02 FE_RC_715_0 ( .a(FE_RN_478_0), .b(FE_RN_479_0), .o(FE_RN_480_0) );
na02s01 TIMEBOOST_cell_39721 ( .a(TIMEBOOST_net_11472), .b(g58410_db), .o(n_9207) );
in01s01 TIMEBOOST_cell_73864 ( .a(n_7895), .o(TIMEBOOST_net_23429) );
in01f10 FE_RC_718_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_), .o(FE_RN_481_0) );
in01f10 FE_RC_720_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_), .o(FE_RN_483_0) );
oa22f08 FE_RC_721_0 ( .a(FE_OCP_RBN2225_n_16322), .b(FE_RN_481_0), .c(FE_RN_483_0), .d(n_16322), .o(n_16368) );
in01m08 FE_RC_722_0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_4__213), .o(FE_RN_484_0) );
na02m06 TIMEBOOST_cell_53457 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_124), .o(TIMEBOOST_net_16946) );
na03f02 TIMEBOOST_cell_69546 ( .a(FE_OFN1797_n_2299), .b(TIMEBOOST_net_20717), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q), .o(TIMEBOOST_net_21981) );
na03f02 FE_RC_726_0 ( .a(n_16594), .b(n_14478), .c(n_16595), .o(n_14614) );
na03f02 FE_RC_728_0 ( .a(n_14551), .b(n_14258), .c(n_14257), .o(n_14596) );
na03f02 FE_RC_729_0 ( .a(n_14426), .b(n_14543), .c(n_14427), .o(n_14588) );
na03f02 FE_RC_731_0 ( .a(n_14271), .b(n_14272), .c(n_14558), .o(n_14603) );
na03f02 FE_RC_732_0 ( .a(n_14544), .b(n_14511), .c(n_14429), .o(n_14589) );
na03f02 FE_RC_733_0 ( .a(n_14564), .b(n_14290), .c(n_14471), .o(n_14609) );
na03f02 FE_RC_736_0 ( .a(n_14301), .b(n_14480), .c(n_14569), .o(n_14613) );
na03f02 FE_RC_737_0 ( .a(n_14442), .b(n_14255), .c(n_14550), .o(n_14595) );
na03f02 FE_RC_738_0 ( .a(n_14251), .b(n_14438), .c(n_14548), .o(n_14593) );
in01f08 FE_RC_73_0 ( .a(conf_w_addr_in_931), .o(FE_RN_39_0) );
no02f02 FE_RC_742_0 ( .a(g53222_p), .b(g53223_p), .o(FE_RN_489_0) );
na02f02 FE_RC_743_0 ( .a(n_14554), .b(FE_RN_489_0), .o(n_14599) );
in01f40 FE_RC_744_0 ( .a(wishbone_slave_unit_wishbone_slave_img_wallow), .o(FE_RN_490_0) );
na02f20 FE_RC_745_0 ( .a(n_15919), .b(FE_RN_490_0), .o(n_15908) );
in01f10 FE_RC_746_0 ( .a(n_16071), .o(FE_RN_491_0) );
in01f10 FE_RC_748_0 ( .a(n_16070), .o(FE_RN_493_0) );
in01f06 FE_RC_74_0 ( .a(parchk_pci_cbe_reg_in_1236), .o(FE_RN_40_0) );
na02f06 FE_RC_751_0 ( .a(FE_OCP_RBN2280_g74996_p), .b(n_16364), .o(FE_RN_494_0) );
na03f02 FE_RC_752_0 ( .a(n_13058), .b(FE_RN_203_0), .c(n_12695), .o(n_13139) );
na04f02 FE_RC_753_0 ( .a(n_13053), .b(n_12899), .c(n_12900), .d(n_12790), .o(n_13136) );
na04f02 FE_RC_754_0 ( .a(n_13117), .b(n_12864), .c(n_12863), .d(n_12778), .o(n_13318) );
na04f04 FE_RC_755_0 ( .a(n_12779), .b(n_12866), .c(n_12867), .d(n_13044), .o(n_13128) );
na04f04 FE_RC_756_0 ( .a(n_13060), .b(n_12797), .c(n_12917), .d(n_12918), .o(n_13140) );
na04f02 FE_RC_759_0 ( .a(n_13045), .b(n_12780), .c(n_12870), .d(n_12869), .o(n_13129) );
no02f10 FE_RC_75_0 ( .a(FE_RN_40_0), .b(FE_RN_39_0), .o(FE_RN_41_0) );
na04f03 FE_RC_760_0 ( .a(n_12781), .b(n_13046), .c(n_12873), .d(n_12872), .o(n_13130) );
na04f04 FE_RC_761_0 ( .a(n_11908), .b(n_11806), .c(n_12349), .d(n_12206), .o(n_12877) );
na04f04 FE_RC_762_0 ( .a(n_12203), .b(n_11903), .c(n_11805), .d(n_12345), .o(n_12874) );
ao22f02 FE_RC_764_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q), .b(FE_OFN1734_n_16317), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q), .d(FE_OFN1739_n_11019), .o(FE_RN_496_0) );
na02m02 TIMEBOOST_cell_50368 ( .a(TIMEBOOST_net_15401), .b(g62658_sb), .o(n_6228) );
in01f02 FE_RC_766_0 ( .a(FE_RN_498_0), .o(n_12912) );
na03f10 FE_RC_76_0 ( .a(FE_RN_41_0), .b(conf_w_addr_in), .c(n_15959), .o(n_16046) );
in01f08 FE_RC_770_0 ( .a(n_8452), .o(FE_RN_500_0) );
na02m08 TIMEBOOST_cell_52947 ( .a(wishbone_slave_unit_pcim_sm_data_in_650), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q), .o(TIMEBOOST_net_16691) );
na02f02 FE_RC_772_0 ( .a(n_4699), .b(n_2963), .o(FE_RN_501_0) );
in01f02 FE_RC_773_0 ( .a(FE_RN_502_0), .o(n_7093) );
oa12f02 FE_RC_774_0 ( .a(FE_RN_501_0), .b(n_4699), .c(n_2963), .o(FE_RN_502_0) );
in01f08 FE_RC_775_0 ( .a(n_1397), .o(FE_RN_503_0) );
na04s02 TIMEBOOST_cell_72919 ( .a(TIMEBOOST_net_10354), .b(g65769_sb), .c(g61742_sb), .d(g61742_db), .o(n_8333) );
na03f02 TIMEBOOST_cell_72682 ( .a(TIMEBOOST_net_16591), .b(FE_OFN784_n_2678), .c(g65220_sb), .o(n_2667) );
in01f20 FE_RC_779_0 ( .a(FE_RN_506_0), .o(n_1679) );
na03f02 FE_RC_77_0 ( .a(n_15593), .b(n_15586), .c(n_15591), .o(n_15594) );
na02f40 FE_RC_780_0 ( .a(wbu_addr_in_252), .b(wbu_addr_in_251), .o(FE_RN_506_0) );
no02f40 FE_RC_781_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_), .o(FE_RN_507_0) );
ao12f20 FE_RC_782_0 ( .a(FE_RN_507_0), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_), .o(FE_RN_508_0) );
no02f40 FE_RC_783_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_), .o(FE_RN_509_0) );
ao12f20 FE_RC_784_0 ( .a(FE_RN_509_0), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_), .o(FE_RN_510_0) );
no02f40 FE_RC_785_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_), .o(FE_RN_511_0) );
ao12f20 FE_RC_786_0 ( .a(FE_RN_511_0), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_), .o(FE_RN_512_0) );
no02f40 FE_RC_787_0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_), .o(FE_RN_513_0) );
ao12f20 FE_RC_788_0 ( .a(FE_RN_513_0), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_), .o(FE_RN_514_0) );
na02s02 TIMEBOOST_cell_38837 ( .a(TIMEBOOST_net_11030), .b(g65892_sb), .o(n_2573) );
in01f02 FE_RC_78_0 ( .a(n_551), .o(FE_RN_42_0) );
na02f06 FE_RC_790_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(FE_RN_515_0) );
oa12f04 FE_RC_791_0 ( .a(FE_RN_515_0), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(FE_RN_516_0) );
na02f06 FE_RC_792_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(FE_RN_517_0) );
oa12f04 FE_RC_793_0 ( .a(FE_RN_517_0), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(FE_RN_518_0) );
in01f08 FE_RC_794_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_), .o(FE_RN_519_0) );
in01f02 FE_RC_795_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .o(FE_RN_520_0) );
oa22f04 FE_RC_796_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .c(FE_RN_519_0), .d(FE_RN_520_0), .o(FE_RN_521_0) );
na03f08 FE_RC_797_0 ( .a(FE_RN_516_0), .b(FE_RN_518_0), .c(FE_RN_521_0), .o(n_3334) );
in01f20 FE_RC_798_0 ( .a(FE_RN_522_0), .o(n_2809) );
na02f80 FE_RC_799_0 ( .a(pciu_am1_in_523), .b(pciu_bar1_in_385), .o(FE_RN_522_0) );
in01f04 FE_RC_79_0 ( .a(n_16690), .o(FE_RN_43_0) );
na03f80 FE_RC_800_0 ( .a(n_16942), .b(n_16635), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(n_15417) );
in01f04 FE_RC_801_0 ( .a(n_2961), .o(FE_RN_523_0) );
in01f06 FE_RC_802_0 ( .a(n_2962), .o(FE_RN_524_0) );
ao22f08 FE_RC_803_0 ( .a(FE_RN_523_0), .b(FE_RN_524_0), .c(n_2961), .d(n_2962), .o(n_4702) );
in01f04 FE_RC_804_0 ( .a(FE_OCPN1852_n_16538), .o(FE_RN_525_0) );
in01f08 FE_RC_805_0 ( .a(FE_OCPN1843_n_16033), .o(FE_RN_526_0) );
na02f08 FE_RC_806_0 ( .a(FE_RN_525_0), .b(FE_RN_526_0), .o(n_16034) );
in01f10 FE_RC_807_0 ( .a(n_15744), .o(FE_RN_527_0) );
in01f10 FE_RC_808_0 ( .a(n_15748), .o(FE_RN_528_0) );
no02f20 FE_RC_809_0 ( .a(FE_OCPN1843_n_16033), .b(FE_OCPN1852_n_16538), .o(FE_RN_529_0) );
no02f08 FE_RC_80_0 ( .a(FE_RN_43_0), .b(FE_RN_42_0), .o(FE_RN_44_0) );
na02s01 TIMEBOOST_cell_38409 ( .a(TIMEBOOST_net_10816), .b(g58037_db), .o(n_9752) );
na02m06 TIMEBOOST_cell_69059 ( .a(TIMEBOOST_net_21737), .b(g64969_sb), .o(TIMEBOOST_net_9755) );
na02m04 FE_RC_812_0 ( .a(parchk_pci_trdy_en_in), .b(n_565), .o(n_1088) );
na02f10 FE_RC_813_0 ( .a(parchk_pci_trdy_en_in), .b(n_565), .o(FE_RN_530_0) );
no02f10 FE_RC_814_0 ( .a(FE_OCP_RBN1930_parchk_pci_trdy_reg_in), .b(FE_RN_530_0), .o(n_1616) );
in01f08 FE_RC_815_0 ( .a(FE_RN_71_0), .o(FE_RN_531_0) );
in01f04 FE_RC_816_0 ( .a(n_1616), .o(FE_RN_532_0) );
no02f10 FE_RC_817_0 ( .a(FE_RN_531_0), .b(FE_RN_532_0), .o(FE_RN_533_0) );
na02m01 TIMEBOOST_cell_68840 ( .a(n_4482), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q), .o(TIMEBOOST_net_21628) );
na02f10 FE_RC_81_0 ( .a(FE_RN_44_0), .b(n_1072), .o(n_2552) );
na02f20 FE_RC_820_0 ( .a(n_16284), .b(n_16285), .o(n_16289) );
na02f04 FE_RC_821_0 ( .a(n_16284), .b(n_16285), .o(FE_OCPN1868_n_16289) );
na02f10 FE_RC_822_0 ( .a(FE_RN_535_0), .b(n_16474), .o(n_16475) );
na02f10 FE_RC_823_0 ( .a(n_16513), .b(FE_OCP_RBN1954_FE_RN_462_0), .o(FE_RN_535_0) );
in01s01 TIMEBOOST_cell_73865 ( .a(TIMEBOOST_net_23429), .o(TIMEBOOST_net_23430) );
na02m02 TIMEBOOST_cell_69947 ( .a(TIMEBOOST_net_22181), .b(g52641_sb), .o(TIMEBOOST_net_5470) );
in01f20 FE_RC_828_0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .o(FE_RN_538_0) );
in01f06 FE_RC_829_0 ( .a(n_15512), .o(FE_RN_539_0) );
in01f10 FE_RC_82_0 ( .a(n_8728), .o(FE_RN_45_0) );
na02f01 TIMEBOOST_cell_26205 ( .a(conf_wb_err_addr_in_949), .b(g53940_sb), .o(TIMEBOOST_net_7207) );
na03s02 TIMEBOOST_cell_73076 ( .a(TIMEBOOST_net_22079), .b(FE_OFN1806_n_4501), .c(TIMEBOOST_net_22249), .o(TIMEBOOST_net_16780) );
na02f02 TIMEBOOST_cell_71616 ( .a(TIMEBOOST_net_13664), .b(n_12099), .o(TIMEBOOST_net_23016) );
in01s01 FE_RC_833_0 ( .a(n_7822), .o(FE_RN_541_0) );
in01f02 FE_RC_834_0 ( .a(n_12983), .o(FE_RN_542_0) );
na03f02 TIMEBOOST_cell_67996 ( .a(TIMEBOOST_net_17022), .b(FE_OFN1194_n_6935), .c(g62937_sb), .o(n_6007) );
na03f02 TIMEBOOST_cell_34957 ( .a(TIMEBOOST_net_9459), .b(FE_OFN1414_n_8567), .c(g57376_sb), .o(n_11372) );
in01f01 FE_RC_837_0 ( .a(n_13354), .o(FE_RN_544_0) );
in01f02 FE_RC_838_0 ( .a(n_12988), .o(FE_RN_545_0) );
na03m02 TIMEBOOST_cell_72645 ( .a(TIMEBOOST_net_21487), .b(g65081_sb), .c(TIMEBOOST_net_21678), .o(TIMEBOOST_net_16785) );
in01f04 FE_RC_83_0 ( .a(n_3334), .o(FE_RN_46_0) );
na03f02 TIMEBOOST_cell_66500 ( .a(TIMEBOOST_net_17100), .b(FE_OFN1312_n_6624), .c(g62948_sb), .o(n_5985) );
in01s01 FE_RC_841_0 ( .a(n_3404), .o(FE_RN_547_0) );
in01f01 FE_RC_842_0 ( .a(n_16000), .o(FE_RN_548_0) );
no02f02 FE_RC_843_0 ( .a(FE_RN_547_0), .b(FE_RN_548_0), .o(FE_RN_549_0) );
no02f02 FE_RC_844_0 ( .a(n_5724), .b(FE_RN_549_0), .o(n_7308) );
in01f80 FE_RC_846_0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_), .o(FE_RN_551_0) );
na02f80 FE_RC_847_0 ( .a(FE_OCP_RBN2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_), .b(FE_RN_551_0), .o(FE_RN_552_0) );
na03f02 TIMEBOOST_cell_34962 ( .a(TIMEBOOST_net_9465), .b(FE_OFN1377_n_8567), .c(g57096_sb), .o(n_10487) );
in01f20 FE_RC_849_0 ( .a(configuration_sync_cache_lsize_to_wb_bits_reg_2__Q), .o(FE_RN_553_0) );
no02f08 FE_RC_84_0 ( .a(FE_RN_45_0), .b(FE_RN_46_0), .o(FE_RN_47_0) );
no02f10 FE_RC_850_0 ( .a(FE_RN_553_0), .b(n_3319), .o(n_3320) );
in01f40 FE_RC_851_0 ( .a(n_681), .o(FE_RN_554_0) );
no02f40 FE_RC_852_0 ( .a(n_1200), .b(FE_RN_554_0), .o(n_16474) );
in01f20 FE_RC_854_0 ( .a(FE_RN_555_0), .o(FE_OFN993_n_15366) );
na02f40 FE_RC_855_0 ( .a(pci_target_unit_pci_target_sm_previous_frame), .b(n_15365), .o(FE_RN_555_0) );
in01f10 FE_RC_856_0 ( .a(FE_RN_556_0), .o(n_16351) );
no02f20 FE_RC_857_0 ( .a(n_16350), .b(parchk_pci_cbe_reg_in_1236), .o(FE_RN_556_0) );
in01f20 FE_RC_858_0 ( .a(FE_RN_557_0), .o(n_16307) );
na02f40 FE_RC_859_0 ( .a(n_16027), .b(n_16390), .o(FE_RN_557_0) );
in01f08 FE_RC_860_0 ( .a(n_15958), .o(FE_RN_558_0) );
na02f10 FE_RC_861_0 ( .a(FE_RN_558_0), .b(n_15959), .o(n_16388) );
no04f40 FE_RC_862_0 ( .a(pciu_cache_line_size_in_776), .b(configuration_sync_cache_lsize_to_wb_bits_reg_4__Q), .c(pciu_cache_line_size_in_777), .d(pciu_cache_line_size_in_775), .o(FE_RN_386_0) );
in01f02 FE_RC_863_0 ( .a(n_12595), .o(FE_RN_559_0) );
in01s01 FE_RC_864_0 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_789), .o(FE_RN_560_0) );
no02f02 FE_RC_865_0 ( .a(FE_RN_560_0), .b(FE_OCPN1909_n_16497), .o(FE_RN_561_0) );
ao12f02 FE_RC_866_0 ( .a(FE_RN_561_0), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q), .c(FE_OCPN1909_n_16497), .o(FE_RN_562_0) );
ao22f02 FE_RC_868_0 ( .a(configuration_pci_err_data_525), .b(FE_OFN1066_n_15808), .c(configuration_wb_err_cs_bit31_24), .d(n_16543), .o(FE_RN_564_0) );
na02f02 FE_RC_869_0 ( .a(FE_RN_564_0), .b(n_2768), .o(FE_RN_565_0) );
ao22f02 FE_RC_870_0 ( .a(configuration_status_bit8), .b(n_3248), .c(n_2815), .d(n_16000), .o(FE_RN_566_0) );
ao22f02 FE_RC_871_0 ( .a(configuration_pci_err_addr_494), .b(FE_OFN1005_n_16288), .c(configuration_pci_err_cs_bit31_24), .d(n_3252), .o(FE_RN_567_0) );
in01s01 TIMEBOOST_cell_73908 ( .a(n_4621), .o(TIMEBOOST_net_23473) );
na04f02 TIMEBOOST_cell_73587 ( .a(n_1967), .b(n_8590), .c(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .d(g59082_sb), .o(n_8591) );
ao22f02 FE_RC_874_0 ( .a(n_14927), .b(n_16810), .c(pciu_am1_in_533), .d(FE_OFN2129_n_16720), .o(FE_RN_570_0) );
ao22f02 FE_RC_875_0 ( .a(configuration_wb_err_data_594), .b(FE_OFN1070_n_15729), .c(n_2815), .d(FE_OCPN1845_n_16427), .o(FE_RN_571_0) );
na02m08 TIMEBOOST_cell_62616 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_150), .o(TIMEBOOST_net_20255) );
na02m02 TIMEBOOST_cell_44906 ( .a(TIMEBOOST_net_13347), .b(g62628_sb), .o(n_6298) );
na03f06 TIMEBOOST_cell_73077 ( .a(TIMEBOOST_net_22055), .b(FE_OFN1936_n_1781), .c(g54239_sb), .o(TIMEBOOST_net_23313) );
na03f02 TIMEBOOST_cell_34981 ( .a(TIMEBOOST_net_9515), .b(FE_OFN1382_n_8567), .c(g57397_sb), .o(n_11344) );
na03f02 TIMEBOOST_cell_34964 ( .a(TIMEBOOST_net_9435), .b(FE_OFN1388_n_8567), .c(g57534_sb), .o(n_11208) );
in01f10 FE_RC_882_0 ( .a(FE_OFN969_n_13784), .o(FE_RN_578_0) );
na02f08 FE_RC_884_0 ( .a(conf_wb_err_addr_in_965), .b(FE_OFN1620_n_1787), .o(FE_RN_580_0) );
na02f02 TIMEBOOST_cell_70839 ( .a(TIMEBOOST_net_22627), .b(g62053_sb), .o(n_7756) );
in01f01 FE_RC_886_0 ( .a(n_504), .o(FE_RN_582_0) );
in01f02 FE_RC_887_0 ( .a(FE_OFN1151_n_13249), .o(FE_RN_583_0) );
ao22f04 FE_RC_888_0 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q), .b(FE_OCPN1911_FE_OFN1152_n_13249), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_407), .d(FE_RN_583_0), .o(FE_RN_584_0) );
na02f01 TIMEBOOST_cell_49718 ( .a(TIMEBOOST_net_15076), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_13462) );
in01f02 FE_RC_88_0 ( .a(n_13754), .o(FE_RN_48_0) );
na02m02 TIMEBOOST_cell_68969 ( .a(TIMEBOOST_net_21692), .b(g65366_sb), .o(TIMEBOOST_net_12596) );
na03m02 TIMEBOOST_cell_64701 ( .a(TIMEBOOST_net_16166), .b(FE_OFN950_n_2055), .c(g65723_sb), .o(n_1748) );
in01f02 FE_RC_893_0 ( .a(FE_RN_589_0), .o(n_14345) );
na03f02 TIMEBOOST_cell_72993 ( .a(TIMEBOOST_net_23223), .b(FE_OFN1049_n_16657), .c(g64093_sb), .o(n_4062) );
in01f08 FE_RC_895_0 ( .a(n_2440), .o(FE_RN_590_0) );
in01f10 FE_RC_896_0 ( .a(FE_OFN2093_n_2301), .o(FE_RN_591_0) );
no02f10 FE_RC_897_0 ( .a(FE_RN_590_0), .b(FE_RN_591_0), .o(FE_RN_592_0) );
no02f01 FE_RC_898_0 ( .a(n_8511), .b(n_16326), .o(FE_RN_593_0) );
in01f08 FE_RC_899_0 ( .a(n_2833), .o(FE_RN_594_0) );
in01f02 FE_RC_89_0 ( .a(n_13654), .o(FE_RN_49_0) );
in01f06 FE_RC_900_0 ( .a(n_307), .o(FE_RN_595_0) );
oa22f06 FE_RC_901_0 ( .a(n_2833), .b(n_307), .c(FE_RN_594_0), .d(FE_RN_595_0), .o(FE_RN_596_0) );
in01f10 FE_RC_902_0 ( .a(n_2841), .o(FE_RN_597_0) );
in01f08 FE_RC_903_0 ( .a(n_385), .o(FE_RN_598_0) );
na02f02 TIMEBOOST_cell_68971 ( .a(TIMEBOOST_net_21693), .b(g64152_sb), .o(n_4013) );
na03m02 TIMEBOOST_cell_72369 ( .a(wishbone_slave_unit_pci_initiator_sm_timeout), .b(wishbone_slave_unit_pci_initiator_sm_transfer), .c(pciu_pciif_stop_reg_in), .o(TIMEBOOST_net_86) );
na02m04 TIMEBOOST_cell_43219 ( .a(FE_OFN642_n_4677), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q), .o(TIMEBOOST_net_12504) );
no02f04 FE_RC_907_0 ( .a(FE_RN_596_0), .b(FE_RN_601_0), .o(FE_RN_602_0) );
na02f01 FE_RC_908_0 ( .a(pciu_am1_in_540), .b(conf_pci_init_complete_out), .o(FE_RN_603_0) );
in01s04 FE_RC_909_0 ( .a(configuration_sync_command_bit0), .o(FE_RN_604_0) );
na03m02 TIMEBOOST_cell_72826 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q), .b(n_3785), .c(FE_OFN671_n_4505), .o(TIMEBOOST_net_10568) );
in01f02 FE_RC_910_0 ( .a(n_2380), .o(FE_RN_605_0) );
in01f10 FE_RC_912_0 ( .a(n_2815), .o(FE_RN_607_0) );
in01f06 FE_RC_913_0 ( .a(n_227), .o(FE_RN_608_0) );
ao22f04 FE_RC_914_0 ( .a(FE_RN_607_0), .b(FE_RN_608_0), .c(n_2815), .d(n_227), .o(FE_RN_609_0) );
na02f08 FE_RC_915_0 ( .a(n_2851), .b(n_233), .o(FE_RN_610_0) );
oa12f04 FE_RC_916_0 ( .a(FE_RN_610_0), .b(n_2851), .c(n_233), .o(FE_RN_611_0) );
na02f20 FE_RC_917_0 ( .a(n_2854), .b(n_277), .o(FE_RN_612_0) );
oa12f08 FE_RC_918_0 ( .a(FE_RN_612_0), .b(n_2854), .c(n_277), .o(FE_RN_613_0) );
na02f20 FE_RC_919_0 ( .a(n_2825), .b(n_302), .o(FE_RN_614_0) );
na04f02 TIMEBOOST_cell_73080 ( .a(TIMEBOOST_net_22062), .b(FE_OFN1807_n_4501), .c(g64870_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q), .o(TIMEBOOST_net_20979) );
oa12f08 FE_RC_920_0 ( .a(FE_RN_614_0), .b(n_2825), .c(n_302), .o(FE_RN_615_0) );
in01f10 FE_RC_921_0 ( .a(n_3592), .o(FE_RN_616_0) );
in01f06 FE_RC_922_0 ( .a(n_372), .o(FE_RN_617_0) );
oa22f04 FE_RC_923_0 ( .a(n_3592), .b(n_372), .c(FE_RN_616_0), .d(FE_RN_617_0), .o(FE_RN_618_0) );
na02f10 FE_RC_925_0 ( .a(n_2856), .b(n_336), .o(FE_RN_620_0) );
oa12f06 FE_RC_926_0 ( .a(FE_RN_620_0), .b(n_2856), .c(n_336), .o(FE_RN_621_0) );
in01f04 FE_RC_927_0 ( .a(n_3404), .o(FE_RN_622_0) );
in01f02 FE_RC_928_0 ( .a(n_290), .o(FE_RN_623_0) );
na02f02 TIMEBOOST_cell_69483 ( .a(TIMEBOOST_net_21949), .b(FE_OFN1797_n_2299), .o(n_2158) );
na03f10 FE_RC_92_0 ( .a(n_16388), .b(n_16389), .c(n_16390), .o(n_16391) );
na02m01 TIMEBOOST_cell_52330 ( .a(TIMEBOOST_net_16382), .b(FE_OFN2021_n_4778), .o(n_7187) );
na02f06 TIMEBOOST_cell_62927 ( .a(TIMEBOOST_net_20410), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_16968) );
in01f06 FE_RC_932_0 ( .a(n_2869), .o(FE_RN_627_0) );
in01f04 FE_RC_933_0 ( .a(n_287), .o(FE_RN_628_0) );
na02m04 TIMEBOOST_cell_69070 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q), .b(g65061_sb), .o(TIMEBOOST_net_21743) );
na02m01 TIMEBOOST_cell_62926 ( .a(pci_target_unit_pcit_if_strd_addr_in_701), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65), .o(TIMEBOOST_net_20410) );
in01f10 FE_RC_937_0 ( .a(n_15598), .o(FE_RN_632_0) );
in01f08 FE_RC_938_0 ( .a(n_360), .o(FE_RN_633_0) );
na02m01 TIMEBOOST_cell_52861 ( .a(TIMEBOOST_net_12783), .b(FE_OFN577_n_9902), .o(TIMEBOOST_net_16648) );
in01f02 FE_RC_93_0 ( .a(n_3365), .o(FE_RN_51_0) );
in01s01 TIMEBOOST_cell_31889 ( .a(conf_wb_err_addr_in_946), .o(TIMEBOOST_net_10053) );
in01f10 FE_RC_942_0 ( .a(n_2866), .o(FE_RN_637_0) );
in01f04 FE_RC_943_0 ( .a(n_300), .o(FE_RN_638_0) );
in01f10 FE_RC_947_0 ( .a(n_2809), .o(FE_RN_642_0) );
in01f10 FE_RC_948_0 ( .a(n_413), .o(FE_RN_643_0) );
na02f10 FE_RC_949_0 ( .a(FE_RN_643_0), .b(FE_RN_642_0), .o(FE_RN_644_0) );
in01f02 FE_RC_94_0 ( .a(n_3046), .o(FE_RN_52_0) );
in01f04 FE_RC_950_0 ( .a(n_2809), .o(FE_RN_645_0) );
in01f04 FE_RC_951_0 ( .a(n_413), .o(FE_RN_646_0) );
oa12f08 FE_RC_952_0 ( .a(FE_RN_644_0), .b(FE_RN_645_0), .c(FE_RN_646_0), .o(FE_RN_647_0) );
in01f10 FE_RC_953_0 ( .a(n_2831), .o(FE_RN_648_0) );
in01f10 FE_RC_954_0 ( .a(n_303), .o(FE_RN_649_0) );
na02f10 FE_RC_955_0 ( .a(FE_RN_648_0), .b(FE_RN_649_0), .o(FE_RN_650_0) );
in01f04 FE_RC_956_0 ( .a(n_2831), .o(FE_RN_651_0) );
oa12f08 FE_RC_958_0 ( .a(FE_RN_650_0), .b(FE_RN_651_0), .c(FE_RN_649_0), .o(FE_RN_653_0) );
in01f10 FE_RC_959_0 ( .a(n_2812), .o(FE_RN_654_0) );
no02f02 FE_RC_95_0 ( .a(FE_RN_51_0), .b(FE_RN_52_0), .o(FE_RN_53_0) );
in01f10 FE_RC_960_0 ( .a(n_389), .o(FE_RN_655_0) );
na02f10 FE_RC_961_0 ( .a(FE_RN_654_0), .b(FE_RN_655_0), .o(FE_RN_656_0) );
in01f04 FE_RC_962_0 ( .a(n_2812), .o(FE_RN_657_0) );
oa12f08 FE_RC_964_0 ( .a(FE_RN_656_0), .b(FE_RN_657_0), .c(FE_RN_655_0), .o(FE_RN_659_0) );
in01f10 FE_RC_965_0 ( .a(n_16428), .o(FE_RN_660_0) );
in01f10 FE_RC_966_0 ( .a(n_297), .o(FE_RN_661_0) );
na02f10 FE_RC_967_0 ( .a(FE_RN_660_0), .b(FE_RN_661_0), .o(FE_RN_662_0) );
in01f04 FE_RC_968_0 ( .a(n_16428), .o(FE_RN_663_0) );
na02f02 FE_RC_96_0 ( .a(n_7697), .b(FE_RN_53_0), .o(n_8488) );
oa12f08 FE_RC_970_0 ( .a(FE_RN_662_0), .b(FE_RN_663_0), .c(FE_RN_661_0), .o(FE_RN_665_0) );
na02f02 TIMEBOOST_cell_70863 ( .a(TIMEBOOST_net_22639), .b(g62831_sb), .o(n_5313) );
in01f10 FE_RC_972_0 ( .a(n_231), .o(FE_RN_667_0) );
in01f10 FE_RC_973_0 ( .a(n_2818), .o(FE_RN_668_0) );
no02f10 FE_RC_974_0 ( .a(FE_RN_667_0), .b(FE_RN_668_0), .o(FE_RN_669_0) );
no02f01 FE_RC_975_0 ( .a(n_2822), .b(n_439), .o(FE_RN_670_0) );
in01f08 FE_RC_977_0 ( .a(n_439), .o(FE_RN_672_0) );
in01f08 FE_RC_978_0 ( .a(n_2822), .o(FE_RN_673_0) );
no02f08 FE_RC_979_0 ( .a(FE_RN_672_0), .b(FE_RN_673_0), .o(FE_RN_674_0) );
na02m40 TIMEBOOST_cell_69470 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_796), .o(TIMEBOOST_net_21943) );
na02s01 TIMEBOOST_cell_31087 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_9648) );
in01f06 FE_RC_982_0 ( .a(n_376), .o(FE_RN_677_0) );
in01f08 FE_RC_983_0 ( .a(n_2844), .o(FE_RN_678_0) );
na02s01 TIMEBOOST_cell_63058 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q), .o(TIMEBOOST_net_20476) );
in01f04 FE_RC_985_0 ( .a(n_298), .o(FE_RN_680_0) );
in01f08 FE_RC_986_0 ( .a(n_2838), .o(FE_RN_681_0) );
oa22f04 FE_RC_987_0 ( .a(n_298), .b(n_2838), .c(FE_RN_680_0), .d(FE_RN_681_0), .o(FE_RN_682_0) );
na03f06 TIMEBOOST_cell_33464 ( .a(TIMEBOOST_net_9127), .b(g63138_sb), .c(FE_OFN1129_g64577_p), .o(n_4973) );
na02f02 FE_RC_989_0 ( .a(FE_RN_675_0), .b(FE_RN_683_0), .o(FE_RN_684_0) );
in01f03 FE_RC_98_0 ( .a(n_15798), .o(FE_RN_55_0) );
in01f10 FE_RC_990_0 ( .a(n_2864), .o(FE_RN_685_0) );
in01f06 FE_RC_991_0 ( .a(n_436), .o(FE_RN_686_0) );
na04f80 TIMEBOOST_cell_72451 ( .a(g58790_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q), .c(FE_OFN2055_n_8831), .d(wbu_addr_in_279), .o(n_9832) );
na02f10 FE_RC_993_0 ( .a(n_204), .b(n_2828), .o(FE_RN_688_0) );
oa12f06 FE_RC_994_0 ( .a(FE_RN_688_0), .b(n_2828), .c(n_204), .o(FE_RN_689_0) );
in01f20 FE_RC_998_0 ( .a(n_357), .o(FE_RN_693_0) );
na02f20 FE_RC_999_0 ( .a(FE_RN_695_0), .b(FE_RN_693_0), .o(FE_RN_694_0) );
no02f06 FE_RC_99_0 ( .a(FE_RN_55_0), .b(parchk_pci_trdy_reg_in), .o(FE_RN_56_0) );
ms00f80 configuration_cache_line_size_reg_reg_0__u0 ( .ck(ispd_clk), .d(n_7598), .o(configuration_cache_line_size_reg) );
ms00f80 configuration_cache_line_size_reg_reg_1__u0 ( .ck(ispd_clk), .d(n_7596), .o(configuration_cache_line_size_reg_2996) );
ms00f80 configuration_cache_line_size_reg_reg_2__u0 ( .ck(ispd_clk), .d(n_7595), .o(wbu_cache_line_size_in_206) );
ms00f80 configuration_cache_line_size_reg_reg_3__u0 ( .ck(ispd_clk), .d(n_8437), .o(wbu_cache_line_size_in_207) );
ms00f80 configuration_cache_line_size_reg_reg_4__u0 ( .ck(ispd_clk), .d(n_8436), .o(wbu_cache_line_size_in_208) );
ms00f80 configuration_cache_line_size_reg_reg_5__u0 ( .ck(ispd_clk), .d(n_8434), .o(wbu_cache_line_size_in_209) );
ms00f80 configuration_cache_line_size_reg_reg_6__u0 ( .ck(ispd_clk), .d(n_7590), .o(wbu_cache_line_size_in_210) );
ms00f80 configuration_cache_line_size_reg_reg_7__u0 ( .ck(ispd_clk), .d(n_8433), .o(wbu_cache_line_size_in_211) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_206), .o(configuration_meta_cache_lsize_to_wb_bits) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_207), .o(configuration_meta_cache_lsize_to_wb_bits_926) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_208), .o(configuration_meta_cache_lsize_to_wb_bits_927) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_3__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_209), .o(configuration_meta_cache_lsize_to_wb_bits_928) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_4__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_210), .o(configuration_meta_cache_lsize_to_wb_bits_929) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_5__u0 ( .ck(ispd_clk), .d(wbu_cache_line_size_in_211), .o(configuration_meta_cache_lsize_to_wb_bits_930) );
ms00f80 configuration_cache_lsize_to_wb_bits_sync_sync_data_out_reg_6__u0 ( .ck(ispd_clk), .d(n_1625), .o(configuration_meta_cache_lsize_to_wb_bits_931) );
ms00f80 configuration_command_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(n_8456), .o(configuration_sync_command_bit0) );
ms00f80 configuration_command_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_8455), .o(configuration_sync_command_bit1) );
ms00f80 configuration_command_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(n_8454), .o(configuration_command_bit) );
ms00f80 configuration_command_bit6_reg_u0 ( .ck(ispd_clk), .d(n_8453), .o(configuration_sync_command_bit6) );
ms00f80 configuration_command_bit8_reg_u0 ( .ck(ispd_clk), .d(n_8464), .o(configuration_sync_command_bit8) );
ms00f80 configuration_command_bit_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_command_bit), .o(configuration_meta_command_bit) );
ms00f80 configuration_i_wb_init_complete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(FE_OFN992_n_2373), .o(configuration_sync_init_complete) );
ms00f80 configuration_icr_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(n_7820), .o(configuration_icr_bit2_0) );
ms00f80 configuration_icr_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_7819), .o(configuration_icr_bit_2961) );
ms00f80 configuration_icr_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(n_7817), .o(configuration_icr_bit_2967) );
ms00f80 configuration_icr_bit31_reg_u0 ( .ck(ispd_clk), .d(n_7627), .o(pci_resi_conf_soft_res_in) );
ms00f80 configuration_init_complete_reg_u0 ( .ck(ispd_clk), .d(n_1385), .o(conf_pci_init_complete_out) );
ms00f80 configuration_int_pin_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23396), .o(configuration_int_meta) );
ms00f80 configuration_interrupt_line_reg_0__u0 ( .ck(ispd_clk), .d(n_8463), .o(configuration_interrupt_line) );
ms00f80 configuration_interrupt_line_reg_1__u0 ( .ck(ispd_clk), .d(n_8462), .o(configuration_interrupt_line_37) );
ms00f80 configuration_interrupt_line_reg_2__u0 ( .ck(ispd_clk), .d(n_8461), .o(configuration_interrupt_line_38) );
ms00f80 configuration_interrupt_line_reg_3__u0 ( .ck(ispd_clk), .d(n_8442), .o(configuration_interrupt_line_39) );
ms00f80 configuration_interrupt_line_reg_4__u0 ( .ck(ispd_clk), .d(n_8441), .o(configuration_interrupt_line_40) );
ms00f80 configuration_interrupt_line_reg_5__u0 ( .ck(ispd_clk), .d(n_8439), .o(configuration_interrupt_line_41) );
ms00f80 configuration_interrupt_line_reg_6__u0 ( .ck(ispd_clk), .d(n_8457), .o(configuration_interrupt_line_42) );
ms00f80 configuration_interrupt_line_reg_7__u0 ( .ck(ispd_clk), .d(n_8438), .o(configuration_interrupt_line_43) );
ms00f80 configuration_interrupt_out_reg_u0 ( .ck(ispd_clk), .d(configuration_int_meta), .o(configuration_interrupt_out_reg_Q) );
in01s01 configuration_interrupt_out_reg_u1 ( .a(configuration_interrupt_out_reg_Q), .o(pci_inti_conf_int_in) );
ms00f80 configuration_isr_bit0_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_536), .o(configuration_isr_bit_1461) );
ms00f80 configuration_isr_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(configuration_isr_bit_1461), .o(configuration_isr_bit_631) );
ms00f80 configuration_isr_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_8508), .o(configuration_isr_bit_2975) );
ms00f80 configuration_isr_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(configuration_isr_bit_1457), .o(configuration_isr_bit_618) );
ms00f80 configuration_isr_bit2_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_1084), .o(configuration_isr_bit_1457) );
ms00f80 configuration_latency_timer_reg_0__u0 ( .ck(ispd_clk), .d(n_7607), .o(wbu_latency_tim_val_in) );
ms00f80 configuration_latency_timer_reg_1__u0 ( .ck(ispd_clk), .d(n_7606), .o(wbu_latency_tim_val_in_243) );
ms00f80 configuration_latency_timer_reg_2__u0 ( .ck(ispd_clk), .d(n_7605), .o(wbu_latency_tim_val_in_244) );
ms00f80 configuration_latency_timer_reg_3__u0 ( .ck(ispd_clk), .d(n_7604), .o(wbu_latency_tim_val_in_245) );
ms00f80 configuration_latency_timer_reg_4__u0 ( .ck(ispd_clk), .d(n_7602), .o(wbu_latency_tim_val_in_246) );
ms00f80 configuration_latency_timer_reg_5__u0 ( .ck(ispd_clk), .d(n_7601), .o(wbu_latency_tim_val_in_247) );
ms00f80 configuration_latency_timer_reg_6__u0 ( .ck(ispd_clk), .d(n_7600), .o(wbu_latency_tim_val_in_248) );
ms00f80 configuration_latency_timer_reg_7__u0 ( .ck(ispd_clk), .d(n_7599), .o(wbu_latency_tim_val_in_249) );
ms00f80 configuration_pci_am1_reg_10__u0 ( .ck(ispd_clk), .d(n_7453), .o(pciu_am1_in_519) );
ms00f80 configuration_pci_am1_reg_11__u0 ( .ck(ispd_clk), .d(n_7452), .o(pciu_am1_in_520) );
ms00f80 configuration_pci_am1_reg_12__u0 ( .ck(ispd_clk), .d(n_7451), .o(pciu_am1_in_521) );
ms00f80 configuration_pci_am1_reg_13__u0 ( .ck(ispd_clk), .d(n_7450), .o(pciu_am1_in_522) );
ms00f80 configuration_pci_am1_reg_14__u0 ( .ck(ispd_clk), .d(n_7449), .o(pciu_am1_in_523) );
ms00f80 configuration_pci_am1_reg_15__u0 ( .ck(ispd_clk), .d(n_7448), .o(pciu_am1_in_524) );
ms00f80 configuration_pci_am1_reg_16__u0 ( .ck(ispd_clk), .d(n_7447), .o(pciu_am1_in_525) );
ms00f80 configuration_pci_am1_reg_17__u0 ( .ck(ispd_clk), .d(n_7446), .o(pciu_am1_in_526) );
ms00f80 configuration_pci_am1_reg_18__u0 ( .ck(ispd_clk), .d(n_7445), .o(pciu_am1_in_527) );
ms00f80 configuration_pci_am1_reg_19__u0 ( .ck(ispd_clk), .d(n_7433), .o(pciu_am1_in_528) );
ms00f80 configuration_pci_am1_reg_20__u0 ( .ck(ispd_clk), .d(n_7444), .o(pciu_am1_in_529) );
ms00f80 configuration_pci_am1_reg_21__u0 ( .ck(ispd_clk), .d(n_7443), .o(pciu_am1_in_530) );
ms00f80 configuration_pci_am1_reg_22__u0 ( .ck(ispd_clk), .d(n_7458), .o(pciu_am1_in_531) );
ms00f80 configuration_pci_am1_reg_23__u0 ( .ck(ispd_clk), .d(n_7439), .o(pciu_am1_in_532) );
ms00f80 configuration_pci_am1_reg_24__u0 ( .ck(ispd_clk), .d(n_7436), .o(pciu_am1_in_533) );
ms00f80 configuration_pci_am1_reg_25__u0 ( .ck(ispd_clk), .d(n_7435), .o(pciu_am1_in_534) );
ms00f80 configuration_pci_am1_reg_26__u0 ( .ck(ispd_clk), .d(n_7456), .o(pciu_am1_in_535) );
ms00f80 configuration_pci_am1_reg_27__u0 ( .ck(ispd_clk), .d(n_7432), .o(pciu_am1_in_536) );
ms00f80 configuration_pci_am1_reg_28__u0 ( .ck(ispd_clk), .d(n_7431), .o(pciu_am1_in_537) );
ms00f80 configuration_pci_am1_reg_29__u0 ( .ck(ispd_clk), .d(n_7470), .o(pciu_am1_in_538) );
ms00f80 configuration_pci_am1_reg_30__u0 ( .ck(ispd_clk), .d(n_7464), .o(pciu_am1_in_539) );
ms00f80 configuration_pci_am1_reg_31__u0 ( .ck(ispd_clk), .d(n_7430), .o(pciu_am1_in_540) );
ms00f80 configuration_pci_am1_reg_8__u0 ( .ck(ispd_clk), .d(n_7460), .o(pciu_am1_in) );
ms00f80 configuration_pci_am1_reg_9__u0 ( .ck(ispd_clk), .d(n_7429), .o(pciu_am1_in_518) );
ms00f80 configuration_pci_ba0_bit31_8_reg_12__u0 ( .ck(ispd_clk), .d(n_7594), .o(pciu_bar0_in) );
ms00f80 configuration_pci_ba0_bit31_8_reg_13__u0 ( .ck(ispd_clk), .d(n_7593), .o(pciu_bar0_in_361) );
ms00f80 configuration_pci_ba0_bit31_8_reg_14__u0 ( .ck(ispd_clk), .d(n_7592), .o(pciu_bar0_in_362) );
ms00f80 configuration_pci_ba0_bit31_8_reg_15__u0 ( .ck(ispd_clk), .d(n_7597), .o(pciu_bar0_in_363) );
ms00f80 configuration_pci_ba0_bit31_8_reg_16__u0 ( .ck(ispd_clk), .d(n_7603), .o(pciu_bar0_in_364) );
ms00f80 configuration_pci_ba0_bit31_8_reg_17__u0 ( .ck(ispd_clk), .d(n_7589), .o(pciu_bar0_in_365) );
ms00f80 configuration_pci_ba0_bit31_8_reg_18__u0 ( .ck(ispd_clk), .d(n_7591), .o(pciu_bar0_in_366) );
ms00f80 configuration_pci_ba0_bit31_8_reg_19__u0 ( .ck(ispd_clk), .d(n_7588), .o(pciu_bar0_in_367) );
ms00f80 configuration_pci_ba0_bit31_8_reg_20__u0 ( .ck(ispd_clk), .d(n_7587), .o(pciu_bar0_in_368) );
ms00f80 configuration_pci_ba0_bit31_8_reg_21__u0 ( .ck(ispd_clk), .d(n_7586), .o(pciu_bar0_in_369) );
ms00f80 configuration_pci_ba0_bit31_8_reg_22__u0 ( .ck(ispd_clk), .d(n_7585), .o(pciu_bar0_in_370) );
ms00f80 configuration_pci_ba0_bit31_8_reg_23__u0 ( .ck(ispd_clk), .d(n_7584), .o(pciu_bar0_in_371) );
ms00f80 configuration_pci_ba0_bit31_8_reg_24__u0 ( .ck(ispd_clk), .d(n_7583), .o(pciu_bar0_in_372) );
ms00f80 configuration_pci_ba0_bit31_8_reg_25__u0 ( .ck(ispd_clk), .d(n_7582), .o(pciu_bar0_in_373) );
ms00f80 configuration_pci_ba0_bit31_8_reg_26__u0 ( .ck(ispd_clk), .d(n_7581), .o(pciu_bar0_in_374) );
ms00f80 configuration_pci_ba0_bit31_8_reg_27__u0 ( .ck(ispd_clk), .d(n_7580), .o(pciu_bar0_in_375) );
ms00f80 configuration_pci_ba0_bit31_8_reg_28__u0 ( .ck(ispd_clk), .d(n_7579), .o(pciu_bar0_in_376) );
ms00f80 configuration_pci_ba0_bit31_8_reg_29__u0 ( .ck(ispd_clk), .d(n_7578), .o(pciu_bar0_in_377) );
ms00f80 configuration_pci_ba0_bit31_8_reg_30__u0 ( .ck(ispd_clk), .d(n_7577), .o(pciu_bar0_in_378) );
ms00f80 configuration_pci_ba0_bit31_8_reg_31__u0 ( .ck(ispd_clk), .d(n_7576), .o(pciu_bar0_in_379) );
ms00f80 configuration_pci_ba1_bit31_8_reg_10__u0 ( .ck(ispd_clk), .d(n_7483), .o(pciu_bar1_in_381) );
ms00f80 configuration_pci_ba1_bit31_8_reg_11__u0 ( .ck(ispd_clk), .d(n_7482), .o(pciu_bar1_in_382) );
ms00f80 configuration_pci_ba1_bit31_8_reg_12__u0 ( .ck(ispd_clk), .d(n_7481), .o(pciu_bar1_in_383) );
ms00f80 configuration_pci_ba1_bit31_8_reg_13__u0 ( .ck(ispd_clk), .d(n_7480), .o(pciu_bar1_in_384) );
ms00f80 configuration_pci_ba1_bit31_8_reg_14__u0 ( .ck(ispd_clk), .d(n_7479), .o(pciu_bar1_in_385) );
ms00f80 configuration_pci_ba1_bit31_8_reg_15__u0 ( .ck(ispd_clk), .d(n_7478), .o(pciu_bar1_in_386) );
ms00f80 configuration_pci_ba1_bit31_8_reg_16__u0 ( .ck(ispd_clk), .d(n_7477), .o(pciu_bar1_in_387) );
ms00f80 configuration_pci_ba1_bit31_8_reg_17__u0 ( .ck(ispd_clk), .d(n_7476), .o(pciu_bar1_in_388) );
ms00f80 configuration_pci_ba1_bit31_8_reg_18__u0 ( .ck(ispd_clk), .d(n_7500), .o(pciu_bar1_in_389) );
ms00f80 configuration_pci_ba1_bit31_8_reg_19__u0 ( .ck(ispd_clk), .d(n_7499), .o(pciu_bar1_in_390) );
ms00f80 configuration_pci_ba1_bit31_8_reg_20__u0 ( .ck(ispd_clk), .d(n_7497), .o(pciu_bar1_in_391) );
ms00f80 configuration_pci_ba1_bit31_8_reg_21__u0 ( .ck(ispd_clk), .d(n_7495), .o(pciu_bar1_in_392) );
ms00f80 configuration_pci_ba1_bit31_8_reg_22__u0 ( .ck(ispd_clk), .d(n_7496), .o(pciu_bar1_in_393) );
ms00f80 configuration_pci_ba1_bit31_8_reg_23__u0 ( .ck(ispd_clk), .d(n_7494), .o(pciu_bar1_in_394) );
ms00f80 configuration_pci_ba1_bit31_8_reg_24__u0 ( .ck(ispd_clk), .d(n_7493), .o(pciu_bar1_in_395) );
ms00f80 configuration_pci_ba1_bit31_8_reg_25__u0 ( .ck(ispd_clk), .d(n_7492), .o(pciu_bar1_in_396) );
ms00f80 configuration_pci_ba1_bit31_8_reg_26__u0 ( .ck(ispd_clk), .d(n_7491), .o(pciu_bar1_in_397) );
ms00f80 configuration_pci_ba1_bit31_8_reg_27__u0 ( .ck(ispd_clk), .d(n_7490), .o(pciu_bar1_in_398) );
ms00f80 configuration_pci_ba1_bit31_8_reg_28__u0 ( .ck(ispd_clk), .d(n_7489), .o(pciu_bar1_in_399) );
ms00f80 configuration_pci_ba1_bit31_8_reg_29__u0 ( .ck(ispd_clk), .d(n_7488), .o(pciu_bar1_in_400) );
ms00f80 configuration_pci_ba1_bit31_8_reg_30__u0 ( .ck(ispd_clk), .d(n_7487), .o(pciu_bar1_in_401) );
ms00f80 configuration_pci_ba1_bit31_8_reg_31__u0 ( .ck(ispd_clk), .d(n_7486), .o(pciu_bar1_in_402) );
ms00f80 configuration_pci_ba1_bit31_8_reg_8__u0 ( .ck(ispd_clk), .d(n_7484), .o(pciu_bar1_in) );
ms00f80 configuration_pci_ba1_bit31_8_reg_9__u0 ( .ck(ispd_clk), .d(n_7485), .o(pciu_bar1_in_380) );
ms00f80 configuration_pci_err_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_4851), .o(configuration_pci_err_addr) );
ms00f80 configuration_pci_err_addr_reg_10__u0 ( .ck(ispd_clk), .d(n_4849), .o(configuration_pci_err_addr_480) );
ms00f80 configuration_pci_err_addr_reg_11__u0 ( .ck(ispd_clk), .d(n_4848), .o(configuration_pci_err_addr_481) );
ms00f80 configuration_pci_err_addr_reg_12__u0 ( .ck(ispd_clk), .d(n_4847), .o(configuration_pci_err_addr_482) );
ms00f80 configuration_pci_err_addr_reg_13__u0 ( .ck(ispd_clk), .d(n_4846), .o(configuration_pci_err_addr_483) );
ms00f80 configuration_pci_err_addr_reg_14__u0 ( .ck(ispd_clk), .d(n_4845), .o(configuration_pci_err_addr_484) );
ms00f80 configuration_pci_err_addr_reg_15__u0 ( .ck(ispd_clk), .d(n_4844), .o(configuration_pci_err_addr_485) );
ms00f80 configuration_pci_err_addr_reg_16__u0 ( .ck(ispd_clk), .d(n_4843), .o(configuration_pci_err_addr_486) );
ms00f80 configuration_pci_err_addr_reg_17__u0 ( .ck(ispd_clk), .d(n_4842), .o(configuration_pci_err_addr_487) );
ms00f80 configuration_pci_err_addr_reg_18__u0 ( .ck(ispd_clk), .d(n_4841), .o(configuration_pci_err_addr_488) );
ms00f80 configuration_pci_err_addr_reg_19__u0 ( .ck(ispd_clk), .d(n_4840), .o(configuration_pci_err_addr_489) );
ms00f80 configuration_pci_err_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_4839), .o(configuration_pci_err_addr_471) );
ms00f80 configuration_pci_err_addr_reg_20__u0 ( .ck(ispd_clk), .d(n_4838), .o(configuration_pci_err_addr_490) );
ms00f80 configuration_pci_err_addr_reg_21__u0 ( .ck(ispd_clk), .d(n_4837), .o(configuration_pci_err_addr_491) );
ms00f80 configuration_pci_err_addr_reg_22__u0 ( .ck(ispd_clk), .d(n_4836), .o(configuration_pci_err_addr_492) );
ms00f80 configuration_pci_err_addr_reg_23__u0 ( .ck(ispd_clk), .d(n_4835), .o(configuration_pci_err_addr_493) );
ms00f80 configuration_pci_err_addr_reg_24__u0 ( .ck(ispd_clk), .d(n_4834), .o(configuration_pci_err_addr_494) );
ms00f80 configuration_pci_err_addr_reg_25__u0 ( .ck(ispd_clk), .d(n_4833), .o(configuration_pci_err_addr_495) );
ms00f80 configuration_pci_err_addr_reg_26__u0 ( .ck(ispd_clk), .d(n_4831), .o(configuration_pci_err_addr_496) );
ms00f80 configuration_pci_err_addr_reg_27__u0 ( .ck(ispd_clk), .d(n_4832), .o(configuration_pci_err_addr_497) );
ms00f80 configuration_pci_err_addr_reg_28__u0 ( .ck(ispd_clk), .d(n_4830), .o(configuration_pci_err_addr_498) );
ms00f80 configuration_pci_err_addr_reg_29__u0 ( .ck(ispd_clk), .d(n_4828), .o(configuration_pci_err_addr_499) );
ms00f80 configuration_pci_err_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_5712), .o(configuration_pci_err_addr_472) );
ms00f80 configuration_pci_err_addr_reg_30__u0 ( .ck(ispd_clk), .d(n_5710), .o(configuration_pci_err_addr_500) );
ms00f80 configuration_pci_err_addr_reg_31__u0 ( .ck(ispd_clk), .d(n_5709), .o(configuration_pci_err_addr_501) );
ms00f80 configuration_pci_err_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_5708), .o(configuration_pci_err_addr_473) );
ms00f80 configuration_pci_err_addr_reg_4__u0 ( .ck(ispd_clk), .d(n_5707), .o(configuration_pci_err_addr_474) );
ms00f80 configuration_pci_err_addr_reg_5__u0 ( .ck(ispd_clk), .d(n_5705), .o(configuration_pci_err_addr_475) );
ms00f80 configuration_pci_err_addr_reg_6__u0 ( .ck(ispd_clk), .d(n_5704), .o(configuration_pci_err_addr_476) );
ms00f80 configuration_pci_err_addr_reg_7__u0 ( .ck(ispd_clk), .d(n_5703), .o(configuration_pci_err_addr_477) );
ms00f80 configuration_pci_err_addr_reg_8__u0 ( .ck(ispd_clk), .d(n_5702), .o(configuration_pci_err_addr_478) );
ms00f80 configuration_pci_err_addr_reg_9__u0 ( .ck(ispd_clk), .d(n_5701), .o(configuration_pci_err_addr_479) );
ms00f80 configuration_pci_err_cs_bit0_reg_u0 ( .ck(ispd_clk), .d(n_8519), .o(configuration_pci_err_cs_bit0) );
ms00f80 configuration_pci_err_cs_bit10_reg_u0 ( .ck(ispd_clk), .d(n_4873), .o(configuration_pci_err_cs_bit10) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_24__u0 ( .ck(ispd_clk), .d(n_5699), .o(configuration_pci_err_cs_bit31_24) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_25__u0 ( .ck(ispd_clk), .d(n_5696), .o(configuration_pci_err_cs_bit_464) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_26__u0 ( .ck(ispd_clk), .d(n_5694), .o(configuration_pci_err_cs_bit_465) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_27__u0 ( .ck(ispd_clk), .d(n_5691), .o(configuration_pci_err_cs_bit_466) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_28__u0 ( .ck(ispd_clk), .d(n_4867), .o(configuration_pci_err_cs_bit_467) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_29__u0 ( .ck(ispd_clk), .d(n_4866), .o(configuration_pci_err_cs_bit_468) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_30__u0 ( .ck(ispd_clk), .d(n_4864), .o(configuration_pci_err_cs_bit_469) );
ms00f80 configuration_pci_err_cs_bit31_24_reg_31__u0 ( .ck(ispd_clk), .d(n_4863), .o(configuration_pci_err_cs_bit_470) );
ms00f80 configuration_pci_err_cs_bit8_reg_u0 ( .ck(ispd_clk), .d(configuration_meta_pci_err_cs_bits), .o(configuration_pci_err_cs_bit8) );
ms00f80 configuration_pci_err_cs_bit9_reg_u0 ( .ck(ispd_clk), .d(n_4872), .o(configuration_pci_err_cs_bit9) );
ms00f80 configuration_pci_err_cs_bits_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_736), .o(configuration_meta_pci_err_cs_bits) );
ms00f80 configuration_pci_err_data_reg_0__u0 ( .ck(ispd_clk), .d(n_5689), .o(configuration_pci_err_data) );
ms00f80 configuration_pci_err_data_reg_10__u0 ( .ck(ispd_clk), .d(n_5688), .o(configuration_pci_err_data_511) );
ms00f80 configuration_pci_err_data_reg_11__u0 ( .ck(ispd_clk), .d(n_5687), .o(configuration_pci_err_data_512) );
ms00f80 configuration_pci_err_data_reg_12__u0 ( .ck(ispd_clk), .d(n_5686), .o(configuration_pci_err_data_513) );
ms00f80 configuration_pci_err_data_reg_13__u0 ( .ck(ispd_clk), .d(n_5684), .o(configuration_pci_err_data_514) );
ms00f80 configuration_pci_err_data_reg_14__u0 ( .ck(ispd_clk), .d(n_5682), .o(configuration_pci_err_data_515) );
ms00f80 configuration_pci_err_data_reg_15__u0 ( .ck(ispd_clk), .d(n_5681), .o(configuration_pci_err_data_516) );
ms00f80 configuration_pci_err_data_reg_16__u0 ( .ck(ispd_clk), .d(n_5679), .o(configuration_pci_err_data_517) );
ms00f80 configuration_pci_err_data_reg_17__u0 ( .ck(ispd_clk), .d(n_5678), .o(configuration_pci_err_data_518) );
ms00f80 configuration_pci_err_data_reg_18__u0 ( .ck(ispd_clk), .d(n_5676), .o(configuration_pci_err_data_519) );
ms00f80 configuration_pci_err_data_reg_19__u0 ( .ck(ispd_clk), .d(n_5675), .o(configuration_pci_err_data_520) );
ms00f80 configuration_pci_err_data_reg_1__u0 ( .ck(ispd_clk), .d(n_5673), .o(configuration_pci_err_data_502) );
ms00f80 configuration_pci_err_data_reg_20__u0 ( .ck(ispd_clk), .d(n_5672), .o(configuration_pci_err_data_521) );
ms00f80 configuration_pci_err_data_reg_21__u0 ( .ck(ispd_clk), .d(n_5670), .o(configuration_pci_err_data_522) );
ms00f80 configuration_pci_err_data_reg_22__u0 ( .ck(ispd_clk), .d(n_5669), .o(configuration_pci_err_data_523) );
ms00f80 configuration_pci_err_data_reg_23__u0 ( .ck(ispd_clk), .d(n_5668), .o(configuration_pci_err_data_524) );
ms00f80 configuration_pci_err_data_reg_24__u0 ( .ck(ispd_clk), .d(n_5666), .o(configuration_pci_err_data_525) );
ms00f80 configuration_pci_err_data_reg_25__u0 ( .ck(ispd_clk), .d(n_5664), .o(configuration_pci_err_data_526) );
ms00f80 configuration_pci_err_data_reg_26__u0 ( .ck(ispd_clk), .d(n_5663), .o(configuration_pci_err_data_527) );
ms00f80 configuration_pci_err_data_reg_27__u0 ( .ck(ispd_clk), .d(n_5662), .o(configuration_pci_err_data_528) );
ms00f80 configuration_pci_err_data_reg_28__u0 ( .ck(ispd_clk), .d(n_5660), .o(configuration_pci_err_data_529) );
ms00f80 configuration_pci_err_data_reg_29__u0 ( .ck(ispd_clk), .d(n_5658), .o(configuration_pci_err_data_530) );
ms00f80 configuration_pci_err_data_reg_2__u0 ( .ck(ispd_clk), .d(n_5648), .o(configuration_pci_err_data_503) );
ms00f80 configuration_pci_err_data_reg_30__u0 ( .ck(ispd_clk), .d(n_5657), .o(configuration_pci_err_data_531) );
ms00f80 configuration_pci_err_data_reg_31__u0 ( .ck(ispd_clk), .d(n_5656), .o(configuration_pci_err_data_532) );
ms00f80 configuration_pci_err_data_reg_3__u0 ( .ck(ispd_clk), .d(n_5655), .o(configuration_pci_err_data_504) );
ms00f80 configuration_pci_err_data_reg_4__u0 ( .ck(ispd_clk), .d(n_5654), .o(configuration_pci_err_data_505) );
ms00f80 configuration_pci_err_data_reg_5__u0 ( .ck(ispd_clk), .d(n_5652), .o(configuration_pci_err_data_506) );
ms00f80 configuration_pci_err_data_reg_6__u0 ( .ck(ispd_clk), .d(n_5646), .o(configuration_pci_err_data_507) );
ms00f80 configuration_pci_err_data_reg_7__u0 ( .ck(ispd_clk), .d(n_5651), .o(configuration_pci_err_data_508) );
ms00f80 configuration_pci_err_data_reg_8__u0 ( .ck(ispd_clk), .d(n_5650), .o(configuration_pci_err_data_509) );
ms00f80 configuration_pci_err_data_reg_9__u0 ( .ck(ispd_clk), .d(n_5649), .o(configuration_pci_err_data_510) );
ms00f80 configuration_pci_img_ctrl1_bit2_1_reg_1__u0 ( .ck(ispd_clk), .d(n_8523), .o(pciu_pref_en_in_320) );
ms00f80 configuration_pci_img_ctrl1_bit2_1_reg_2__u0 ( .ck(ispd_clk), .d(n_8522), .o(n_14910) );
ms00f80 configuration_pci_ta1_reg_10__u0 ( .ck(ispd_clk), .d(n_7271), .o(n_14913) );
ms00f80 configuration_pci_ta1_reg_11__u0 ( .ck(ispd_clk), .d(n_7264), .o(n_14914) );
ms00f80 configuration_pci_ta1_reg_12__u0 ( .ck(ispd_clk), .d(n_7263), .o(n_14915) );
ms00f80 configuration_pci_ta1_reg_13__u0 ( .ck(ispd_clk), .d(n_7262), .o(n_14916) );
ms00f80 configuration_pci_ta1_reg_14__u0 ( .ck(ispd_clk), .d(n_7261), .o(n_14917) );
ms00f80 configuration_pci_ta1_reg_15__u0 ( .ck(ispd_clk), .d(n_7228), .o(n_14918) );
ms00f80 configuration_pci_ta1_reg_16__u0 ( .ck(ispd_clk), .d(n_7258), .o(n_14919) );
ms00f80 configuration_pci_ta1_reg_17__u0 ( .ck(ispd_clk), .d(n_7257), .o(n_14920) );
ms00f80 configuration_pci_ta1_reg_18__u0 ( .ck(ispd_clk), .d(n_7256), .o(n_14921) );
ms00f80 configuration_pci_ta1_reg_19__u0 ( .ck(ispd_clk), .d(n_7298), .o(n_14922) );
ms00f80 configuration_pci_ta1_reg_20__u0 ( .ck(ispd_clk), .d(n_7253), .o(n_14923) );
ms00f80 configuration_pci_ta1_reg_21__u0 ( .ck(ispd_clk), .d(n_7252), .o(n_14924) );
ms00f80 configuration_pci_ta1_reg_22__u0 ( .ck(ispd_clk), .d(n_7251), .o(n_14925) );
ms00f80 configuration_pci_ta1_reg_23__u0 ( .ck(ispd_clk), .d(n_7248), .o(n_14926) );
ms00f80 configuration_pci_ta1_reg_24__u0 ( .ck(ispd_clk), .d(n_7247), .o(n_14927) );
ms00f80 configuration_pci_ta1_reg_25__u0 ( .ck(ispd_clk), .d(n_7246), .o(n_14928) );
ms00f80 configuration_pci_ta1_reg_26__u0 ( .ck(ispd_clk), .d(n_7243), .o(n_14929) );
ms00f80 configuration_pci_ta1_reg_27__u0 ( .ck(ispd_clk), .d(n_7281), .o(n_14930) );
ms00f80 configuration_pci_ta1_reg_28__u0 ( .ck(ispd_clk), .d(n_7229), .o(n_14931) );
ms00f80 configuration_pci_ta1_reg_29__u0 ( .ck(ispd_clk), .d(n_7297), .o(n_14932) );
ms00f80 configuration_pci_ta1_reg_30__u0 ( .ck(ispd_clk), .d(n_7227), .o(n_14933) );
ms00f80 configuration_pci_ta1_reg_31__u0 ( .ck(ispd_clk), .d(n_7238), .o(n_14934) );
ms00f80 configuration_pci_ta1_reg_8__u0 ( .ck(ispd_clk), .d(n_7237), .o(n_14911) );
ms00f80 configuration_pci_ta1_reg_9__u0 ( .ck(ispd_clk), .d(n_7236), .o(n_14912) );
ms00f80 configuration_rst_inactive_reg_u0 ( .ck(ispd_clk), .d(configuration_rst_inactive_sync), .o(configuration_rst_inactive) );
ms00f80 configuration_rst_inactive_sync_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23398), .o(configuration_rst_inactive_sync) );
ms00f80 configuration_set_isr_bit2_reg_u0 ( .ck(ispd_clk), .d(n_5730), .o(configuration_set_isr_bit2_reg_Q) );
in01s01 configuration_set_isr_bit2_reg_u1 ( .a(configuration_set_isr_bit2_reg_Q), .o(configuration_set_isr_bit2) );
ms00f80 configuration_set_pci_err_cs_bit8_reg_u0 ( .ck(ispd_clk), .d(n_4695), .o(configuration_set_pci_err_cs_bit8_reg_Q) );
in01s01 configuration_set_pci_err_cs_bit8_reg_u1 ( .a(configuration_set_pci_err_cs_bit8_reg_Q), .o(configuration_set_pci_err_cs_bit8) );
ms00f80 configuration_status_bit15_11_reg_11__u0 ( .ck(ispd_clk), .d(n_8472), .o(configuration_status_bit_435) );
ms00f80 configuration_status_bit15_11_reg_12__u0 ( .ck(ispd_clk), .d(n_8509), .o(configuration_status_bit_407) );
ms00f80 configuration_status_bit15_11_reg_13__u0 ( .ck(ispd_clk), .d(n_8506), .o(configuration_status_bit_379) );
ms00f80 configuration_status_bit15_11_reg_14__u0 ( .ck(ispd_clk), .d(n_14080), .o(configuration_status_bit_351) );
ms00f80 configuration_status_bit15_11_reg_15__u0 ( .ck(ispd_clk), .d(n_14491), .o(configuration_status_bit_322) );
ms00f80 configuration_status_bit8_reg_u0 ( .ck(ispd_clk), .d(n_14901), .o(configuration_status_bit8) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_2__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits), .o(configuration_sync_cache_lsize_to_wb_bits_reg_2__Q) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_3__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_926), .o(configuration_sync_cache_lsize_to_wb_bits_reg_3__Q) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_4__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_927), .o(configuration_sync_cache_lsize_to_wb_bits_reg_4__Q) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_5__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_928), .o(pciu_cache_line_size_in_775) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_6__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_929), .o(pciu_cache_line_size_in_776) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_7__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_930), .o(pciu_cache_line_size_in_777) );
ms00f80 configuration_sync_cache_lsize_to_wb_bits_reg_8__u0 ( .ck(ispd_clk), .d(configuration_meta_cache_lsize_to_wb_bits_931), .o(pciu_cache_lsize_not_zero_in) );
ms00f80 configuration_sync_command_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_meta_command_bit), .o(configuration_sync_command_bit2) );
ms00f80 configuration_sync_isr_2_clear_delete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_sync_del_bit), .o(configuration_sync_isr_2_meta_bckp_bit) );
ms00f80 configuration_sync_isr_2_del_bit_reg_u0 ( .ck(ispd_clk), .d(n_8432), .o(configuration_sync_isr_2_del_bit_reg_Q) );
ms00f80 configuration_sync_isr_2_delayed_bckp_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_sync_bckp_bit), .o(configuration_sync_isr_2_delayed_bckp_bit_reg_Q) );
in01s01 configuration_sync_isr_2_delayed_bckp_bit_reg_u1 ( .a(configuration_sync_isr_2_delayed_bckp_bit_reg_Q), .o(configuration_sync_isr_2_delayed_bckp_bit) );
ms00f80 configuration_sync_isr_2_delayed_del_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_sync_del_bit), .o(configuration_sync_isr_2_delayed_del_bit_reg_Q) );
in01s01 configuration_sync_isr_2_delayed_del_bit_reg_u1 ( .a(configuration_sync_isr_2_delayed_del_bit_reg_Q), .o(configuration_sync_isr_2_delayed_del_bit) );
ms00f80 configuration_sync_isr_2_delete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_del_bit_reg_Q), .o(configuration_sync_isr_2_meta_del_bit) );
ms00f80 configuration_sync_isr_2_sync_bckp_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_meta_bckp_bit), .o(TIMEBOOST_net_13833) );
ms00f80 configuration_sync_isr_2_sync_del_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_isr_2_meta_del_bit), .o(configuration_sync_isr_2_sync_del_bit) );
ms00f80 configuration_sync_pci_err_cs_8_clear_delete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_sync_del_bit), .o(configuration_sync_pci_err_cs_8_meta_bckp_bit) );
ms00f80 configuration_sync_pci_err_cs_8_del_bit_reg_u0 ( .ck(ispd_clk), .d(n_8431), .o(configuration_sync_pci_err_cs_8_del_bit_reg_Q) );
ms00f80 configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_sync_bckp_bit), .o(configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_Q) );
in01s01 configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_u1 ( .a(configuration_sync_pci_err_cs_8_delayed_bckp_bit_reg_Q), .o(configuration_sync_pci_err_cs_8_delayed_bckp_bit) );
ms00f80 configuration_sync_pci_err_cs_8_delayed_del_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_sync_del_bit), .o(configuration_sync_pci_err_cs_8_delayed_del_bit_reg_Q) );
in01s01 configuration_sync_pci_err_cs_8_delayed_del_bit_reg_u1 ( .a(configuration_sync_pci_err_cs_8_delayed_del_bit_reg_Q), .o(configuration_sync_pci_err_cs_8_delayed_del_bit) );
ms00f80 configuration_sync_pci_err_cs_8_delete_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_del_bit_reg_Q), .o(configuration_sync_pci_err_cs_8_meta_del_bit) );
ms00f80 configuration_sync_pci_err_cs_8_sync_bckp_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_meta_bckp_bit), .o(TIMEBOOST_net_13835) );
ms00f80 configuration_sync_pci_err_cs_8_sync_del_bit_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_pci_err_cs_8_meta_del_bit), .o(configuration_sync_pci_err_cs_8_sync_del_bit) );
ms00f80 configuration_wb_am1_reg_31__u0 ( .ck(ispd_clk), .d(n_8542), .o(wbu_am1_in) );
ms00f80 configuration_wb_am2_reg_31__u0 ( .ck(ispd_clk), .d(n_8541), .o(wbu_am2_in) );
ms00f80 configuration_wb_ba1_bit0_reg_u0 ( .ck(ispd_clk), .d(n_8470), .o(wbu_map_in_131) );
ms00f80 configuration_wb_ba1_bit31_12_reg_31__u0 ( .ck(ispd_clk), .d(n_8469), .o(wbu_bar1_in) );
ms00f80 configuration_wb_ba2_bit0_reg_u0 ( .ck(ispd_clk), .d(n_8467), .o(wbu_map_in_132) );
ms00f80 configuration_wb_ba2_bit31_12_reg_31__u0 ( .ck(ispd_clk), .d(n_8466), .o(wbu_bar2_in) );
ms00f80 configuration_wb_err_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_5718), .o(configuration_wb_err_addr) );
ms00f80 configuration_wb_err_addr_reg_10__u0 ( .ck(ispd_clk), .d(n_5587), .o(configuration_wb_err_addr_542) );
ms00f80 configuration_wb_err_addr_reg_11__u0 ( .ck(ispd_clk), .d(n_5585), .o(configuration_wb_err_addr_543) );
ms00f80 configuration_wb_err_addr_reg_12__u0 ( .ck(ispd_clk), .d(n_5583), .o(configuration_wb_err_addr_544) );
ms00f80 configuration_wb_err_addr_reg_13__u0 ( .ck(ispd_clk), .d(n_5582), .o(configuration_wb_err_addr_545) );
ms00f80 configuration_wb_err_addr_reg_14__u0 ( .ck(ispd_clk), .d(n_5581), .o(configuration_wb_err_addr_546) );
ms00f80 configuration_wb_err_addr_reg_15__u0 ( .ck(ispd_clk), .d(n_5580), .o(configuration_wb_err_addr_547) );
ms00f80 configuration_wb_err_addr_reg_16__u0 ( .ck(ispd_clk), .d(n_5579), .o(configuration_wb_err_addr_548) );
ms00f80 configuration_wb_err_addr_reg_17__u0 ( .ck(ispd_clk), .d(n_5578), .o(configuration_wb_err_addr_549) );
ms00f80 configuration_wb_err_addr_reg_18__u0 ( .ck(ispd_clk), .d(n_5577), .o(configuration_wb_err_addr_550) );
ms00f80 configuration_wb_err_addr_reg_19__u0 ( .ck(ispd_clk), .d(n_5576), .o(configuration_wb_err_addr_551) );
ms00f80 configuration_wb_err_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_4891), .o(configuration_wb_err_addr_533) );
ms00f80 configuration_wb_err_addr_reg_20__u0 ( .ck(ispd_clk), .d(n_5575), .o(configuration_wb_err_addr_552) );
ms00f80 configuration_wb_err_addr_reg_21__u0 ( .ck(ispd_clk), .d(n_5574), .o(configuration_wb_err_addr_553) );
ms00f80 configuration_wb_err_addr_reg_22__u0 ( .ck(ispd_clk), .d(n_5573), .o(configuration_wb_err_addr_554) );
ms00f80 configuration_wb_err_addr_reg_23__u0 ( .ck(ispd_clk), .d(n_5572), .o(configuration_wb_err_addr_555) );
ms00f80 configuration_wb_err_addr_reg_24__u0 ( .ck(ispd_clk), .d(n_5571), .o(configuration_wb_err_addr_556) );
ms00f80 configuration_wb_err_addr_reg_25__u0 ( .ck(ispd_clk), .d(n_5570), .o(configuration_wb_err_addr_557) );
ms00f80 configuration_wb_err_addr_reg_26__u0 ( .ck(ispd_clk), .d(n_5569), .o(configuration_wb_err_addr_558) );
ms00f80 configuration_wb_err_addr_reg_27__u0 ( .ck(ispd_clk), .d(n_5568), .o(configuration_wb_err_addr_559) );
ms00f80 configuration_wb_err_addr_reg_28__u0 ( .ck(ispd_clk), .d(n_5567), .o(configuration_wb_err_addr_560) );
ms00f80 configuration_wb_err_addr_reg_29__u0 ( .ck(ispd_clk), .d(n_5566), .o(configuration_wb_err_addr_561) );
ms00f80 configuration_wb_err_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_5565), .o(configuration_wb_err_addr_534) );
ms00f80 configuration_wb_err_addr_reg_30__u0 ( .ck(ispd_clk), .d(n_5563), .o(configuration_wb_err_addr_562) );
ms00f80 configuration_wb_err_addr_reg_31__u0 ( .ck(ispd_clk), .d(n_5561), .o(configuration_wb_err_addr_563) );
ms00f80 configuration_wb_err_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_5559), .o(configuration_wb_err_addr_535) );
ms00f80 configuration_wb_err_addr_reg_4__u0 ( .ck(ispd_clk), .d(n_5558), .o(configuration_wb_err_addr_536) );
ms00f80 configuration_wb_err_addr_reg_5__u0 ( .ck(ispd_clk), .d(n_5557), .o(configuration_wb_err_addr_537) );
ms00f80 configuration_wb_err_addr_reg_6__u0 ( .ck(ispd_clk), .d(n_5556), .o(configuration_wb_err_addr_538) );
ms00f80 configuration_wb_err_addr_reg_7__u0 ( .ck(ispd_clk), .d(n_5555), .o(configuration_wb_err_addr_539) );
ms00f80 configuration_wb_err_addr_reg_8__u0 ( .ck(ispd_clk), .d(n_5554), .o(configuration_wb_err_addr_540) );
ms00f80 configuration_wb_err_addr_reg_9__u0 ( .ck(ispd_clk), .d(n_5553), .o(configuration_wb_err_addr_541) );
ms00f80 configuration_wb_err_cs_bit0_reg_u0 ( .ck(ispd_clk), .d(n_8518), .o(configuration_wb_err_cs_bit0) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_24__u0 ( .ck(ispd_clk), .d(n_5552), .o(configuration_wb_err_cs_bit31_24) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_25__u0 ( .ck(ispd_clk), .d(n_5639), .o(configuration_wb_err_cs_bit_564) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_26__u0 ( .ck(ispd_clk), .d(n_5638), .o(configuration_wb_err_cs_bit_565) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_27__u0 ( .ck(ispd_clk), .d(n_5637), .o(configuration_wb_err_cs_bit_566) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_28__u0 ( .ck(ispd_clk), .d(n_5636), .o(configuration_wb_err_cs_bit_567) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_29__u0 ( .ck(ispd_clk), .d(n_5635), .o(configuration_wb_err_cs_bit_568) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_30__u0 ( .ck(ispd_clk), .d(n_5634), .o(configuration_wb_err_cs_bit_569) );
ms00f80 configuration_wb_err_cs_bit31_24_reg_31__u0 ( .ck(ispd_clk), .d(n_5632), .o(configuration_wb_err_cs_bit_570) );
ms00f80 configuration_wb_err_cs_bit8_reg_u0 ( .ck(ispd_clk), .d(n_8510), .o(configuration_wb_err_cs_bit8) );
ms00f80 configuration_wb_err_cs_bit9_reg_u0 ( .ck(ispd_clk), .d(n_6218), .o(configuration_wb_err_cs_bit9) );
ms00f80 configuration_wb_err_data_reg_0__u0 ( .ck(ispd_clk), .d(n_5631), .o(configuration_wb_err_data) );
ms00f80 configuration_wb_err_data_reg_10__u0 ( .ck(ispd_clk), .d(n_5630), .o(configuration_wb_err_data_580) );
ms00f80 configuration_wb_err_data_reg_11__u0 ( .ck(ispd_clk), .d(n_5628), .o(configuration_wb_err_data_581) );
ms00f80 configuration_wb_err_data_reg_12__u0 ( .ck(ispd_clk), .d(n_5627), .o(configuration_wb_err_data_582) );
ms00f80 configuration_wb_err_data_reg_13__u0 ( .ck(ispd_clk), .d(n_5626), .o(configuration_wb_err_data_583) );
ms00f80 configuration_wb_err_data_reg_14__u0 ( .ck(ispd_clk), .d(n_5625), .o(configuration_wb_err_data_584) );
ms00f80 configuration_wb_err_data_reg_15__u0 ( .ck(ispd_clk), .d(n_5623), .o(configuration_wb_err_data_585) );
ms00f80 configuration_wb_err_data_reg_16__u0 ( .ck(ispd_clk), .d(n_5622), .o(configuration_wb_err_data_586) );
ms00f80 configuration_wb_err_data_reg_17__u0 ( .ck(ispd_clk), .d(n_5620), .o(configuration_wb_err_data_587) );
ms00f80 configuration_wb_err_data_reg_18__u0 ( .ck(ispd_clk), .d(n_5619), .o(configuration_wb_err_data_588) );
ms00f80 configuration_wb_err_data_reg_19__u0 ( .ck(ispd_clk), .d(n_5618), .o(configuration_wb_err_data_589) );
ms00f80 configuration_wb_err_data_reg_1__u0 ( .ck(ispd_clk), .d(n_5617), .o(configuration_wb_err_data_571) );
ms00f80 configuration_wb_err_data_reg_20__u0 ( .ck(ispd_clk), .d(n_5616), .o(configuration_wb_err_data_590) );
ms00f80 configuration_wb_err_data_reg_21__u0 ( .ck(ispd_clk), .d(n_5614), .o(configuration_wb_err_data_591) );
ms00f80 configuration_wb_err_data_reg_22__u0 ( .ck(ispd_clk), .d(n_5612), .o(configuration_wb_err_data_592) );
ms00f80 configuration_wb_err_data_reg_23__u0 ( .ck(ispd_clk), .d(n_5611), .o(configuration_wb_err_data_593) );
ms00f80 configuration_wb_err_data_reg_24__u0 ( .ck(ispd_clk), .d(n_5609), .o(configuration_wb_err_data_594) );
ms00f80 configuration_wb_err_data_reg_25__u0 ( .ck(ispd_clk), .d(n_5608), .o(configuration_wb_err_data_595) );
ms00f80 configuration_wb_err_data_reg_26__u0 ( .ck(ispd_clk), .d(n_5607), .o(configuration_wb_err_data_596) );
ms00f80 configuration_wb_err_data_reg_27__u0 ( .ck(ispd_clk), .d(n_5606), .o(configuration_wb_err_data_597) );
ms00f80 configuration_wb_err_data_reg_28__u0 ( .ck(ispd_clk), .d(n_5604), .o(configuration_wb_err_data_598) );
ms00f80 configuration_wb_err_data_reg_29__u0 ( .ck(ispd_clk), .d(n_5603), .o(configuration_wb_err_data_599) );
ms00f80 configuration_wb_err_data_reg_2__u0 ( .ck(ispd_clk), .d(n_5601), .o(configuration_wb_err_data_572) );
ms00f80 configuration_wb_err_data_reg_30__u0 ( .ck(ispd_clk), .d(n_5600), .o(configuration_wb_err_data_600) );
ms00f80 configuration_wb_err_data_reg_31__u0 ( .ck(ispd_clk), .d(n_5598), .o(configuration_wb_err_data_601) );
ms00f80 configuration_wb_err_data_reg_3__u0 ( .ck(ispd_clk), .d(n_5597), .o(configuration_wb_err_data_573) );
ms00f80 configuration_wb_err_data_reg_4__u0 ( .ck(ispd_clk), .d(n_5595), .o(configuration_wb_err_data_574) );
ms00f80 configuration_wb_err_data_reg_5__u0 ( .ck(ispd_clk), .d(n_5594), .o(configuration_wb_err_data_575) );
ms00f80 configuration_wb_err_data_reg_6__u0 ( .ck(ispd_clk), .d(n_5593), .o(configuration_wb_err_data_576) );
ms00f80 configuration_wb_err_data_reg_7__u0 ( .ck(ispd_clk), .d(n_5591), .o(configuration_wb_err_data_577) );
ms00f80 configuration_wb_err_data_reg_8__u0 ( .ck(ispd_clk), .d(n_5589), .o(configuration_wb_err_data_578) );
ms00f80 configuration_wb_err_data_reg_9__u0 ( .ck(ispd_clk), .d(n_5588), .o(configuration_wb_err_data_579) );
ms00f80 configuration_wb_img_ctrl1_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(n_8478), .o(wbu_mrl_en_in_141) );
ms00f80 configuration_wb_img_ctrl1_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_8474), .o(wbu_pref_en_in_136) );
ms00f80 configuration_wb_img_ctrl1_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(n_8477), .o(n_14907) );
ms00f80 configuration_wb_img_ctrl2_bit2_0_reg_0__u0 ( .ck(ispd_clk), .d(n_8460), .o(wbu_mrl_en_in_142) );
ms00f80 configuration_wb_img_ctrl2_bit2_0_reg_1__u0 ( .ck(ispd_clk), .d(n_8459), .o(wbu_pref_en_in_137) );
ms00f80 configuration_wb_img_ctrl2_bit2_0_reg_2__u0 ( .ck(ispd_clk), .d(n_8458), .o(n_14906) );
ms00f80 configuration_wb_init_complete_out_reg_u0 ( .ck(ispd_clk), .d(configuration_sync_init_complete), .o(wbu_wb_init_complete_in) );
ms00f80 configuration_wb_ta1_reg_31__u0 ( .ck(ispd_clk), .d(n_8520), .o(n_14909) );
ms00f80 configuration_wb_ta2_reg_31__u0 ( .ck(ispd_clk), .d(n_8516), .o(n_14908) );
na02f80 g10_u0 ( .a(wbs_cti_i_0_), .b(wbs_cti_i_2_), .o(n_16963) );
na02f10 g13_u0 ( .a(parchk_pci_cbe_reg_in_1238), .b(parchk_pci_cbe_reg_in_1236), .o(n_15958) );
in01f08 g14_u0 ( .a(n_15959), .o(n_15960) );
na02f10 g15_u0 ( .a(parchk_pci_cbe_reg_in_1237), .b(parchk_pci_cbe_reg_in), .o(g15_p) );
in01f10 g15_u1 ( .a(g15_p), .o(n_15959) );
in01f80 g16_u0 ( .a(parchk_pci_cbe_reg_in_1238), .o(n_1061) );
na02f20 g17_u0 ( .a(wishbone_slave_unit_pcim_sm_rdy_in), .b(n_15262), .o(g17_p) );
in01f10 g17_u1 ( .a(g17_p), .o(n_15054) );
na02s01 TIMEBOOST_cell_31089 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_9649) );
no02m10 g20_u0 ( .a(n_15999), .b(n_15998), .o(n_16001) );
in01f06 g21_u0 ( .a(n_16577), .o(n_16578) );
no02f20 g22_u0 ( .a(n_1323), .b(n_15371), .o(g22_p) );
in01f10 g22_u1 ( .a(g22_p), .o(n_15055) );
na02f10 g23_dup_u0 ( .a(n_16487), .b(n_16089), .o(n_16576) );
in01f20 g23_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_), .o(n_16071) );
no02f10 g25_u0 ( .a(FE_OCPN1852_n_16538), .b(n_15210), .o(n_15065) );
no02f10 g27_u0 ( .a(n_15924), .b(n_15998), .o(n_15231) );
na02f10 g28_dup74417_u0 ( .a(n_15746), .b(n_15924), .o(n_15748) );
no02f10 g28_dup_u0 ( .a(n_15403), .b(n_15397), .o(n_15512) );
ao22f06 g31_u0 ( .a(configuration_pci_err_data_510), .b(FE_OFN1063_n_15808), .c(n_16810), .d(n_14912), .o(n_15813) );
na03f02 TIMEBOOST_cell_66431 ( .a(TIMEBOOST_net_16782), .b(FE_OFN1315_n_6624), .c(g62906_sb), .o(n_6065) );
no02f40 g33_u0 ( .a(n_16460), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_16914) );
na02f20 g34_u0 ( .a(n_931), .b(n_370), .o(n_16021) );
na03f02 TIMEBOOST_cell_34885 ( .a(TIMEBOOST_net_9373), .b(FE_OFN1374_n_8567), .c(g57350_sb), .o(n_11399) );
na04f04 TIMEBOOST_cell_24236 ( .a(n_9045), .b(g57386_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q), .d(FE_OFN1406_n_8567), .o(n_10377) );
na02s01 TIMEBOOST_cell_45363 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q), .o(TIMEBOOST_net_13576) );
na02m02 TIMEBOOST_cell_54222 ( .a(TIMEBOOST_net_17328), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_15882) );
no02f40 g46_u0 ( .a(n_1177), .b(n_906), .o(n_16154) );
in01f20 g47_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_control_in_86), .o(n_16157) );
oa12m02 g52241_u0 ( .a(n_7740), .b(n_14888), .c(parity_checker_master_perr_report), .o(n_14901) );
na03f02 g52244_u0 ( .a(n_14900), .b(n_14306), .c(n_14902), .o(n_14904) );
na03f02 g52245_u0 ( .a(n_14899), .b(n_14304), .c(n_14902), .o(n_14903) );
ao12s01 g52246_u0 ( .a(parity_checker_pci_perr_en_reg), .b(parity_checker_perr_sampled), .c(n_13766), .o(n_14888) );
no02f02 g52252_u0 ( .a(n_14892), .b(n_14898), .o(g52252_p) );
in01f02 g52252_u1 ( .a(g52252_p), .o(n_14900) );
no02f02 g52253_u0 ( .a(n_14891), .b(n_14898), .o(g52253_p) );
in01f02 g52253_u1 ( .a(g52253_p), .o(n_14899) );
na03m06 TIMEBOOST_cell_72771 ( .a(n_4482), .b(FE_OFN640_n_4669), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q), .o(TIMEBOOST_net_23229) );
na04m06 TIMEBOOST_cell_73189 ( .a(FE_OFN1807_n_4501), .b(g64867_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q), .d(TIMEBOOST_net_14602), .o(TIMEBOOST_net_17507) );
in01s03 TIMEBOOST_cell_45904 ( .a(TIMEBOOST_net_13864), .o(TIMEBOOST_net_13865) );
na03f02 TIMEBOOST_cell_34789 ( .a(TIMEBOOST_net_9542), .b(FE_OFN1404_n_8567), .c(g57329_sb), .o(n_11420) );
ao12f02 g52353_u0 ( .a(n_14889), .b(n_14890), .c(wbm_cti_o_0_), .o(n_14892) );
ao12f02 g52354_u0 ( .a(n_14889), .b(n_14890), .c(wbm_cti_o_2_), .o(n_14891) );
oa12f02 g52390_u0 ( .a(n_14308), .b(n_14586), .c(n_9178), .o(n_14630) );
no02s01 g52391_u0 ( .a(n_14662), .b(parity_checker_check_perr), .o(n_14765) );
ao12f02 g52392_u0 ( .a(n_14806), .b(n_14764), .c(n_14967), .o(n_14889) );
in01f02 g52393_u0 ( .a(n_8757), .o(g52393_sb) );
na02f01 TIMEBOOST_cell_3640 ( .a(n_2367), .b(n_3498), .o(TIMEBOOST_net_380) );
in01m02 g52394_u0 ( .a(n_8757), .o(g52394_sb) );
na02s01 TIMEBOOST_cell_3618 ( .a(n_14079), .b(parchk_pci_serr_out_in), .o(TIMEBOOST_net_369) );
na02m02 TIMEBOOST_cell_62615 ( .a(TIMEBOOST_net_20254), .b(FE_OFN1011_n_4734), .o(TIMEBOOST_net_16926) );
in01f02 g52395_u0 ( .a(n_14839), .o(g52395_sb) );
na02f01 TIMEBOOST_cell_70346 ( .a(TIMEBOOST_net_17288), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_22381) );
na03f02 TIMEBOOST_cell_34883 ( .a(TIMEBOOST_net_9372), .b(FE_OFN1387_n_8567), .c(g57183_sb), .o(n_11571) );
na02f06 g54202_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_393), .b(g54202_sb), .o(g54202_da) );
in01f02 g52396_u0 ( .a(n_8757), .o(g52396_sb) );
na02f02 TIMEBOOST_cell_71637 ( .a(TIMEBOOST_net_23026), .b(FE_OFN1584_n_12306), .o(n_12764) );
na02s01 TIMEBOOST_cell_52373 ( .a(parchk_pci_ad_out_in_1195), .b(configuration_wb_err_data_598), .o(TIMEBOOST_net_16404) );
in01f02 g52397_u0 ( .a(n_14839), .o(g52397_sb) );
na02m04 TIMEBOOST_cell_53805 ( .a(n_4327), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q), .o(TIMEBOOST_net_17120) );
na03f02 TIMEBOOST_cell_66939 ( .a(FE_OFN1753_n_12086), .b(FE_OFN1568_n_11027), .c(TIMEBOOST_net_13613), .o(n_12664) );
in01f02 g52398_u0 ( .a(n_14839), .o(g52398_sb) );
na02f02 TIMEBOOST_cell_70751 ( .a(TIMEBOOST_net_22583), .b(n_1848), .o(n_3298) );
in01m02 g52399_u0 ( .a(n_8757), .o(g52399_sb) );
na02m10 TIMEBOOST_cell_3945 ( .a(TIMEBOOST_net_532), .b(n_1616), .o(n_1617) );
na02m04 g52399_u2 ( .a(n_14751), .b(n_8757), .o(g52399_db) );
in01m04 TIMEBOOST_cell_47506 ( .a(TIMEBOOST_net_13969), .o(TIMEBOOST_net_13968) );
in01m02 g52400_u0 ( .a(n_14839), .o(g52400_sb) );
na02m01 TIMEBOOST_cell_38238 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_10731) );
na03s06 TIMEBOOST_cell_68402 ( .a(TIMEBOOST_net_21187), .b(g65794_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_21409) );
in01f02 g52401_u0 ( .a(n_8757), .o(g52401_sb) );
na04f04 TIMEBOOST_cell_33806 ( .a(n_2203), .b(g61722_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q), .d(FE_OFN2081_n_8176), .o(n_8379) );
na04f02 TIMEBOOST_cell_36834 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q), .b(FE_OFN1394_n_8567), .c(n_9090), .d(g57203_sb), .o(n_10444) );
in01f02 g52402_u0 ( .a(n_14837), .o(g52402_sb) );
no02f01 TIMEBOOST_cell_3972 ( .a(wbu_pciif_frame_out_in), .b(wishbone_slave_unit_pci_initiator_sm_timeout), .o(TIMEBOOST_net_546) );
na02f01 g52402_u2 ( .a(n_14747), .b(n_14837), .o(g52402_db) );
na02f02 TIMEBOOST_cell_71727 ( .a(TIMEBOOST_net_23071), .b(FE_OCP_RBN1961_FE_OFN1591_n_13741), .o(n_14401) );
in01f02 g52403_u0 ( .a(n_8757), .o(g52403_sb) );
na04f04 TIMEBOOST_cell_24618 ( .a(n_9701), .b(g57137_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q), .d(FE_OFN2173_n_8567), .o(n_11613) );
na02m04 TIMEBOOST_cell_62426 ( .a(TIMEBOOST_net_10205), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q), .o(TIMEBOOST_net_20160) );
in01m02 g52404_u0 ( .a(n_14839), .o(g52404_sb) );
na02f01 TIMEBOOST_cell_3646 ( .a(n_4743), .b(n_2308), .o(TIMEBOOST_net_383) );
na03m02 TIMEBOOST_cell_72920 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(FE_OFN1042_n_2037), .c(TIMEBOOST_net_23232), .o(n_1881) );
in01f02 g52405_u0 ( .a(n_14839), .o(g52405_sb) );
na02m01 TIMEBOOST_cell_3974 ( .a(pciu_cache_lsize_not_zero_in), .b(n_16818), .o(TIMEBOOST_net_547) );
na03f02 TIMEBOOST_cell_64647 ( .a(TIMEBOOST_net_14136), .b(g64188_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q), .o(TIMEBOOST_net_17313) );
oa12m02 g52406_u0 ( .a(n_13398), .b(n_14802), .c(FE_OFN2163_n_16301), .o(n_14887) );
oa12m02 g52408_u0 ( .a(n_13395), .b(n_14799), .c(FE_OFN2165_n_16301), .o(n_14885) );
oa12m02 g52409_u0 ( .a(n_13394), .b(n_14798), .c(FE_OFN2165_n_16301), .o(n_14884) );
oa12m02 g52410_u0 ( .a(n_13393), .b(n_14797), .c(FE_OFN2165_n_16301), .o(n_14883) );
oa12m02 g52411_u0 ( .a(n_13392), .b(n_14796), .c(FE_OFN2165_n_16301), .o(n_14881) );
oa12m02 g52412_u0 ( .a(n_13391), .b(n_14763), .c(n_16305), .o(n_14851) );
oa12m02 g52413_u0 ( .a(n_13389), .b(n_14793), .c(FE_OFN2165_n_16301), .o(n_14880) );
oa12m02 g52414_u0 ( .a(n_13390), .b(n_14794), .c(FE_OFN2165_n_16301), .o(n_14879) );
oa12m02 g52415_u0 ( .a(n_13388), .b(n_14762), .c(FE_OFN2165_n_16301), .o(n_14850) );
oa12m02 g52416_u0 ( .a(n_13387), .b(n_14792), .c(FE_OFN2165_n_16301), .o(n_14877) );
oa12f02 g52417_u0 ( .a(n_13386), .b(n_14791), .c(FE_OFN2163_n_16301), .o(n_14875) );
oa12m02 g52418_u0 ( .a(n_13384), .b(n_14790), .c(FE_OFN2165_n_16301), .o(n_14873) );
oa12m02 g52419_u0 ( .a(n_13383), .b(n_14789), .c(FE_OFN2165_n_16301), .o(n_14871) );
oa12m02 g52421_u0 ( .a(n_13381), .b(n_14786), .c(FE_OFN2165_n_16301), .o(n_14869) );
oa12m02 g52422_u0 ( .a(n_13380), .b(n_14784), .c(FE_OFN2162_n_16301), .o(n_14867) );
oa12m02 g52423_u0 ( .a(n_13379), .b(n_14783), .c(FE_OFN2162_n_16301), .o(n_14866) );
oa12m02 g52424_u0 ( .a(n_13378), .b(n_14781), .c(FE_OFN2164_n_16301), .o(n_14865) );
oa12m02 g52425_u0 ( .a(n_13376), .b(n_14778), .c(FE_OFN2162_n_16301), .o(n_14864) );
oa12m02 g52426_u0 ( .a(n_13377), .b(n_14780), .c(FE_OFN2164_n_16301), .o(n_14863) );
oa12m02 g52427_u0 ( .a(n_13375), .b(n_14777), .c(FE_OFN2162_n_16301), .o(n_14862) );
oa12f02 g52428_u0 ( .a(n_13374), .b(n_14776), .c(FE_OFN2162_n_16301), .o(n_14861) );
oa12m02 g52429_u0 ( .a(n_13373), .b(n_14775), .c(FE_OFN2162_n_16301), .o(n_14860) );
oa12m02 g52430_u0 ( .a(n_13371), .b(n_14772), .c(FE_OFN2163_n_16301), .o(n_14859) );
oa12m02 g52431_u0 ( .a(n_13370), .b(n_14770), .c(n_16305), .o(n_14858) );
oa12m02 g52432_u0 ( .a(n_13372), .b(n_14773), .c(n_16305), .o(n_14856) );
oa12m02 g52433_u0 ( .a(n_13369), .b(n_14769), .c(n_16305), .o(n_14855) );
oa12f02 g52434_u0 ( .a(n_13368), .b(n_14768), .c(FE_OFN2163_n_16301), .o(n_14854) );
oa12f02 g52435_u0 ( .a(n_13367), .b(n_14761), .c(FE_OFN2164_n_16301), .o(n_14849) );
oa12m02 g52436_u0 ( .a(n_13366), .b(n_14767), .c(FE_OFN2164_n_16301), .o(n_14853) );
oa12m02 g52437_u0 ( .a(n_13365), .b(n_14766), .c(FE_OFN2164_n_16301), .o(n_14852) );
na02m10 TIMEBOOST_cell_52949 ( .a(wishbone_slave_unit_pcim_sm_data_in_646), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q), .o(TIMEBOOST_net_16692) );
na02f02 g52439_u2 ( .a(n_14682), .b(n_14837), .o(g52439_db) );
in01s01 TIMEBOOST_cell_73909 ( .a(TIMEBOOST_net_23473), .o(TIMEBOOST_net_23474) );
in01f02 g52440_u0 ( .a(n_14839), .o(g52440_sb) );
na04f04 TIMEBOOST_cell_67485 ( .a(TIMEBOOST_net_14570), .b(g65909_sb), .c(TIMEBOOST_net_20381), .d(g62016_sb), .o(n_7863) );
na03s02 TIMEBOOST_cell_70470 ( .a(FE_OFN592_n_9694), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q), .c(FE_OFN219_n_9853), .o(TIMEBOOST_net_22443) );
in01f02 g52441_u0 ( .a(n_14839), .o(g52441_sb) );
na02s01 TIMEBOOST_cell_39765 ( .a(TIMEBOOST_net_11494), .b(g57973_db), .o(n_9115) );
na02f02 g54200_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_391), .b(g54200_sb), .o(g54200_da) );
in01f02 g52442_u0 ( .a(n_8757), .o(g52442_sb) );
na03m04 TIMEBOOST_cell_73002 ( .a(TIMEBOOST_net_22001), .b(FE_OFN1051_n_16657), .c(TIMEBOOST_net_23259), .o(TIMEBOOST_net_21063) );
in01f02 TIMEBOOST_cell_47508 ( .a(TIMEBOOST_net_13971), .o(TIMEBOOST_net_13970) );
in01f02 g52443_u0 ( .a(n_8757), .o(g52443_sb) );
na04f04 TIMEBOOST_cell_24588 ( .a(n_9777), .b(g57146_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q), .d(FE_OFN2182_n_8567), .o(n_11604) );
na03f08 TIMEBOOST_cell_72401 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_397), .b(n_13447), .c(n_13781), .o(TIMEBOOST_net_22055) );
na04f40 TIMEBOOST_cell_67135 ( .a(FE_OFN2055_n_8831), .b(g58774_sb), .c(wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q), .d(wbu_addr_in_271), .o(n_9122) );
in01f02 g52444_u0 ( .a(n_14839), .o(g52444_sb) );
na02s01 TIMEBOOST_cell_38307 ( .a(TIMEBOOST_net_10765), .b(g52479_sb), .o(TIMEBOOST_net_712) );
na04f04 TIMEBOOST_cell_36836 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q), .b(FE_OFN1414_n_8567), .c(n_9763), .d(g57158_sb), .o(n_11592) );
na04f04 TIMEBOOST_cell_36106 ( .a(parchk_pci_ad_out_in_1182), .b(g62085_sb), .c(configuration_wb_err_data_585), .d(FE_OFN1173_n_5592), .o(n_5623) );
na02f02 g52445_u2 ( .a(n_14678), .b(n_14837), .o(g52445_db) );
na02s01 TIMEBOOST_cell_43013 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q), .b(FE_OFN585_n_9692), .o(TIMEBOOST_net_12401) );
in01f01 g52446_u0 ( .a(n_8757), .o(g52446_sb) );
in01s01 TIMEBOOST_cell_45994 ( .a(TIMEBOOST_net_13954), .o(TIMEBOOST_net_13955) );
na02s02 TIMEBOOST_cell_63892 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q), .o(TIMEBOOST_net_20932) );
na02f02 TIMEBOOST_cell_39483 ( .a(TIMEBOOST_net_11353), .b(g59373_sb), .o(n_7687) );
in01m02 g52447_u0 ( .a(n_14839), .o(g52447_sb) );
na02f02 g52447_u2 ( .a(n_14750), .b(n_14839), .o(g52447_db) );
in01f02 g52448_u0 ( .a(n_14839), .o(g52448_sb) );
na02f02 TIMEBOOST_cell_3249 ( .a(TIMEBOOST_net_184), .b(n_3313), .o(n_3436) );
na02m02 TIMEBOOST_cell_68973 ( .a(TIMEBOOST_net_21694), .b(g64153_sb), .o(TIMEBOOST_net_8800) );
na04f02 TIMEBOOST_cell_25259 ( .a(n_16616), .b(n_13923), .c(n_16617), .d(n_13846), .o(n_14577) );
in01f02 g52449_u0 ( .a(n_14839), .o(g52449_sb) );
na03m04 TIMEBOOST_cell_72724 ( .a(g64361_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q), .c(TIMEBOOST_net_14286), .o(TIMEBOOST_net_17317) );
na03m02 TIMEBOOST_cell_72723 ( .a(g64348_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q), .c(TIMEBOOST_net_21992), .o(TIMEBOOST_net_13063) );
na02f02 TIMEBOOST_cell_39607 ( .a(TIMEBOOST_net_11415), .b(g63118_sb), .o(n_5021) );
in01f02 g52450_u0 ( .a(n_14839), .o(g52450_sb) );
na02s02 TIMEBOOST_cell_28190 ( .a(TIMEBOOST_net_8199), .b(g65774_sb), .o(n_2193) );
na03f02 TIMEBOOST_cell_34889 ( .a(TIMEBOOST_net_9377), .b(FE_OFN1391_n_8567), .c(g57185_sb), .o(n_11568) );
in01f02 g52451_u0 ( .a(n_14839), .o(g52451_sb) );
na02m20 TIMEBOOST_cell_3448 ( .a(n_2316), .b(n_2308), .o(TIMEBOOST_net_284) );
na03f02 TIMEBOOST_cell_34905 ( .a(TIMEBOOST_net_9484), .b(FE_OFN1368_n_8567), .c(g57161_sb), .o(n_10460) );
in01f02 g52452_u0 ( .a(n_14839), .o(g52452_sb) );
na03s01 TIMEBOOST_cell_72453 ( .a(n_2512), .b(FE_OFN2094_n_2520), .c(g66419_db), .o(n_2513) );
na02s01 TIMEBOOST_cell_39769 ( .a(TIMEBOOST_net_11496), .b(g58034_db), .o(n_9097) );
na02m03 TIMEBOOST_cell_3644 ( .a(n_4743), .b(n_2742), .o(TIMEBOOST_net_382) );
na03m02 TIMEBOOST_cell_72371 ( .a(configuration_sync_command_bit2), .b(wbu_wb_init_complete_in), .c(wishbone_slave_unit_wishbone_slave_img_wallow), .o(TIMEBOOST_net_16412) );
in01f02 g52454_u0 ( .a(n_14839), .o(g52454_sb) );
na02s01 TIMEBOOST_cell_45365 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q), .o(TIMEBOOST_net_13577) );
na03f02 TIMEBOOST_cell_34887 ( .a(TIMEBOOST_net_9340), .b(FE_OFN1390_n_8567), .c(g57418_sb), .o(n_11322) );
na03f02 TIMEBOOST_cell_67934 ( .a(n_3917), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q), .c(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_15179) );
in01f02 g52455_u0 ( .a(n_8757), .o(g52455_sb) );
na02m02 TIMEBOOST_cell_70865 ( .a(TIMEBOOST_net_22640), .b(g58196_sb), .o(n_9590) );
in01s01 g52456_u0 ( .a(FE_OFN1021_n_11877), .o(g52456_sb) );
na02s01 g52456_u1 ( .a(wbs_adr_i_10_), .b(g52456_sb), .o(g52456_da) );
in01m08 g52457_u0 ( .a(FE_OFN1022_n_11877), .o(g52457_sb) );
na02s01 TIMEBOOST_cell_53437 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q), .o(TIMEBOOST_net_16936) );
na03s02 TIMEBOOST_cell_73334 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q), .c(TIMEBOOST_net_20506), .o(TIMEBOOST_net_16427) );
in01f04 g52458_u0 ( .a(FE_OFN1022_n_11877), .o(g52458_sb) );
na02f02 TIMEBOOST_cell_50362 ( .a(TIMEBOOST_net_15398), .b(g62336_sb), .o(n_6926) );
na02m01 TIMEBOOST_cell_42781 ( .a(pci_ad_i_5_), .b(parchk_pci_ad_reg_in_1209), .o(TIMEBOOST_net_12285) );
na04s02 TIMEBOOST_cell_73081 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q), .b(g65841_sb), .c(TIMEBOOST_net_23392), .d(FE_OFN1042_n_2037), .o(n_1879) );
in01f02 g52459_u0 ( .a(FE_OFN1022_n_11877), .o(g52459_sb) );
na02s01 g52459_u1 ( .a(wbs_adr_i_13_), .b(g52459_sb), .o(g52459_da) );
na03m04 TIMEBOOST_cell_72856 ( .a(n_3785), .b(FE_OFN642_n_4677), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q), .o(TIMEBOOST_net_23256) );
na03f02 TIMEBOOST_cell_72373 ( .a(TIMEBOOST_net_21228), .b(pci_target_unit_del_sync_comp_cycle_count_0_), .c(n_1187), .o(n_1425) );
in01m02 g52460_u0 ( .a(FE_OFN1021_n_11877), .o(g52460_sb) );
na02m01 TIMEBOOST_cell_53438 ( .a(TIMEBOOST_net_16936), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_14736) );
na02m02 TIMEBOOST_cell_49721 ( .a(g58384_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q), .o(TIMEBOOST_net_15078) );
in01m04 g52461_u0 ( .a(FE_OFN1022_n_11877), .o(g52461_sb) );
in01s01 TIMEBOOST_cell_67748 ( .a(TIMEBOOST_net_21174), .o(TIMEBOOST_net_21175) );
na04f04 TIMEBOOST_cell_34714 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q), .b(FE_OFN1349_n_8567), .c(n_9713), .d(g57222_sb), .o(n_11533) );
in01f01 g52462_u0 ( .a(FE_OFN1022_n_11877), .o(g52462_sb) );
na02s01 g52462_u1 ( .a(wbs_adr_i_16_), .b(g52462_sb), .o(g52462_da) );
na02m02 TIMEBOOST_cell_62614 ( .a(TIMEBOOST_net_12407), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q), .o(TIMEBOOST_net_20254) );
na02f02 TIMEBOOST_cell_49954 ( .a(TIMEBOOST_net_15194), .b(g63087_sb), .o(n_5080) );
in01f04 g52463_u0 ( .a(FE_OFN1022_n_11877), .o(g52463_sb) );
no03f04 TIMEBOOST_cell_34717 ( .a(FE_RN_565_0), .b(n_7552), .c(FE_RN_569_0), .o(TIMEBOOST_net_463) );
in01s01 g52464_u0 ( .a(FE_OFN1021_n_11877), .o(g52464_sb) );
na02s01 g52464_u1 ( .a(wbs_adr_i_18_), .b(g52464_sb), .o(g52464_da) );
na02f02 TIMEBOOST_cell_40847 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_12035), .o(n_12527) );
na02m10 TIMEBOOST_cell_72348 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q), .o(TIMEBOOST_net_23382) );
na04f02 TIMEBOOST_cell_35123 ( .a(wbs_dat_o_0_), .b(g52504_sb), .c(wbs_wbb3_2_wbb2_dat_o_i), .d(FE_OFN1471_g52675_p), .o(n_13727) );
na03f02 TIMEBOOST_cell_34966 ( .a(TIMEBOOST_net_9476), .b(FE_OFN1374_n_8567), .c(g57590_sb), .o(n_10289) );
in01f01 g52466_u0 ( .a(FE_OFN1021_n_11877), .o(g52466_sb) );
na02s01 g52466_u1 ( .a(wbs_adr_i_20_), .b(g52466_sb), .o(g52466_da) );
na03f02 TIMEBOOST_cell_34987 ( .a(TIMEBOOST_net_9516), .b(FE_OFN1401_n_8567), .c(g57302_sb), .o(n_10407) );
na03f02 TIMEBOOST_cell_34968 ( .a(TIMEBOOST_net_9537), .b(FE_OFN1414_n_8567), .c(g57427_sb), .o(n_11307) );
na02m10 TIMEBOOST_cell_69406 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q), .o(TIMEBOOST_net_21911) );
na03m02 TIMEBOOST_cell_73082 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q), .b(g58298_sb), .c(TIMEBOOST_net_11146), .o(TIMEBOOST_net_9488) );
na02s01 g52468_u1 ( .a(wbs_adr_i_22_), .b(g52463_sb), .o(g52468_da) );
na03f02 TIMEBOOST_cell_34959 ( .a(TIMEBOOST_net_9561), .b(FE_OFN1391_n_8567), .c(g57407_sb), .o(n_10366) );
na02m06 TIMEBOOST_cell_70242 ( .a(TIMEBOOST_net_9986), .b(FE_OFN881_g64577_p), .o(TIMEBOOST_net_22329) );
na02m02 TIMEBOOST_cell_69386 ( .a(g64958_sb), .b(n_119), .o(TIMEBOOST_net_21901) );
na02m02 TIMEBOOST_cell_53414 ( .a(TIMEBOOST_net_16924), .b(g58332_sb), .o(n_9022) );
in01m08 g52470_u0 ( .a(FE_OFN1023_n_11877), .o(g52470_sb) );
na04m06 TIMEBOOST_cell_72774 ( .a(n_4452), .b(g64901_sb), .c(n_4410), .d(g64901_db), .o(TIMEBOOST_net_13360) );
na03f02 TIMEBOOST_cell_34967 ( .a(TIMEBOOST_net_9477), .b(FE_OFN1368_n_8567), .c(g57126_sb), .o(n_10474) );
na03f02 TIMEBOOST_cell_34970 ( .a(TIMEBOOST_net_9460), .b(FE_OFN1382_n_8567), .c(g57476_sb), .o(n_10336) );
na02m02 TIMEBOOST_cell_51000 ( .a(TIMEBOOST_net_15717), .b(g62383_sb), .o(n_6835) );
na03m04 TIMEBOOST_cell_73190 ( .a(g64760_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q), .c(TIMEBOOST_net_16378), .o(TIMEBOOST_net_17369) );
na02s01 g52472_u1 ( .a(wbs_adr_i_26_), .b(g52458_sb), .o(g52472_da) );
na03f02 TIMEBOOST_cell_34781 ( .a(TIMEBOOST_net_9420), .b(FE_OFN1404_n_8567), .c(g57105_sb), .o(n_11640) );
na02s01 TIMEBOOST_cell_44445 ( .a(g58377_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q), .o(TIMEBOOST_net_13117) );
na02m02 TIMEBOOST_cell_49722 ( .a(TIMEBOOST_net_15078), .b(TIMEBOOST_net_11197), .o(TIMEBOOST_net_9360) );
na02s02 TIMEBOOST_cell_49723 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q), .b(FE_OFN539_n_9690), .o(TIMEBOOST_net_15079) );
na02s01 TIMEBOOST_cell_42737 ( .a(wbu_addr_in_254), .b(n_8831), .o(TIMEBOOST_net_12263) );
na02m04 TIMEBOOST_cell_69824 ( .a(g64832_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q), .o(TIMEBOOST_net_22120) );
na03m02 TIMEBOOST_cell_70108 ( .a(g65828_db), .b(TIMEBOOST_net_12760), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q), .o(TIMEBOOST_net_22262) );
na02f02 TIMEBOOST_cell_45430 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13609), .o(TIMEBOOST_net_12041) );
in01s01 g52476_u0 ( .a(FE_OFN1021_n_11877), .o(g52476_sb) );
na02s01 g52476_u1 ( .a(wbs_adr_i_30_), .b(g52476_sb), .o(g52476_da) );
na03f02 TIMEBOOST_cell_67038 ( .a(FE_OFN1606_n_13997), .b(TIMEBOOST_net_13754), .c(FE_OFN1599_n_13995), .o(n_14469) );
no03f06 TIMEBOOST_cell_66820 ( .a(TIMEBOOST_net_20659), .b(TIMEBOOST_net_771), .c(n_7823), .o(g53078_p) );
in01m04 g52477_u0 ( .a(FE_OFN1025_n_11877), .o(g52477_sb) );
na02m01 g52477_u1 ( .a(wbs_adr_i_29_), .b(g52477_sb), .o(g52477_da) );
na03f02 TIMEBOOST_cell_34972 ( .a(TIMEBOOST_net_9478), .b(FE_OFN1377_n_8567), .c(g57131_sb), .o(n_10473) );
na02m10 TIMEBOOST_cell_50013 ( .a(wishbone_slave_unit_pcim_sm_data_in_663), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q), .o(TIMEBOOST_net_15224) );
in01m02 g52478_u0 ( .a(FE_OFN8_n_11877), .o(g52478_sb) );
na02m01 g52478_u1 ( .a(wbs_adr_i_31_), .b(g52478_sb), .o(g52478_da) );
in01f01 g52479_u0 ( .a(FE_OFN1024_n_11877), .o(g52479_sb) );
na02s01 g52479_u1 ( .a(wbs_adr_i_3_), .b(g52479_sb), .o(g52479_da) );
na03m02 TIMEBOOST_cell_64646 ( .a(TIMEBOOST_net_12342), .b(n_3744), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q), .o(TIMEBOOST_net_17062) );
na04s02 TIMEBOOST_cell_72955 ( .a(TIMEBOOST_net_10712), .b(g65748_sb), .c(g61798_sb), .d(g61798_db), .o(n_8200) );
na02f02 TIMEBOOST_cell_71059 ( .a(TIMEBOOST_net_22737), .b(g63151_sb), .o(n_5838) );
na02f01 TIMEBOOST_cell_62613 ( .a(TIMEBOOST_net_20253), .b(FE_OFN908_n_4734), .o(TIMEBOOST_net_16254) );
na02s01 TIMEBOOST_cell_45431 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q), .o(TIMEBOOST_net_13610) );
in01s01 g52482_u0 ( .a(FE_OFN8_n_11877), .o(g52482_sb) );
na02s02 g52482_u1 ( .a(wbs_adr_i_6_), .b(g52482_sb), .o(g52482_da) );
na03f02 TIMEBOOST_cell_34985 ( .a(TIMEBOOST_net_9388), .b(FE_OFN1380_n_8567), .c(g57121_sb), .o(n_10476) );
na03f02 TIMEBOOST_cell_34974 ( .a(TIMEBOOST_net_9565), .b(FE_OFN1388_n_8567), .c(g57490_sb), .o(n_11246) );
na03f02 TIMEBOOST_cell_34965 ( .a(TIMEBOOST_net_9436), .b(FE_OFN1388_n_8567), .c(g57317_sb), .o(n_11434) );
na03f02 TIMEBOOST_cell_34976 ( .a(TIMEBOOST_net_9438), .b(FE_OFN1413_n_8567), .c(g57497_sb), .o(n_10329) );
na03f02 TIMEBOOST_cell_66684 ( .a(TIMEBOOST_net_17562), .b(FE_OFN1270_n_4095), .c(g62510_sb), .o(n_6558) );
na03f02 TIMEBOOST_cell_34971 ( .a(TIMEBOOST_net_9483), .b(FE_OFN1401_n_8567), .c(g57503_sb), .o(n_11235) );
na04f04 TIMEBOOST_cell_67930 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q), .b(FE_OFN2212_n_8407), .c(n_2177), .d(g62017_sb), .o(n_7861) );
na02f02 TIMEBOOST_cell_50422 ( .a(TIMEBOOST_net_15428), .b(g62621_sb), .o(n_6315) );
na02m08 TIMEBOOST_cell_52863 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q), .b(wbs_dat_i_13_), .o(TIMEBOOST_net_16649) );
na02f02 TIMEBOOST_cell_71199 ( .a(TIMEBOOST_net_22807), .b(g62403_sb), .o(n_6793) );
no02f02 g52495_u0 ( .a(n_14760), .b(FE_OFN2163_n_16301), .o(g52495_p) );
in01f02 g52495_u1 ( .a(g52495_p), .o(n_14833) );
no02f02 g52496_u0 ( .a(n_14759), .b(FE_OFN2163_n_16301), .o(g52496_p) );
in01f02 g52496_u1 ( .a(g52496_p), .o(n_14832) );
no02f02 g52497_u0 ( .a(n_14757), .b(FE_OFN2163_n_16301), .o(g52497_p) );
in01f02 g52497_u1 ( .a(g52497_p), .o(n_14830) );
no02f02 g52498_u0 ( .a(n_14756), .b(FE_OFN2163_n_16301), .o(g52498_p) );
in01f02 g52498_u1 ( .a(g52498_p), .o(n_14829) );
oa12f01 g52499_u0 ( .a(n_10793), .b(FE_OFN3_n_4778), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(n_11844) );
na02f02 g52500_u0 ( .a(n_8880), .b(n_14691), .o(n_14804) );
na02f02 g52501_u0 ( .a(n_8879), .b(n_14690), .o(n_14805) );
ao12s01 g52502_u0 ( .a(n_14624), .b(parchk_pci_perr_out_in), .c(out_bckp_perr_en_out), .o(n_14662) );
in01f02 g52503_u0 ( .a(FE_OFN2243_g52675_p), .o(g52503_sb) );
na04f04 TIMEBOOST_cell_24661 ( .a(n_9094), .b(g57179_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q), .d(FE_OFN2180_n_8567), .o(n_10450) );
na03f02 TIMEBOOST_cell_34969 ( .a(TIMEBOOST_net_9437), .b(FE_OFN1414_n_8567), .c(g57499_sb), .o(n_11239) );
na04f02 TIMEBOOST_cell_73691 ( .a(wishbone_slave_unit_wishbone_slave_del_completion_allow), .b(n_7115), .c(FE_OFN1189_n_5742), .d(g59350_sb), .o(n_7701) );
in01f02 g52504_u0 ( .a(FE_OFN1471_g52675_p), .o(g52504_sb) );
na04f04 TIMEBOOST_cell_24655 ( .a(n_9714), .b(g57221_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q), .d(FE_OFN2177_n_8567), .o(n_11534) );
na02s02 TIMEBOOST_cell_52892 ( .a(TIMEBOOST_net_16663), .b(TIMEBOOST_net_10825), .o(TIMEBOOST_net_9459) );
na03s02 TIMEBOOST_cell_72560 ( .a(pci_target_unit_del_sync_addr_in_216), .b(g66403_sb), .c(g66405_db), .o(n_2534) );
in01f02 g52505_u0 ( .a(FE_OFN2243_g52675_p), .o(g52505_sb) );
na02s02 TIMEBOOST_cell_37251 ( .a(TIMEBOOST_net_10237), .b(g65718_sb), .o(n_2197) );
na03f02 TIMEBOOST_cell_34953 ( .a(TIMEBOOST_net_9500), .b(FE_OFN1412_n_8567), .c(g57196_sb), .o(n_10446) );
na03f02 TIMEBOOST_cell_34978 ( .a(TIMEBOOST_net_9385), .b(FE_OFN1404_n_8567), .c(g57429_sb), .o(n_11305) );
in01f02 g52506_u0 ( .a(FE_OFN1471_g52675_p), .o(g52506_sb) );
na02f01 TIMEBOOST_cell_37034 ( .a(pci_target_unit_pci_target_sm_wr_to_fifo), .b(n_565), .o(TIMEBOOST_net_10129) );
in01s01 TIMEBOOST_cell_45882 ( .a(TIMEBOOST_net_13842), .o(TIMEBOOST_net_13843) );
na02m02 TIMEBOOST_cell_26309 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q), .b(g65352_sb), .o(TIMEBOOST_net_7259) );
in01f02 g52507_u0 ( .a(FE_OFN2243_g52675_p), .o(g52507_sb) );
na03f10 TIMEBOOST_cell_41271 ( .a(n_15680), .b(n_16871), .c(n_16860), .o(n_1805) );
na04f02 TIMEBOOST_cell_67660 ( .a(TIMEBOOST_net_20594), .b(g59234_sb), .c(TIMEBOOST_net_12861), .d(FE_OFN1145_n_15261), .o(n_13508) );
in01f02 g52508_u0 ( .a(FE_OFN2242_g52675_p), .o(g52508_sb) );
na02s01 TIMEBOOST_cell_47510 ( .a(TIMEBOOST_net_13972), .b(g67042_sb), .o(n_1431) );
na03f02 TIMEBOOST_cell_34979 ( .a(TIMEBOOST_net_9417), .b(FE_OFN1383_n_8567), .c(g57052_sb), .o(n_11684) );
na03f02 TIMEBOOST_cell_66227 ( .a(TIMEBOOST_net_20543), .b(FE_OFN1294_n_4098), .c(g62463_sb), .o(n_6670) );
in01f01 g52509_u0 ( .a(FE_OFN1472_g52675_p), .o(g52509_sb) );
na02f01 TIMEBOOST_cell_37035 ( .a(TIMEBOOST_net_10129), .b(n_5755), .o(FE_RN_268_0) );
na02s01 TIMEBOOST_cell_45429 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q), .o(TIMEBOOST_net_13609) );
na03f02 TIMEBOOST_cell_35142 ( .a(TIMEBOOST_net_8596), .b(n_13621), .c(g54337_sb), .o(n_13482) );
in01f02 g52510_u0 ( .a(FE_OFN2243_g52675_p), .o(g52510_sb) );
na04f04 TIMEBOOST_cell_24609 ( .a(n_9208), .b(g57542_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q), .d(FE_OFN2175_n_8567), .o(n_10812) );
na02m02 TIMEBOOST_cell_52320 ( .a(TIMEBOOST_net_16377), .b(TIMEBOOST_net_8311), .o(n_9509) );
na02m08 TIMEBOOST_cell_45281 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q), .o(TIMEBOOST_net_13535) );
in01f02 g52511_u0 ( .a(FE_OFN2243_g52675_p), .o(g52511_sb) );
na04f04 TIMEBOOST_cell_24611 ( .a(n_9436), .b(g57540_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q), .d(FE_OFN2167_n_8567), .o(n_11202) );
in01s01 TIMEBOOST_cell_45905 ( .a(TIMEBOOST_net_13866), .o(wbs_dat_i_17_) );
in01f02 g52512_u0 ( .a(FE_OFN2243_g52675_p), .o(g52512_sb) );
na04f04 TIMEBOOST_cell_24613 ( .a(n_9441), .b(g57532_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q), .d(FE_OFN2187_n_8567), .o(n_11209) );
in01s01 TIMEBOOST_cell_45906 ( .a(TIMEBOOST_net_13867), .o(TIMEBOOST_net_13866) );
na02f01 TIMEBOOST_cell_26115 ( .a(pci_target_unit_pcit_if_strd_addr_in_712), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7162) );
in01f02 g52513_u0 ( .a(FE_OFN2243_g52675_p), .o(g52513_sb) );
na04f04 TIMEBOOST_cell_24615 ( .a(n_9450), .b(g57522_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q), .d(FE_OFN2168_n_8567), .o(n_11219) );
na02f02 TIMEBOOST_cell_18713 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_do_del_request), .o(TIMEBOOST_net_5720) );
in01f02 g52514_u0 ( .a(FE_OFN2243_g52675_p), .o(g52514_sb) );
na04f04 TIMEBOOST_cell_24617 ( .a(n_9102), .b(g57144_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q), .d(FE_OFN2167_n_8567), .o(n_10464) );
na02s01 TIMEBOOST_cell_42815 ( .a(TIMEBOOST_net_10131), .b(n_574), .o(TIMEBOOST_net_12302) );
in01f01 g52515_u0 ( .a(FE_OFN1472_g52675_p), .o(g52515_sb) );
na04f04 TIMEBOOST_cell_24693 ( .a(wishbone_slave_unit_fifos_wbr_be_in_265), .b(g58840_sb), .c(TIMEBOOST_net_13855), .d(FE_OFN1438_n_9372), .o(n_8674) );
in01f02 g52516_u0 ( .a(FE_OFN2243_g52675_p), .o(g52516_sb) );
na04f04 TIMEBOOST_cell_24629 ( .a(n_9869), .b(g57067_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q), .d(FE_OFN2175_n_8567), .o(n_11675) );
na02s01 TIMEBOOST_cell_43573 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_121), .o(TIMEBOOST_net_12681) );
na02s01 TIMEBOOST_cell_43567 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_12678) );
in01f01 g52517_u0 ( .a(FE_OFN1472_g52675_p), .o(g52517_sb) );
na04f04 TIMEBOOST_cell_24695 ( .a(wishbone_slave_unit_fifos_wbr_be_in), .b(g58838_sb), .c(TIMEBOOST_net_13859), .d(FE_OFN1438_n_9372), .o(n_8676) );
in01s01 TIMEBOOST_cell_45883 ( .a(conf_wb_err_bc_in_848), .o(TIMEBOOST_net_13844) );
na02s01 TIMEBOOST_cell_43651 ( .a(pci_target_unit_del_sync_addr_in_229), .b(parchk_pci_ad_reg_in_1230), .o(TIMEBOOST_net_12720) );
in01f02 g52518_u0 ( .a(FE_OFN2241_g52675_p), .o(g52518_sb) );
na04f04 TIMEBOOST_cell_24627 ( .a(n_9855), .b(g57076_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q), .d(FE_OFN2182_n_8567), .o(n_11667) );
in01f02 g52519_u0 ( .a(FE_OFN1471_g52675_p), .o(g52519_sb) );
na03f02 TIMEBOOST_cell_73191 ( .a(TIMEBOOST_net_22222), .b(g61884_sb), .c(TIMEBOOST_net_22354), .o(n_8062) );
na02m04 TIMEBOOST_cell_43569 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_136), .o(TIMEBOOST_net_12679) );
na02m01 TIMEBOOST_cell_62612 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_144), .o(TIMEBOOST_net_20253) );
in01f02 g52520_u0 ( .a(FE_OFN2242_g52675_p), .o(g52520_sb) );
na04f04 TIMEBOOST_cell_24631 ( .a(n_9879), .b(g57050_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q), .d(FE_OFN2189_n_8567), .o(n_11685) );
na03m02 TIMEBOOST_cell_72966 ( .a(TIMEBOOST_net_23212), .b(g65423_sb), .c(TIMEBOOST_net_22020), .o(TIMEBOOST_net_17123) );
na02m02 TIMEBOOST_cell_64046 ( .a(TIMEBOOST_net_7595), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_21009) );
in01f02 g52521_u0 ( .a(FE_OFN2242_g52675_p), .o(g52521_sb) );
na04f04 TIMEBOOST_cell_24633 ( .a(n_9883), .b(g57046_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q), .d(FE_OFN2177_n_8567), .o(n_11688) );
na02f02 g60682_u1 ( .a(wbu_latency_tim_val_in_246), .b(g60682_sb), .o(g60682_da) );
in01f02 g52522_u0 ( .a(FE_OFN2243_g52675_p), .o(g52522_sb) );
na04f04 TIMEBOOST_cell_24635 ( .a(n_9134), .b(g57039_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q), .d(FE_OFN2168_n_8567), .o(n_10513) );
na02f01 TIMEBOOST_cell_52273 ( .a(TIMEBOOST_net_12712), .b(FE_OFN1051_n_16657), .o(TIMEBOOST_net_16354) );
in01f02 g52523_u0 ( .a(FE_OFN2241_g52675_p), .o(g52523_sb) );
na04f04 TIMEBOOST_cell_24637 ( .a(n_9648), .b(g57284_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q), .d(FE_OFN2188_n_8567), .o(n_11470) );
na03m08 TIMEBOOST_cell_69736 ( .a(g65394_sb), .b(FE_OFN1677_n_4655), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q), .o(TIMEBOOST_net_22076) );
in01f02 g52524_u0 ( .a(FE_OFN2242_g52675_p), .o(g52524_sb) );
na04f04 TIMEBOOST_cell_24639 ( .a(n_9069), .b(g57281_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q), .d(FE_OFN2169_n_8567), .o(n_10412) );
na02f02 TIMEBOOST_cell_50900 ( .a(TIMEBOOST_net_15667), .b(g62642_sb), .o(n_6264) );
in01f01 g52525_u0 ( .a(FE_OFN1472_g52675_p), .o(g52525_sb) );
na04m02 TIMEBOOST_cell_72972 ( .a(n_4452), .b(g64983_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q), .d(g64983_db), .o(TIMEBOOST_net_13371) );
na02f02 TIMEBOOST_cell_70246 ( .a(TIMEBOOST_net_14834), .b(FE_OFN1094_g64577_p), .o(TIMEBOOST_net_22331) );
na02s01 TIMEBOOST_cell_25283 ( .a(pci_ad_i_28_), .b(parchk_pci_ad_reg_in_1232), .o(TIMEBOOST_net_6746) );
in01f02 g52526_u0 ( .a(FE_OFN2243_g52675_p), .o(g52526_sb) );
na04f04 TIMEBOOST_cell_24641 ( .a(n_9663), .b(g57268_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q), .d(FE_OFN2170_n_8567), .o(n_11484) );
na03m02 TIMEBOOST_cell_65888 ( .a(n_3993), .b(g62858_sb), .c(g62858_db), .o(n_5251) );
in01f02 g52527_u0 ( .a(FE_OFN2243_g52675_p), .o(g52527_sb) );
na04f04 TIMEBOOST_cell_24643 ( .a(n_9076), .b(g57258_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q), .d(FE_OFN2179_n_8567), .o(n_10421) );
na02s01 TIMEBOOST_cell_25282 ( .a(TIMEBOOST_net_6745), .b(n_574), .o(TIMEBOOST_net_536) );
in01f01 g52528_u0 ( .a(FE_OFN1472_g52675_p), .o(g52528_sb) );
na03s02 TIMEBOOST_cell_72916 ( .a(n_2159), .b(g61812_sb), .c(g62004_db), .o(n_7887) );
in01s01 TIMEBOOST_cell_73866 ( .a(n_7883), .o(TIMEBOOST_net_23431) );
na02s01 TIMEBOOST_cell_37449 ( .a(TIMEBOOST_net_10336), .b(g65716_db), .o(n_1943) );
in01f02 g52529_u0 ( .a(FE_OFN1471_g52675_p), .o(g52529_sb) );
na02s01 TIMEBOOST_cell_37037 ( .a(TIMEBOOST_net_10130), .b(n_1817), .o(TIMEBOOST_net_558) );
na02f04 TIMEBOOST_cell_26209 ( .a(conf_wb_err_addr_in_951), .b(g53897_sb), .o(TIMEBOOST_net_7209) );
na03s01 TIMEBOOST_cell_64389 ( .a(TIMEBOOST_net_14021), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_410), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q), .o(TIMEBOOST_net_17567) );
in01f01 g52530_u0 ( .a(FE_OFN1472_g52675_p), .o(g52530_sb) );
na02f01 TIMEBOOST_cell_62611 ( .a(TIMEBOOST_net_20252), .b(FE_OFN908_n_4734), .o(TIMEBOOST_net_16252) );
na02m06 TIMEBOOST_cell_63656 ( .a(FE_OFN679_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q), .o(TIMEBOOST_net_20814) );
in01f02 g52531_u0 ( .a(FE_OFN1471_g52675_p), .o(g52531_sb) );
na04f04 TIMEBOOST_cell_36838 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q), .b(FE_OFN1404_n_8567), .c(n_9060), .d(g57322_sb), .o(n_10400) );
na02s01 TIMEBOOST_cell_48819 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q), .b(FE_OFN235_n_9834), .o(TIMEBOOST_net_14627) );
in01f02 g52532_u0 ( .a(FE_OFN1471_g52675_p), .o(g52532_sb) );
na04f04 TIMEBOOST_cell_36839 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q), .b(FE_OFN1373_n_8567), .c(n_9412), .d(g57404_sb), .o(n_11337) );
na02s01 TIMEBOOST_cell_52375 ( .a(configuration_wb_err_addr_538), .b(conf_wb_err_addr_in_947), .o(TIMEBOOST_net_16405) );
na02f02 TIMEBOOST_cell_62742 ( .a(FE_OFN1011_n_4734), .b(TIMEBOOST_net_12404), .o(TIMEBOOST_net_20318) );
in01f02 g52533_u0 ( .a(FE_OFN1471_g52675_p), .o(g52533_sb) );
na02f01 TIMEBOOST_cell_51911 ( .a(TIMEBOOST_net_12339), .b(FE_OFN989_n_574), .o(TIMEBOOST_net_16173) );
na02m02 TIMEBOOST_cell_53807 ( .a(n_3667), .b(n_65), .o(TIMEBOOST_net_17121) );
na03f02 TIMEBOOST_cell_70250 ( .a(n_4728), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q), .c(FE_OFN1097_g64577_p), .o(TIMEBOOST_net_22333) );
in01f02 g52534_u0 ( .a(FE_OFN1471_g52675_p), .o(g52534_sb) );
na03s01 TIMEBOOST_cell_67600 ( .a(TIMEBOOST_net_14631), .b(FE_OFN247_n_9112), .c(TIMEBOOST_net_14862), .o(TIMEBOOST_net_9518) );
na03f02 TIMEBOOST_cell_34980 ( .a(TIMEBOOST_net_9418), .b(FE_OFN1381_n_8567), .c(g57107_sb), .o(n_10479) );
ao12f02 g52543_u0 ( .a(pci_target_unit_pci_target_sm_backoff), .b(n_14529), .c(FE_OFN191_n_1193), .o(n_14586) );
no02f01 g52544_u0 ( .a(n_14663), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in), .o(n_14764) );
no02s01 g52545_u0 ( .a(pci_perr_i), .b(out_bckp_perr_en_out), .o(n_14624) );
na04f04 TIMEBOOST_cell_24836 ( .a(wbu_addr_in_265), .b(g52600_sb), .c(g52600_db), .d(TIMEBOOST_net_773), .o(n_11871) );
ao12f02 g52547_u0 ( .a(n_8564), .b(n_1185), .c(pci_target_unit_wbm_sm_pciw_fifo_control_in_84), .o(n_14694) );
na02m02 TIMEBOOST_cell_71151 ( .a(TIMEBOOST_net_22783), .b(FE_OFN1634_n_9531), .o(TIMEBOOST_net_21014) );
ao12f02 g52549_u0 ( .a(n_8582), .b(n_1101), .c(FE_OFN2198_n_10256), .o(n_10281) );
ao12f02 g52550_u0 ( .a(wishbone_slave_unit_del_sync_req_comp_pending_sample), .b(n_14620), .c(wishbone_slave_unit_del_sync_req_done_reg), .o(n_14623) );
ao22f02 g52551_u0 ( .a(n_671), .b(n_14689), .c(n_14688), .d(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in), .o(n_14691) );
ao22f02 g52552_u0 ( .a(n_661), .b(n_14689), .c(n_14688), .d(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50), .o(n_14690) );
ao12f02 g52554_u0 ( .a(n_14731), .b(n_14800), .c(wbm_dat_o_0_), .o(n_14802) );
ao12f02 g52556_u0 ( .a(n_14728), .b(n_16306), .c(wbm_dat_o_11_), .o(n_14799) );
ao12f02 g52557_u0 ( .a(n_14727), .b(n_14800), .c(wbm_dat_o_12_), .o(n_14798) );
ao12f02 g52558_u0 ( .a(n_14726), .b(n_16306), .c(wbm_dat_o_13_), .o(n_14797) );
ao12f02 g52559_u0 ( .a(n_14724), .b(n_16306), .c(wbm_dat_o_14_), .o(n_14796) );
ao12f02 g52560_u0 ( .a(n_14670), .b(n_14800), .c(wbm_dat_o_15_), .o(n_14763) );
ao12f02 g52561_u0 ( .a(n_14723), .b(n_14800), .c(wbm_dat_o_16_), .o(n_14794) );
ao12f02 g52562_u0 ( .a(n_14722), .b(n_14800), .c(wbm_dat_o_17_), .o(n_14793) );
ao12m02 g52563_u0 ( .a(n_14669), .b(n_16306), .c(wbm_dat_o_18_), .o(n_14762) );
ao12f02 g52564_u0 ( .a(n_14721), .b(n_16306), .c(wbm_dat_o_19_), .o(n_14792) );
ao12f02 g52565_u0 ( .a(n_14719), .b(n_14800), .c(wbm_dat_o_1_), .o(n_14791) );
ao12f02 g52566_u0 ( .a(n_14717), .b(n_16306), .c(wbm_dat_o_20_), .o(n_14790) );
ao12f02 g52567_u0 ( .a(n_14715), .b(n_14800), .c(wbm_dat_o_21_), .o(n_14789) );
ao12f02 g52569_u0 ( .a(n_14713), .b(n_14800), .c(wbm_dat_o_23_), .o(n_14786) );
ao12f02 g52570_u0 ( .a(n_14711), .b(n_14800), .c(wbm_dat_o_24_), .o(n_14784) );
ao12f02 g52571_u0 ( .a(n_14710), .b(n_16306), .c(wbm_dat_o_25_), .o(n_14783) );
ao12f02 g52572_u0 ( .a(n_14709), .b(n_16306), .c(wbm_dat_o_26_), .o(n_14781) );
ao12f02 g52573_u0 ( .a(n_14708), .b(n_16306), .c(wbm_dat_o_27_), .o(n_14780) );
ao12f02 g52574_u0 ( .a(n_14706), .b(n_16306), .c(wbm_dat_o_28_), .o(n_14778) );
ao12f02 g52575_u0 ( .a(n_14705), .b(n_16306), .c(wbm_dat_o_29_), .o(n_14777) );
ao12f02 g52576_u0 ( .a(n_14703), .b(n_16306), .c(wbm_dat_o_2_), .o(n_14776) );
ao12m02 g52577_u0 ( .a(n_14702), .b(n_16306), .c(wbm_dat_o_30_), .o(n_14775) );
ao12f02 g52578_u0 ( .a(n_14701), .b(n_16306), .c(wbm_dat_o_31_), .o(n_14773) );
ao12f02 g52579_u0 ( .a(n_14700), .b(n_14800), .c(wbm_dat_o_3_), .o(n_14772) );
ao12f02 g52580_u0 ( .a(n_14699), .b(n_14800), .c(wbm_dat_o_4_), .o(n_14770) );
ao12f02 g52581_u0 ( .a(n_14698), .b(n_14800), .c(wbm_dat_o_5_), .o(n_14769) );
ao12f02 g52582_u0 ( .a(n_14697), .b(n_14800), .c(wbm_dat_o_6_), .o(n_14768) );
ao12f02 g52583_u0 ( .a(n_14668), .b(n_16306), .c(wbm_dat_o_7_), .o(n_14761) );
ao12f02 g52584_u0 ( .a(n_14696), .b(n_16306), .c(wbm_dat_o_8_), .o(n_14767) );
ao12m02 g52585_u0 ( .a(n_14695), .b(n_14800), .c(wbm_dat_o_9_), .o(n_14766) );
ao12f02 g52586_u0 ( .a(n_14667), .b(n_16306), .c(wbm_sel_o_0_), .o(n_14760) );
ao12f02 g52587_u0 ( .a(n_14666), .b(n_16306), .c(wbm_sel_o_1_), .o(n_14759) );
ao12f02 g52588_u0 ( .a(n_14665), .b(n_16306), .c(wbm_sel_o_2_), .o(n_14757) );
ao12f02 g52589_u0 ( .a(n_14664), .b(n_16306), .c(wbm_sel_o_3_), .o(n_14756) );
in01m01 g52590_u0 ( .a(n_8757), .o(g52590_sb) );
na03m08 TIMEBOOST_cell_72676 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q), .b(g57991_sb), .c(TIMEBOOST_net_14386), .o(TIMEBOOST_net_16844) );
na02f01 TIMEBOOST_cell_68541 ( .a(TIMEBOOST_net_21478), .b(FE_OFN651_n_4508), .o(TIMEBOOST_net_14442) );
na02f02 TIMEBOOST_cell_49868 ( .a(TIMEBOOST_net_15151), .b(g63571_sb), .o(n_4111) );
in01m01 g52591_u0 ( .a(n_8757), .o(g52591_sb) );
na04s04 TIMEBOOST_cell_72664 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(FE_OFN1015_n_2053), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q), .d(g65877_sb), .o(n_1867) );
na02s01 TIMEBOOST_cell_68239 ( .a(TIMEBOOST_net_21327), .b(g63590_db), .o(n_3315) );
in01m01 g52592_u0 ( .a(n_8757), .o(g52592_sb) );
na02s02 TIMEBOOST_cell_48944 ( .a(TIMEBOOST_net_14689), .b(g63601_db), .o(TIMEBOOST_net_13016) );
in01m01 g52593_u0 ( .a(n_8757), .o(g52593_sb) );
na02s01 TIMEBOOST_cell_28945 ( .a(n_2273), .b(wbu_addr_in_254), .o(TIMEBOOST_net_8577) );
na04f02 TIMEBOOST_cell_73679 ( .a(n_8569), .b(wishbone_slave_unit_pcim_if_del_burst_in), .c(TIMEBOOST_net_400), .d(n_8568), .o(n_8843) );
in01f02 g52594_u0 ( .a(n_10256), .o(g52594_sb) );
na03m02 TIMEBOOST_cell_73192 ( .a(TIMEBOOST_net_23289), .b(g62029_sb), .c(TIMEBOOST_net_22358), .o(n_7838) );
na02f01 TIMEBOOST_cell_70686 ( .a(TIMEBOOST_net_13095), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_22551) );
in01f02 g52595_u0 ( .a(FE_OFN2198_n_10256), .o(g52595_sb) );
in01s01 TIMEBOOST_cell_73867 ( .a(TIMEBOOST_net_23431), .o(TIMEBOOST_net_23432) );
na02m01 TIMEBOOST_cell_69116 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_21766) );
na02m01 TIMEBOOST_cell_62710 ( .a(n_3739), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q), .o(TIMEBOOST_net_20302) );
in01f02 g52596_u0 ( .a(FE_OFN2198_n_10256), .o(g52596_sb) );
na03m04 TIMEBOOST_cell_72725 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q), .b(g64879_sb), .c(TIMEBOOST_net_14288), .o(TIMEBOOST_net_17511) );
na03f02 TIMEBOOST_cell_72956 ( .a(pci_target_unit_del_sync_addr_in_227), .b(g65222_sb), .c(TIMEBOOST_net_5410), .o(n_2665) );
in01f01 g52597_u0 ( .a(n_8935), .o(g52597_sb) );
na04f02 TIMEBOOST_cell_36833 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q), .b(FE_OFN1394_n_8567), .c(n_9082), .d(g57238_sb), .o(n_10430) );
na02f02 g52597_u2 ( .a(n_3169), .b(n_8935), .o(g52597_db) );
na04f04 TIMEBOOST_cell_36840 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q), .b(FE_OFN1394_n_8567), .c(n_9696), .d(g57347_sb), .o(n_11403) );
in01f02 g52598_u0 ( .a(FE_OFN2200_n_10256), .o(g52598_sb) );
na03f02 TIMEBOOST_cell_73143 ( .a(TIMEBOOST_net_23244), .b(g64246_sb), .c(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_22483) );
na02m01 TIMEBOOST_cell_68940 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q), .o(TIMEBOOST_net_21678) );
in01f02 g52599_u0 ( .a(FE_OFN2200_n_10256), .o(g52599_sb) );
na02s02 TIMEBOOST_cell_63820 ( .a(configuration_wb_err_cs_bit_566), .b(TIMEBOOST_net_13845), .o(TIMEBOOST_net_20896) );
na02s02 TIMEBOOST_cell_49438 ( .a(TIMEBOOST_net_14936), .b(g58049_db), .o(TIMEBOOST_net_9377) );
in01f01 g52600_u0 ( .a(n_8935), .o(g52600_sb) );
na02m01 TIMEBOOST_cell_62610 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_151), .o(TIMEBOOST_net_20252) );
na02f02 g52600_u2 ( .a(n_3151), .b(n_8935), .o(g52600_db) );
in01f02 g52601_u0 ( .a(FE_OFN2200_n_10256), .o(g52601_sb) );
no02s01 TIMEBOOST_cell_45481 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360), .b(FE_RN_728_0), .o(TIMEBOOST_net_13635) );
na03f02 TIMEBOOST_cell_73193 ( .a(TIMEBOOST_net_23293), .b(FE_OFN1092_g64577_p), .c(g63560_sb), .o(n_4114) );
in01f02 g52602_u0 ( .a(FE_OFN2200_n_10256), .o(g52602_sb) );
na04m06 TIMEBOOST_cell_72976 ( .a(n_4470), .b(g64947_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q), .d(g64947_db), .o(TIMEBOOST_net_13372) );
na03f02 TIMEBOOST_cell_64641 ( .a(TIMEBOOST_net_14141), .b(g64202_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q), .o(TIMEBOOST_net_13071) );
in01f02 g52603_u0 ( .a(FE_OFN2200_n_10256), .o(g52603_sb) );
na02m04 TIMEBOOST_cell_43571 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_140), .o(TIMEBOOST_net_12680) );
no04f04 TIMEBOOST_cell_73692 ( .a(FE_RN_396_0), .b(FE_OFN1710_n_4868), .c(FE_RN_130_0), .d(n_13577), .o(g53017_p) );
na03s02 TIMEBOOST_cell_72901 ( .a(n_1586), .b(g61925_sb), .c(g61925_db), .o(n_7973) );
in01f02 g52604_u0 ( .a(n_10256), .o(g52604_sb) );
na04f02 TIMEBOOST_cell_36841 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q), .b(FE_OFN1394_n_8567), .c(n_9500), .d(g57448_sb), .o(n_11285) );
na02s01 TIMEBOOST_cell_47875 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q), .o(TIMEBOOST_net_14155) );
na03s02 TIMEBOOST_cell_41912 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q), .b(g58345_sb), .c(g58345_db), .o(n_9475) );
in01f02 g52605_u0 ( .a(FE_OFN2200_n_10256), .o(g52605_sb) );
na03f02 TIMEBOOST_cell_66517 ( .a(g53909_sb), .b(FE_OFN1326_n_13547), .c(TIMEBOOST_net_16810), .o(n_13532) );
na03f02 TIMEBOOST_cell_64639 ( .a(TIMEBOOST_net_14139), .b(g64128_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_13072) );
na02m04 TIMEBOOST_cell_68652 ( .a(g64840_sb), .b(n_75), .o(TIMEBOOST_net_21534) );
in01f01 g52606_u0 ( .a(n_8935), .o(g52606_sb) );
na02f02 g52606_u2 ( .a(n_3487), .b(n_8935), .o(g52606_db) );
na03s02 TIMEBOOST_cell_41914 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q), .b(g58361_sb), .c(g58361_db), .o(n_9462) );
in01f02 g52607_u0 ( .a(FE_OFN2200_n_10256), .o(g52607_sb) );
na02f02 TIMEBOOST_cell_27788 ( .a(TIMEBOOST_net_7998), .b(n_14390), .o(n_14396) );
no03f10 TIMEBOOST_cell_68084 ( .a(n_16538), .b(n_15744), .c(n_16290), .o(TIMEBOOST_net_21250) );
in01f02 g52608_u0 ( .a(FE_OFN2198_n_10256), .o(g52608_sb) );
in01s01 TIMEBOOST_cell_45907 ( .a(TIMEBOOST_net_13919), .o(TIMEBOOST_net_13868) );
na02s01 TIMEBOOST_cell_26409 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_793), .b(n_12595), .o(TIMEBOOST_net_7309) );
in01f02 g52609_u0 ( .a(FE_OFN2198_n_10256), .o(g52609_sb) );
na03f02 TIMEBOOST_cell_65890 ( .a(n_4013), .b(g62805_sb), .c(g62805_db), .o(n_5371) );
in01s01 TIMEBOOST_cell_45908 ( .a(TIMEBOOST_net_13868), .o(TIMEBOOST_net_13869) );
in01f02 g52610_u0 ( .a(FE_OFN2200_n_10256), .o(g52610_sb) );
na03f02 TIMEBOOST_cell_65884 ( .a(n_4001), .b(g62773_sb), .c(g62773_db), .o(n_5448) );
na03f02 TIMEBOOST_cell_71064 ( .a(n_1871), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q), .c(FE_OFN1215_n_4151), .o(TIMEBOOST_net_22740) );
in01f02 g52611_u0 ( .a(FE_OFN2200_n_10256), .o(g52611_sb) );
na03m02 TIMEBOOST_cell_72559 ( .a(TIMEBOOST_net_21376), .b(FE_OFN628_n_4454), .c(TIMEBOOST_net_21534), .o(TIMEBOOST_net_20524) );
in01f02 g52612_u0 ( .a(FE_OFN2200_n_10256), .o(g52612_sb) );
na02f01 TIMEBOOST_cell_40257 ( .a(TIMEBOOST_net_11740), .b(FE_OFN1082_n_13221), .o(TIMEBOOST_net_645) );
na02f01 TIMEBOOST_cell_26417 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_794), .b(n_12595), .o(TIMEBOOST_net_7313) );
oa22f02 g52613_u0 ( .a(FE_OFN2198_n_10256), .b(wbu_addr_in_278), .c(n_10155), .d(n_4208), .o(n_10170) );
in01f01 g52614_u0 ( .a(n_8935), .o(g52614_sb) );
in01s01 TIMEBOOST_cell_45909 ( .a(TIMEBOOST_net_13870), .o(TIMEBOOST_net_5289) );
na03m02 TIMEBOOST_cell_72806 ( .a(n_4476), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q), .c(TIMEBOOST_net_9704), .o(TIMEBOOST_net_17433) );
na03m02 TIMEBOOST_cell_72576 ( .a(TIMEBOOST_net_17212), .b(FE_OFN664_n_4495), .c(TIMEBOOST_net_21532), .o(TIMEBOOST_net_13236) );
oa22f02 g52615_u0 ( .a(FE_OFN2198_n_10256), .b(wbu_addr_in_280), .c(n_10155), .d(n_4196), .o(n_10157) );
in01f02 g52616_u0 ( .a(FE_OFN2198_n_10256), .o(g52616_sb) );
in01s01 TIMEBOOST_cell_45910 ( .a(TIMEBOOST_net_13871), .o(TIMEBOOST_net_13870) );
in01f02 g52617_u0 ( .a(n_10256), .o(g52617_sb) );
in01s01 TIMEBOOST_cell_45911 ( .a(pci_target_unit_fifos_pcir_data_in_174), .o(TIMEBOOST_net_13872) );
na02s02 TIMEBOOST_cell_63305 ( .a(TIMEBOOST_net_20599), .b(g58207_db), .o(TIMEBOOST_net_9373) );
in01f02 g52618_u0 ( .a(n_10256), .o(g52618_sb) );
in01s01 TIMEBOOST_cell_45912 ( .a(TIMEBOOST_net_13872), .o(TIMEBOOST_net_13873) );
na02f02 TIMEBOOST_cell_40549 ( .a(TIMEBOOST_net_11886), .b(g52645_sb), .o(TIMEBOOST_net_5667) );
na02m02 TIMEBOOST_cell_72122 ( .a(TIMEBOOST_net_16307), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_23269) );
in01f02 g52619_u0 ( .a(n_10256), .o(g52619_sb) );
na02s01 TIMEBOOST_cell_47723 ( .a(TIMEBOOST_net_10175), .b(FE_OFN945_n_2248), .o(TIMEBOOST_net_14079) );
na02f01 TIMEBOOST_cell_37344 ( .a(n_2171), .b(FE_OFN992_n_2373), .o(TIMEBOOST_net_10284) );
in01f02 g52620_u0 ( .a(FE_OFN2198_n_10256), .o(g52620_sb) );
na04f04 TIMEBOOST_cell_24799 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q), .b(g58803_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q), .d(FE_OFN2157_n_16439), .o(n_8638) );
na02m04 TIMEBOOST_cell_68691 ( .a(TIMEBOOST_net_21553), .b(n_3755), .o(TIMEBOOST_net_10727) );
na02f01 TIMEBOOST_cell_69894 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(g63547_sb), .o(TIMEBOOST_net_22155) );
in01f02 g52621_u0 ( .a(n_10256), .o(g52621_sb) );
na02s01 TIMEBOOST_cell_47725 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q), .b(FE_OFN205_n_9140), .o(TIMEBOOST_net_14080) );
na04m04 TIMEBOOST_cell_73278 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q), .b(FE_OFN1812_n_7845), .c(n_1602), .d(g61828_sb), .o(n_8130) );
na02s02 TIMEBOOST_cell_43149 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q), .o(TIMEBOOST_net_12469) );
in01f02 g52622_u0 ( .a(FE_OFN2198_n_10256), .o(g52622_sb) );
na04f04 TIMEBOOST_cell_24801 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q), .b(g58801_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q), .d(FE_OFN2153_n_16439), .o(n_8641) );
no02f04 g52623_u0 ( .a(wbu_addr_in_251), .b(FE_OFN2198_n_10256), .o(g52623_p) );
ao12f02 g52623_u1 ( .a(g52623_p), .b(wbu_addr_in_251), .c(FE_OFN2198_n_10256), .o(n_10106) );
in01f04 g52624_u0 ( .a(n_16748), .o(g52624_sb) );
na02s01 TIMEBOOST_cell_29009 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q), .o(TIMEBOOST_net_8609) );
na02f02 TIMEBOOST_cell_70239 ( .a(TIMEBOOST_net_22327), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_16820) );
na03m02 TIMEBOOST_cell_72590 ( .a(TIMEBOOST_net_21433), .b(g64771_sb), .c(TIMEBOOST_net_21633), .o(TIMEBOOST_net_20534) );
in01f01 g52625_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52625_sb) );
na02f01 TIMEBOOST_cell_71552 ( .a(TIMEBOOST_net_13568), .b(n_11977), .o(TIMEBOOST_net_22984) );
na03s02 TIMEBOOST_cell_72375 ( .a(TIMEBOOST_net_10425), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q), .c(FE_OFN955_n_1699), .o(TIMEBOOST_net_17244) );
na02s01 TIMEBOOST_cell_47936 ( .a(TIMEBOOST_net_14185), .b(g58026_sb), .o(TIMEBOOST_net_12770) );
in01f01 g52626_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52626_sb) );
na04f04 TIMEBOOST_cell_24814 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q), .b(g58823_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q), .d(FE_OFN2157_n_16439), .o(n_8618) );
in01m02 g52627_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52627_sb) );
na04f04 TIMEBOOST_cell_24816 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q), .b(g58821_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q), .d(FE_OFN2153_n_16439), .o(n_8620) );
in01f02 g52628_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52628_sb) );
na04f04 TIMEBOOST_cell_24181 ( .a(n_9725), .b(g57208_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q), .d(FE_OFN1423_n_8567), .o(n_11548) );
na04m04 TIMEBOOST_cell_73068 ( .a(n_2209), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q), .c(FE_OFN702_n_7845), .d(g61711_sb), .o(n_8404) );
in01f02 g52629_u0 ( .a(n_16748), .o(g52629_sb) );
in01f04 g52630_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52630_sb) );
in01s01 TIMEBOOST_cell_45913 ( .a(TIMEBOOST_net_13923), .o(TIMEBOOST_net_13874) );
na03f06 TIMEBOOST_cell_73335 ( .a(TIMEBOOST_net_20485), .b(FE_OCPN1911_FE_OFN1152_n_13249), .c(g54143_sb), .o(n_13361) );
na03s02 TIMEBOOST_cell_41916 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q), .b(g58364_sb), .c(g58364_db), .o(n_9460) );
in01f02 g52631_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52631_sb) );
na03f02 TIMEBOOST_cell_66908 ( .a(FE_OFN1736_n_16317), .b(TIMEBOOST_net_16003), .c(FE_OFN1742_n_11019), .o(n_12523) );
in01f04 g52632_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52632_sb) );
na03f02 TIMEBOOST_cell_35053 ( .a(TIMEBOOST_net_9605), .b(FE_OFN1436_n_9372), .c(g58467_sb), .o(n_9381) );
na02m04 TIMEBOOST_cell_69518 ( .a(g65001_sb), .b(n_84), .o(TIMEBOOST_net_21967) );
in01f01 g52633_u0 ( .a(n_16748), .o(g52633_sb) );
na02f01 TIMEBOOST_cell_54070 ( .a(TIMEBOOST_net_17252), .b(FE_OFN1049_n_16657), .o(TIMEBOOST_net_14710) );
in01m02 g52634_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52634_sb) );
na04f04 TIMEBOOST_cell_24818 ( .a(n_16984), .b(n_16985), .c(n_9997), .d(n_10584), .o(n_12139) );
na02f02 TIMEBOOST_cell_71078 ( .a(TIMEBOOST_net_17389), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_22747) );
na02f02 TIMEBOOST_cell_50226 ( .a(TIMEBOOST_net_15330), .b(g62959_sb), .o(n_5964) );
in01f02 g52635_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52635_sb) );
na02s02 TIMEBOOST_cell_54057 ( .a(g65751_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q), .o(TIMEBOOST_net_17246) );
na02s01 TIMEBOOST_cell_47512 ( .a(TIMEBOOST_net_13973), .b(g67042_sb), .o(n_1275) );
na03f02 TIMEBOOST_cell_72377 ( .a(n_13784), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_392), .c(TIMEBOOST_net_11103), .o(TIMEBOOST_net_21413) );
in01m02 g52636_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52636_sb) );
na04f04 TIMEBOOST_cell_36862 ( .a(TIMEBOOST_net_8578), .b(n_10256), .c(g52617_sb), .d(TIMEBOOST_net_712), .o(n_11853) );
in01m06 g52637_u0 ( .a(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52637_sb) );
in01s01 TIMEBOOST_cell_45914 ( .a(TIMEBOOST_net_13874), .o(TIMEBOOST_net_13875) );
na03f02 TIMEBOOST_cell_66941 ( .a(FE_OFN1753_n_12086), .b(FE_OFN1568_n_11027), .c(TIMEBOOST_net_13619), .o(n_12635) );
in01m02 g52638_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52638_sb) );
na02s01 TIMEBOOST_cell_29371 ( .a(parchk_pci_ad_out_in_1193), .b(configuration_wb_err_data_596), .o(TIMEBOOST_net_8790) );
na02f01 g52638_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52638_db) );
na03f02 TIMEBOOST_cell_47428 ( .a(FE_OFN1587_n_13736), .b(TIMEBOOST_net_13742), .c(FE_OCP_RBN1997_n_13971), .o(n_14256) );
in01f01 g52639_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52639_sb) );
na04f04 TIMEBOOST_cell_34715 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q), .b(FE_OFN1349_n_8567), .c(n_9737), .d(g57187_sb), .o(n_11565) );
na02m04 TIMEBOOST_cell_53133 ( .a(n_3754), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q), .o(TIMEBOOST_net_16784) );
na03m02 TIMEBOOST_cell_70374 ( .a(FE_OFN2021_n_4778), .b(TIMEBOOST_net_16649), .c(TIMEBOOST_net_637), .o(TIMEBOOST_net_22395) );
in01m01 g52641_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52641_sb) );
in01f01 g52642_u0 ( .a(n_16748), .o(g52642_sb) );
na02s02 TIMEBOOST_cell_48898 ( .a(TIMEBOOST_net_14666), .b(g58106_sb), .o(TIMEBOOST_net_9431) );
in01s01 TIMEBOOST_cell_72355 ( .a(TIMEBOOST_net_23387), .o(TIMEBOOST_net_23388) );
in01f02 g52643_u0 ( .a(n_16748), .o(g52643_sb) );
na04m04 TIMEBOOST_cell_67585 ( .a(TIMEBOOST_net_20419), .b(FE_OFN580_n_9531), .c(g58376_sb), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q), .o(TIMEBOOST_net_9467) );
in01f01 g52644_u0 ( .a(n_16748), .o(g52644_sb) );
na02s02 TIMEBOOST_cell_37362 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(g65755_sb), .o(TIMEBOOST_net_10293) );
na04f04 TIMEBOOST_cell_73116 ( .a(FE_OFN2052_n_6965), .b(FE_OFN2121_n_2687), .c(n_4084), .d(FE_OFN2245_n_4792), .o(n_7210) );
in01m01 g52645_u0 ( .a(n_16748), .o(g52645_sb) );
na03f02 TIMEBOOST_cell_24998 ( .a(n_11002), .b(FE_RN_468_0), .c(n_12590), .o(n_12852) );
na03m02 TIMEBOOST_cell_72915 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q), .b(g65868_sb), .c(g65868_db), .o(n_2054) );
in01m01 g52646_u0 ( .a(n_16748), .o(g52646_sb) );
na03m02 TIMEBOOST_cell_68544 ( .a(TIMEBOOST_net_16880), .b(g65269_sb), .c(wishbone_slave_unit_pcim_sm_be_in_557), .o(TIMEBOOST_net_21480) );
na02m04 TIMEBOOST_cell_69468 ( .a(g64990_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q), .o(TIMEBOOST_net_21942) );
na03f02 TIMEBOOST_cell_73766 ( .a(TIMEBOOST_net_13704), .b(FE_OFN1774_n_13800), .c(FE_OFN1771_n_14054), .o(g74879_p) );
in01m01 g52647_u0 ( .a(FE_OFN697_n_16760), .o(g52647_sb) );
na02m02 TIMEBOOST_cell_68824 ( .a(FE_OFN620_n_4490), .b(n_36), .o(TIMEBOOST_net_21620) );
na02f01 TIMEBOOST_cell_54444 ( .a(TIMEBOOST_net_17439), .b(FE_OFN1242_n_4092), .o(TIMEBOOST_net_15529) );
na03f20 TIMEBOOST_cell_72400 ( .a(TIMEBOOST_net_12251), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in_417), .c(n_398), .o(n_13541) );
in01f01 g52648_u0 ( .a(n_16748), .o(g52648_sb) );
na03m02 TIMEBOOST_cell_72648 ( .a(TIMEBOOST_net_21490), .b(g64914_sb), .c(TIMEBOOST_net_21671), .o(TIMEBOOST_net_17098) );
na03f02 TIMEBOOST_cell_73069 ( .a(TIMEBOOST_net_22035), .b(FE_OFN2084_n_8407), .c(g61826_sb), .o(n_8135) );
na02m01 TIMEBOOST_cell_68545 ( .a(TIMEBOOST_net_21480), .b(n_5641), .o(TIMEBOOST_net_20895) );
na02s01 TIMEBOOST_cell_68187 ( .a(TIMEBOOST_net_21301), .b(FE_OFN938_n_2292), .o(TIMEBOOST_net_10254) );
na03f01 TIMEBOOST_cell_66290 ( .a(n_3763), .b(g62366_sb), .c(g62366_db), .o(n_6869) );
in01f04 g52650_u0 ( .a(n_16748), .o(g52650_sb) );
na02f02 TIMEBOOST_cell_70639 ( .a(TIMEBOOST_net_22527), .b(g54320_sb), .o(n_13287) );
na02f04 g52650_u2 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55), .b(n_16748), .o(g52650_db) );
in01f01 g52651_u0 ( .a(n_16748), .o(g52651_sb) );
na02m02 TIMEBOOST_cell_68131 ( .a(TIMEBOOST_net_21273), .b(g54219_sb), .o(TIMEBOOST_net_14037) );
in01f02 g52652_u0 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(g52652_sb) );
na03f02 TIMEBOOST_cell_24014 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q), .b(g59113_sb), .c(TIMEBOOST_net_5533), .o(n_8699) );
na03m08 TIMEBOOST_cell_64810 ( .a(n_3777), .b(FE_OFN620_n_4490), .c(n_17), .o(TIMEBOOST_net_16241) );
na02f02 TIMEBOOST_cell_70681 ( .a(TIMEBOOST_net_22548), .b(g62739_sb), .o(n_5501) );
in01f01 g52653_u0 ( .a(n_16748), .o(g52653_sb) );
na02m02 TIMEBOOST_cell_68408 ( .a(n_3780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q), .o(TIMEBOOST_net_21412) );
na02m04 TIMEBOOST_cell_72102 ( .a(g64210_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q), .o(TIMEBOOST_net_23259) );
no02f08 g52675_u0 ( .a(n_8872), .b(n_16945), .o(g52675_p) );
na02f02 g52677_u0 ( .a(n_14517), .b(n_14615), .o(n_14629) );
no02f02 g52678_u0 ( .a(n_14725), .b(n_14659), .o(n_14731) );
no02f02 g52679_u0 ( .a(n_14725), .b(n_14658), .o(n_14730) );
no02m02 g52680_u0 ( .a(n_14725), .b(n_14657), .o(n_14728) );
no02m02 g52681_u0 ( .a(n_14725), .b(n_14656), .o(n_14727) );
no02f02 g52682_u0 ( .a(n_14725), .b(n_14655), .o(n_14726) );
no02f02 g52683_u0 ( .a(n_14725), .b(n_14654), .o(n_14724) );
no02f02 g52684_u0 ( .a(n_14725), .b(n_14627), .o(n_14670) );
no02f02 g52685_u0 ( .a(n_14725), .b(n_14653), .o(n_14723) );
no02f02 g52686_u0 ( .a(n_14725), .b(n_14652), .o(n_14722) );
no02m02 g52687_u0 ( .a(n_14725), .b(n_14626), .o(n_14669) );
no02m02 g52688_u0 ( .a(n_14725), .b(n_14651), .o(n_14721) );
no02m02 g52689_u0 ( .a(n_14725), .b(n_14650), .o(n_14719) );
no02m03 g52690_u0 ( .a(n_14725), .b(n_14649), .o(n_14717) );
no02f02 g52691_u0 ( .a(n_14725), .b(n_14648), .o(n_14715) );
no02f02 g52693_u0 ( .a(n_14725), .b(n_14646), .o(n_14713) );
no02f02 g52694_u0 ( .a(n_14725), .b(n_14645), .o(n_14711) );
no02f02 g52695_u0 ( .a(n_14725), .b(n_14644), .o(n_14710) );
no02f02 g52696_u0 ( .a(n_14725), .b(n_14643), .o(n_14709) );
no02f02 g52697_u0 ( .a(n_14725), .b(n_14642), .o(n_14708) );
no02f02 g52698_u0 ( .a(n_14725), .b(n_14641), .o(n_14706) );
no02f02 g52699_u0 ( .a(n_14725), .b(n_14640), .o(n_14705) );
no02f02 g52700_u0 ( .a(n_14725), .b(n_14639), .o(n_14703) );
no02f02 g52701_u0 ( .a(n_14725), .b(n_14638), .o(n_14702) );
no02m03 g52702_u0 ( .a(n_14725), .b(n_14637), .o(n_14701) );
no02f02 g52703_u0 ( .a(n_14725), .b(n_14636), .o(n_14700) );
no02m03 g52704_u0 ( .a(n_14725), .b(n_14635), .o(n_14699) );
no02f02 g52705_u0 ( .a(n_14725), .b(n_14634), .o(n_14698) );
no02f02 g52706_u0 ( .a(n_14725), .b(n_14633), .o(n_14697) );
no02f02 g52707_u0 ( .a(n_14725), .b(n_14625), .o(n_14668) );
no02m02 g52708_u0 ( .a(n_14725), .b(n_14632), .o(n_14696) );
no02m02 g52709_u0 ( .a(n_14725), .b(n_14631), .o(n_14695) );
no02f04 g52710_u0 ( .a(n_16306), .b(pci_target_unit_wbm_sm_pciw_fifo_cbe_in), .o(n_14667) );
no02f04 g52711_u0 ( .a(n_16306), .b(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81), .o(n_14666) );
no02f04 g52712_u0 ( .a(n_16306), .b(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82), .o(n_14665) );
no02f04 g52713_u0 ( .a(n_16306), .b(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83), .o(n_14664) );
na02f02 g52714_u0 ( .a(n_1532), .b(n_14620), .o(g52714_p) );
in01f02 g52714_u1 ( .a(g52714_p), .o(n_14621) );
oa12f01 g52715_u0 ( .a(n_10155), .b(wbs_stb_i), .c(n_779), .o(n_10441) );
na02s06 TIMEBOOST_cell_53951 ( .a(wbs_dat_i_3_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q), .o(TIMEBOOST_net_17193) );
na04f04 TIMEBOOST_cell_24161 ( .a(n_9751), .b(g57173_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q), .d(FE_OFN1425_n_8567), .o(n_11583) );
ao12f02 g52718_u0 ( .a(n_14485), .b(n_13920), .c(n_2285), .o(n_14617) );
oa12f02 g52719_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_control_in_84), .b(n_1541), .c(n_1086), .o(n_14663) );
oa22f01 g52720_u0 ( .a(n_10792), .b(wbs_err_o), .c(wbs_stb_i), .d(n_471), .o(n_8874) );
in01s01 g52778_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in), .o(n_14659) );
in01s01 g52780_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59), .o(n_14658) );
in01s01 g52782_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60), .o(n_14657) );
in01s01 g52784_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61), .o(n_14656) );
in01s01 g52786_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62), .o(n_14655) );
in01s01 g52788_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63), .o(n_14654) );
in01s01 g52790_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64), .o(n_14627) );
in01s01 g52792_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65), .o(n_14653) );
in01s01 g52794_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66), .o(n_14652) );
in01s01 g52796_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67), .o(n_14626) );
in01s01 g52798_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68), .o(n_14651) );
in01s01 g52800_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50), .o(n_14650) );
in01s01 g52802_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69), .o(n_14649) );
in01s01 g52804_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70), .o(n_14648) );
in01s01 g52808_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72), .o(n_14646) );
in01s01 g52810_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73), .o(n_14645) );
in01s01 g52812_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74), .o(n_14644) );
in01s01 g52814_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75), .o(n_14643) );
in01s01 g52816_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76), .o(n_14642) );
in01s01 g52818_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77), .o(n_14641) );
in01s01 g52820_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78), .o(n_14640) );
in01s01 g52822_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51), .o(n_14639) );
in01s01 g52824_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79), .o(n_14638) );
in01s01 g52826_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80), .o(n_14637) );
in01s01 g52836_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52), .o(n_14636) );
in01s01 g52838_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53), .o(n_14635) );
in01s01 g52840_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54), .o(n_14634) );
in01s01 g52842_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55), .o(n_14633) );
in01s01 g52844_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56), .o(n_14625) );
in01s01 g52846_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57), .o(n_14632) );
in01s01 g52848_u0 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58), .o(n_14631) );
in01f20 g52853_u0 ( .a(n_10155), .o(n_10256) );
in01f20 g52862_u0 ( .a(n_8935), .o(n_10155) );
in01f10 g52863_u0 ( .a(n_8872), .o(n_8935) );
no02f10 g52864_u0 ( .a(n_17031), .b(n_17032), .o(n_8872) );
na02f02 g52865_u0 ( .a(n_14074), .b(n_14486), .o(g52865_p) );
in01f02 g52865_u1 ( .a(g52865_p), .o(n_14616) );
in01f01 g52866_u0 ( .a(n_14571), .o(n_14572) );
no02f02 g52867_u0 ( .a(n_14386), .b(parity_checker_pci_perr_en_reg), .o(n_14571) );
no02f04 g52869_u0 ( .a(n_14528), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .o(n_14620) );
in01f02 g52870_u0 ( .a(n_14490), .o(n_14531) );
ao12f02 g52871_u0 ( .a(n_14487), .b(FE_OFN1709_n_4868), .c(parchk_pci_ad_out_in_1198), .o(n_14490) );
in01f02 g52872_u0 ( .a(n_14489), .o(n_14530) );
ao12f02 g52873_u0 ( .a(n_14487), .b(FE_OFN1709_n_4868), .c(pci_ad_o_31_), .o(n_14489) );
ao12f02 g52874_u0 ( .a(n_14570), .b(n_14518), .c(n_14898), .o(n_14615) );
ao12f02 g52875_u0 ( .a(n_14385), .b(n_12168), .c(n_2629), .o(n_14529) );
in01f01 g52876_u0 ( .a(FE_OFN1705_n_4868), .o(g52876_sb) );
na02s01 TIMEBOOST_cell_43151 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q), .o(TIMEBOOST_net_12470) );
in01f01 g52877_u0 ( .a(FE_OFN1705_n_4868), .o(g52877_sb) );
na02f04 TIMEBOOST_cell_3611 ( .a(TIMEBOOST_net_365), .b(n_3221), .o(n_7818) );
na02m02 TIMEBOOST_cell_68890 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q), .b(FE_OFN1624_n_4438), .o(TIMEBOOST_net_21653) );
na02s02 TIMEBOOST_cell_71153 ( .a(TIMEBOOST_net_22784), .b(FE_OFN597_n_9694), .o(TIMEBOOST_net_10863) );
in01f01 g52878_u0 ( .a(FE_OFN1705_n_4868), .o(g52878_sb) );
na02m02 TIMEBOOST_cell_69391 ( .a(TIMEBOOST_net_21903), .b(g65048_sb), .o(TIMEBOOST_net_12688) );
na02f06 TIMEBOOST_cell_3604 ( .a(n_16524), .b(FE_OCPN1823_n_16560), .o(TIMEBOOST_net_362) );
in01m01 g52879_u0 ( .a(n_14389), .o(g52879_sb) );
na02m06 TIMEBOOST_cell_68662 ( .a(FE_OFN686_n_4417), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q), .o(TIMEBOOST_net_21539) );
na02m02 TIMEBOOST_cell_50707 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_387), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_15571) );
na02m02 TIMEBOOST_cell_70185 ( .a(TIMEBOOST_net_22300), .b(TIMEBOOST_net_20871), .o(TIMEBOOST_net_14739) );
in01m01 g52880_u0 ( .a(n_14389), .o(g52880_sb) );
na03f10 TIMEBOOST_cell_64310 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q), .b(n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_396), .o(TIMEBOOST_net_20878) );
in01m01 g52881_u0 ( .a(n_14389), .o(g52881_sb) );
na02f08 TIMEBOOST_cell_3605 ( .a(n_15915), .b(TIMEBOOST_net_362), .o(n_16273) );
na02f02 TIMEBOOST_cell_70418 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_22417) );
no02f02 g52890_u0 ( .a(n_13843), .b(n_14075), .o(n_14486) );
ao12f04 g52891_u0 ( .a(FE_OFN1709_n_4868), .b(n_13787), .c(n_13286), .o(n_14487) );
na02f02 g52892_u0 ( .a(n_13910), .b(n_1196), .o(n_14385) );
oa12f02 g52893_u0 ( .a(n_14073), .b(n_14484), .c(n_15370), .o(n_14528) );
in01f02 g52894_u0 ( .a(n_14104), .o(n_14384) );
na03m02 TIMEBOOST_cell_72896 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q), .b(g64293_sb), .c(TIMEBOOST_net_23235), .o(TIMEBOOST_net_22253) );
na02f02 g52897_u0 ( .a(n_14357), .b(n_7673), .o(n_14383) );
na02f02 g52898_u0 ( .a(n_14355), .b(n_7672), .o(n_14382) );
na02f02 g52899_u0 ( .a(n_14353), .b(n_7671), .o(n_14381) );
na02f02 g52900_u0 ( .a(n_14351), .b(n_7669), .o(n_14380) );
na02f02 g52901_u0 ( .a(n_7667), .b(n_14085), .o(n_14094) );
na02f02 g52902_u0 ( .a(n_14349), .b(n_7666), .o(n_14379) );
na02f02 g52903_u0 ( .a(n_14083), .b(n_7664), .o(n_14093) );
na02f02 g52904_u0 ( .a(n_14347), .b(n_7663), .o(n_14378) );
na02f02 g52905_u0 ( .a(n_14341), .b(n_7661), .o(n_14377) );
na02f02 g52907_u0 ( .a(n_14343), .b(n_7656), .o(n_14375) );
na02f02 g52908_u0 ( .a(n_14337), .b(n_7655), .o(n_14374) );
na02f02 g52909_u0 ( .a(n_14339), .b(n_7654), .o(n_14373) );
na02f02 g52910_u0 ( .a(n_14335), .b(n_7653), .o(n_14372) );
na02f02 g52911_u0 ( .a(n_14081), .b(n_7652), .o(n_14088) );
na02f02 g52912_u0 ( .a(n_7651), .b(n_14333), .o(n_14371) );
na02f02 g52913_u0 ( .a(n_7650), .b(n_14331), .o(n_14370) );
na02f02 g52914_u0 ( .a(n_7649), .b(n_14329), .o(n_14369) );
na02f02 g52915_u0 ( .a(n_7648), .b(n_14327), .o(n_14368) );
na02f02 g52916_u0 ( .a(n_7647), .b(n_14325), .o(n_14367) );
na02f02 g52917_u0 ( .a(n_14323), .b(n_7528), .o(n_14366) );
na02f02 g52918_u0 ( .a(n_14321), .b(n_7646), .o(n_14365) );
na02m04 TIMEBOOST_cell_72197 ( .a(TIMEBOOST_net_23306), .b(g64214_sb), .o(n_3955) );
na02f02 g52920_u0 ( .a(n_14319), .b(n_7636), .o(n_14364) );
na02f02 g52921_u0 ( .a(n_14315), .b(n_7509), .o(n_14363) );
na02f02 g52922_u0 ( .a(n_14317), .b(n_7505), .o(n_14362) );
na02f02 g52923_u0 ( .a(n_14313), .b(n_7522), .o(n_14361) );
na02f02 g52924_u0 ( .a(n_14311), .b(n_7521), .o(n_14360) );
na02f02 g52925_u0 ( .a(n_14309), .b(n_7519), .o(n_14359) );
na02f02 g52926_u0 ( .a(n_14357), .b(n_7629), .o(n_14358) );
na02f02 g52927_u0 ( .a(n_14355), .b(n_7518), .o(n_14356) );
na02f02 g52928_u0 ( .a(n_14353), .b(n_7645), .o(n_14354) );
na02f02 g52929_u0 ( .a(n_7517), .b(n_14085), .o(n_14086) );
na02f02 g52930_u0 ( .a(n_14351), .b(n_7643), .o(n_14352) );
na02f02 g52931_u0 ( .a(n_14349), .b(n_7524), .o(n_14350) );
na02f02 g52932_u0 ( .a(n_14083), .b(n_7516), .o(n_14084) );
na02f02 g52933_u0 ( .a(n_14347), .b(n_7515), .o(n_14348) );
na02f02 g52934_u0 ( .a(n_7514), .b(n_14345), .o(n_14346) );
na02f02 g52935_u0 ( .a(n_7640), .b(n_14343), .o(n_14344) );
na02f02 g52936_u0 ( .a(n_14341), .b(n_7525), .o(n_14342) );
na02f02 g52937_u0 ( .a(n_14339), .b(n_7665), .o(n_14340) );
na02f02 g52938_u0 ( .a(n_14337), .b(n_7639), .o(n_14338) );
na02f02 g52939_u0 ( .a(n_14335), .b(n_7532), .o(n_14336) );
na02f02 g52940_u0 ( .a(n_14081), .b(n_7513), .o(n_14082) );
na02f02 g52941_u0 ( .a(n_7512), .b(n_14333), .o(n_14334) );
na02f02 g52942_u0 ( .a(n_7534), .b(n_14331), .o(n_14332) );
na02f02 g52943_u0 ( .a(n_7535), .b(n_14329), .o(n_14330) );
na02f02 g52944_u0 ( .a(n_7511), .b(n_14327), .o(n_14328) );
na02f02 g52945_u0 ( .a(n_7638), .b(n_14325), .o(n_14326) );
na02f02 g52946_u0 ( .a(n_14323), .b(n_7510), .o(n_14324) );
na02f02 g52947_u0 ( .a(n_14321), .b(n_7637), .o(n_14322) );
na02f02 g52948_u0 ( .a(n_7735), .b(parchk_pci_serr_en_in), .o(n_14080) );
na02f02 g52949_u0 ( .a(n_14319), .b(n_7634), .o(n_14320) );
na02m04 TIMEBOOST_cell_70229 ( .a(TIMEBOOST_net_22322), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_15056) );
na02f02 g52951_u0 ( .a(n_14317), .b(n_7632), .o(n_14318) );
na02f02 g52952_u0 ( .a(n_14315), .b(n_7633), .o(n_14316) );
na02f02 g52953_u0 ( .a(n_14313), .b(n_7631), .o(n_14314) );
na02f02 g52954_u0 ( .a(n_14311), .b(n_7630), .o(n_14312) );
na02f02 g52955_u0 ( .a(n_14309), .b(n_7628), .o(n_14310) );
ao12f04 g52956_u0 ( .a(n_8595), .b(n_1979), .c(n_7567), .o(n_10792) );
ao12f02 g52957_u0 ( .a(n_14898), .b(n_14890), .c(n_112), .o(n_14570) );
na03f02 g52966_u0 ( .a(n_16610), .b(n_14283), .c(n_16611), .o(n_14607) );
na02f02 g52990_u0 ( .a(n_14539), .b(n_14521), .o(n_14583) );
na03f02 g52991_u0 ( .a(n_16615), .b(n_14413), .c(n_16614), .o(n_14582) );
na02f02 TIMEBOOST_cell_18226 ( .a(TIMEBOOST_net_5476), .b(n_4659), .o(n_6982) );
na02f40 g52_u0 ( .a(pciu_am1_in_528), .b(pciu_bar1_in_390), .o(g52_p) );
in01f20 g52_u1 ( .a(g52_p), .o(n_15598) );
in01s01 g53004_u0 ( .a(parchk_pci_perr_out_in), .o(n_14079) );
na02f02 g53010_u0 ( .a(n_14484), .b(n_1684), .o(n_14618) );
no02f04 g53011_u0 ( .a(n_13731), .b(FE_OFN1709_n_4868), .o(g53011_p) );
in01f02 g53011_u1 ( .a(g53011_p), .o(n_14085) );
in01f06 TIMEBOOST_cell_42691 ( .a(TIMEBOOST_net_12239), .o(n_545) );
in01f02 g53012_u1 ( .a(g53012_p), .o(n_14341) );
no02f02 g53014_u0 ( .a(n_13776), .b(FE_OFN1710_n_4868), .o(g53014_p) );
in01f02 g53014_u1 ( .a(g53014_p), .o(n_14343) );
no02f04 g53015_u0 ( .a(n_13775), .b(FE_OFN1709_n_4868), .o(g53015_p) );
in01f02 g53015_u1 ( .a(g53015_p), .o(n_14337) );
no02f04 g53016_u0 ( .a(n_13774), .b(FE_OFN1709_n_4868), .o(g53016_p) );
in01f02 g53016_u1 ( .a(g53016_p), .o(n_14339) );
in01f02 g53017_u1 ( .a(g53017_p), .o(n_14335) );
no02f04 g53018_u0 ( .a(n_13728), .b(FE_OFN1709_n_4868), .o(g53018_p) );
in01f02 g53018_u1 ( .a(g53018_p), .o(n_14081) );
no02f02 g53019_u0 ( .a(n_14481), .b(n_14302), .o(n_14569) );
no02f02 g53020_u0 ( .a(n_14479), .b(n_14300), .o(n_16594) );
no02f02 g53021_u0 ( .a(n_14298), .b(n_14477), .o(n_14567) );
no02f02 g53022_u0 ( .a(n_13772), .b(FE_OFN1705_n_4868), .o(g53022_p) );
in01f02 g53022_u1 ( .a(g53022_p), .o(n_14333) );
no02f02 g53023_u0 ( .a(n_14295), .b(n_14476), .o(n_14566) );
no02f02 g53024_u0 ( .a(n_14293), .b(n_14474), .o(n_14565) );
no02f02 g53025_u0 ( .a(n_14472), .b(n_14291), .o(n_14564) );
no02f02 g53026_u0 ( .a(n_13756), .b(FE_OFN1705_n_4868), .o(g53026_p) );
in01f02 g53026_u1 ( .a(g53026_p), .o(n_14331) );
no02f02 g53028_u0 ( .a(n_14285), .b(n_14469), .o(n_14563) );
no02f02 g53029_u0 ( .a(n_14284), .b(n_14467), .o(n_16611) );
no02f02 g53031_u0 ( .a(n_13771), .b(FE_OFN1710_n_4868), .o(g53031_p) );
in01f02 g53031_u1 ( .a(g53031_p), .o(n_14329) );
no02f02 g53033_u0 ( .a(n_14462), .b(n_14277), .o(n_14560) );
no02f02 g53034_u0 ( .a(n_14274), .b(n_14461), .o(n_14559) );
no02f02 g53035_u0 ( .a(n_13770), .b(FE_OFN1705_n_4868), .o(g53035_p) );
in01f02 g53035_u1 ( .a(g53035_p), .o(n_14327) );
no02f02 g53036_u0 ( .a(n_14458), .b(n_14459), .o(n_14558) );
no02f02 g53037_u0 ( .a(n_14270), .b(n_14457), .o(n_14557) );
no02f02 g53039_u0 ( .a(n_13755), .b(FE_OFN1705_n_4868), .o(g53039_p) );
in01f02 g53039_u1 ( .a(g53039_p), .o(n_14325) );
no02f02 g53041_u0 ( .a(n_14451), .b(n_14264), .o(n_14554) );
no02f02 g53042_u0 ( .a(n_14449), .b(n_14448), .o(n_16623) );
no02f02 g53044_u0 ( .a(n_14447), .b(n_14260), .o(n_16625) );
no02f02 g53045_u0 ( .a(n_14445), .b(n_14444), .o(n_14551) );
no02f02 g53046_u0 ( .a(n_14256), .b(n_14443), .o(n_14550) );
no02f02 g53047_u0 ( .a(n_14254), .b(n_14441), .o(n_14549) );
no02f02 g53048_u0 ( .a(n_14439), .b(n_14252), .o(n_14548) );
no02f02 g53049_u0 ( .a(n_14436), .b(n_14437), .o(n_14547) );
no02f02 g53051_u0 ( .a(n_14432), .b(n_14514), .o(n_14545) );
no02f02 g53052_u0 ( .a(n_14430), .b(n_14512), .o(n_14544) );
no02f02 g53053_u0 ( .a(n_14510), .b(n_14428), .o(n_14543) );
no02f02 g53056_u0 ( .a(n_14508), .b(n_14422), .o(n_14541) );
no02f02 g53060_u0 ( .a(n_14415), .b(n_14416), .o(n_14521) );
no02f02 g53061_u0 ( .a(n_14414), .b(n_14504), .o(n_16615) );
no02f02 g53063_u0 ( .a(n_14500), .b(n_14410), .o(n_14536) );
no02f02 g53064_u0 ( .a(n_14498), .b(n_14408), .o(n_14535) );
no02f02 g53066_u0 ( .a(n_14495), .b(n_14403), .o(n_14534) );
no02f02 g53067_u0 ( .a(n_14493), .b(n_14401), .o(n_16617) );
no02f02 g53068_u0 ( .a(n_13767), .b(n_13332), .o(n_14386) );
no02f02 g53069_u0 ( .a(n_2446), .b(n_8524), .o(g53069_p) );
in01f02 g53069_u1 ( .a(g53069_p), .o(n_8595) );
na02m20 TIMEBOOST_cell_42875 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_141), .o(TIMEBOOST_net_12332) );
no02f02 g53071_u0 ( .a(n_14303), .b(n_14518), .o(g53071_p) );
in01f02 g53071_u1 ( .a(g53071_p), .o(n_14902) );
no02f02 g53072_u0 ( .a(n_14307), .b(n_14518), .o(g53072_p) );
in01f02 g53072_u1 ( .a(g53072_p), .o(n_14517) );
no02f02 g53073_u0 ( .a(n_13764), .b(FE_OFN1708_n_4868), .o(g53073_p) );
in01f02 g53073_u1 ( .a(g53073_p), .o(n_14315) );
no02f02 g53074_u0 ( .a(n_13761), .b(FE_OFN1708_n_4868), .o(g53074_p) );
in01f02 g53074_u1 ( .a(g53074_p), .o(n_14313) );
no02f04 g53075_u0 ( .a(n_13760), .b(FE_OFN1707_n_4868), .o(g53075_p) );
in01f02 g53075_u1 ( .a(g53075_p), .o(n_14311) );
no02f02 g53076_u0 ( .a(n_13759), .b(FE_OFN1706_n_4868), .o(g53076_p) );
in01f02 g53076_u1 ( .a(g53076_p), .o(n_14309) );
na02m02 TIMEBOOST_cell_69123 ( .a(TIMEBOOST_net_21769), .b(g65067_sb), .o(TIMEBOOST_net_12559) );
in01f02 g53077_u1 ( .a(g53077_p), .o(n_14317) );
in01s01 TIMEBOOST_cell_73963 ( .a(TIMEBOOST_net_23527), .o(TIMEBOOST_net_23528) );
in01f02 g53078_u1 ( .a(g53078_p), .o(n_14357) );
no02f02 g53079_u0 ( .a(n_13785), .b(FE_OFN1706_n_4868), .o(g53079_p) );
in01f02 g53079_u1 ( .a(g53079_p), .o(n_14355) );
no02f02 g53080_u0 ( .a(n_13783), .b(FE_OFN1706_n_4868), .o(g53080_p) );
in01f02 g53080_u1 ( .a(g53080_p), .o(n_14353) );
no02f02 g53082_u0 ( .a(n_13780), .b(FE_OFN1706_n_4868), .o(g53082_p) );
in01f02 g53082_u1 ( .a(g53082_p), .o(n_14349) );
no02f02 g53083_u0 ( .a(n_13729), .b(FE_OFN1706_n_4868), .o(g53083_p) );
in01f02 g53083_u1 ( .a(g53083_p), .o(n_14083) );
in01f02 g53084_u1 ( .a(g53084_p), .o(n_14347) );
na02f02 g53085_u0 ( .a(n_13829), .b(n_7658), .o(n_13831) );
na02f02 g53086_u0 ( .a(n_14076), .b(n_7657), .o(n_14078) );
no02f02 g53087_u0 ( .a(FE_OFN1708_n_4868), .b(n_13768), .o(g53087_p) );
in01f02 g53087_u1 ( .a(g53087_p), .o(n_14321) );
na02f02 g53088_u0 ( .a(n_13753), .b(n_1112), .o(n_14392) );
na02f02 g53089_u0 ( .a(n_13752), .b(n_1108), .o(n_14390) );
na02f02 g53090_u0 ( .a(n_13750), .b(n_1202), .o(n_14387) );
na02f02 g53091_u0 ( .a(n_13907), .b(n_7523), .o(n_13911) );
na02f02 g53092_u0 ( .a(n_13829), .b(n_7642), .o(n_13830) );
na02f02 g53093_u0 ( .a(n_14076), .b(n_7527), .o(n_14077) );
ao12f02 g53094_u0 ( .a(n_1551), .b(n_13749), .c(FE_OCPN1836_n_16798), .o(n_13910) );
na02m02 TIMEBOOST_cell_68733 ( .a(TIMEBOOST_net_21574), .b(TIMEBOOST_net_14319), .o(TIMEBOOST_net_17141) );
no02f01 g53096_u0 ( .a(n_4796), .b(n_14484), .o(n_14483) );
na02f02 g53097_u0 ( .a(n_13907), .b(n_7635), .o(n_13908) );
no02m02 g53098_u0 ( .a(n_13765), .b(FE_OFN1708_n_4868), .o(g53098_p) );
in01f02 g53098_u1 ( .a(g53098_p), .o(n_14319) );
ao12f02 g53099_u0 ( .a(n_1551), .b(n_2619), .c(n_13819), .o(n_14075) );
ao12f02 g53102_u0 ( .a(n_13592), .b(n_13671), .c(n_13784), .o(n_13785) );
ao12f02 g53103_u0 ( .a(n_13591), .b(n_13670), .c(n_13781), .o(n_13783) );
na03f02 TIMEBOOST_cell_73448 ( .a(TIMEBOOST_net_17047), .b(FE_OFN1258_n_4143), .c(g62888_sb), .o(n_6101) );
na02m08 TIMEBOOST_cell_52747 ( .a(pci_target_unit_pcit_if_strd_addr_in_693), .b(n_2507), .o(TIMEBOOST_net_16591) );
ao12f02 g53106_u0 ( .a(n_13587), .b(n_13668), .c(n_13784), .o(n_13780) );
ao12f02 g53107_u0 ( .a(n_13585), .b(n_13562), .c(n_13784), .o(n_13729) );
ao12f02 g53111_u0 ( .a(n_13581), .b(n_13664), .c(FE_OFN1946_n_13784), .o(n_13776) );
ao12f02 g53112_u0 ( .a(n_13579), .b(n_13663), .c(n_13781), .o(n_13775) );
ao12f02 g53113_u0 ( .a(n_13578), .b(n_13662), .c(FE_OFN969_n_13784), .o(n_13774) );
ao12f02 g53115_u0 ( .a(n_13576), .b(n_13560), .c(n_13763), .o(n_13728) );
ao12f02 g53116_u0 ( .a(n_13575), .b(n_13659), .c(FE_OFN1946_n_13784), .o(n_13772) );
ao12f02 g53117_u0 ( .a(n_13574), .b(n_13658), .c(FE_OFN1946_n_13784), .o(n_13771) );
ao12f02 g53118_u0 ( .a(n_13573), .b(n_13657), .c(n_13784), .o(n_13770) );
ao12f02 g53121_u0 ( .a(n_16331), .b(n_13810), .c(n_7310), .o(n_14074) );
na02f02 g53122_u0 ( .a(n_13716), .b(n_13766), .o(n_13767) );
na02f02 g53123_u0 ( .a(n_13716), .b(n_13333), .o(n_13918) );
na02f02 g53124_u0 ( .a(n_13716), .b(n_7396), .o(n_13917) );
no02f02 g53125_u0 ( .a(n_1100), .b(n_13748), .o(n_13828) );
no02s01 g53126_u0 ( .a(n_14305), .b(wbm_cti_o_1_), .o(n_14307) );
ao12f02 g53127_u0 ( .a(n_13569), .b(n_13653), .c(n_13784), .o(n_13765) );
no02f04 g53129_u0 ( .a(n_13844), .b(n_15371), .o(n_14484) );
ao12f02 g53133_u0 ( .a(n_13678), .b(n_13673), .c(n_13784), .o(n_13759) );
ao12f02 g53134_u0 ( .a(n_13680), .b(n_13754), .c(n_13561), .o(n_13829) );
ao12f02 g53135_u0 ( .a(n_13582), .b(n_13754), .c(n_13704), .o(n_14076) );
in01f01 g53136_u0 ( .a(n_13757), .o(n_13758) );
no02f02 g53137_u0 ( .a(n_13715), .b(n_7397), .o(n_13757) );
ao12f02 g53138_u0 ( .a(n_13722), .b(n_13334), .c(n_13721), .o(n_13756) );
ao12f02 g53139_u0 ( .a(FE_OFN1335_n_13720), .b(n_13414), .c(n_13721), .o(n_13755) );
ao12f02 g53140_u0 ( .a(n_1522), .b(n_7043), .c(n_7726), .o(n_8524) );
no02f02 g53141_u0 ( .a(n_13412), .b(n_14305), .o(g53141_p) );
in01f02 g53141_u1 ( .a(g53141_p), .o(n_14306) );
no02f02 g53142_u0 ( .a(n_13411), .b(n_14305), .o(g53142_p) );
in01f02 g53142_u1 ( .a(g53142_p), .o(n_14304) );
na02f01 TIMEBOOST_cell_26103 ( .a(pci_target_unit_pcit_if_strd_addr_in_704), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7156) );
oa12f02 g53145_u0 ( .a(n_6941), .b(n_13691), .c(n_13825), .o(n_13827) );
oa12f02 g53146_u0 ( .a(n_6940), .b(n_13689), .c(n_13825), .o(n_13826) );
oa12f02 g53147_u0 ( .a(n_6942), .b(n_13692), .c(n_13825), .o(n_13824) );
oa12f02 g53148_u0 ( .a(n_14305), .b(n_14965), .c(n_3164), .o(n_14303) );
in01f02 g53149_u0 ( .a(n_14890), .o(n_14482) );
ao12f04 g53150_u0 ( .a(n_14305), .b(n_824), .c(wbm_cyc_o_1378), .o(n_14890) );
na04f04 TIMEBOOST_cell_24238 ( .a(n_9021), .b(g57474_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q), .d(FE_OFN1396_n_8567), .o(n_10340) );
in01f02 g53154_u1 ( .a(g53154_p), .o(n_14301) );
na02f10 TIMEBOOST_cell_62880 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_783), .o(TIMEBOOST_net_20387) );
in01f02 g53155_u1 ( .a(g53155_p), .o(n_14480) );
na03f02 TIMEBOOST_cell_73532 ( .a(TIMEBOOST_net_17565), .b(FE_OFN2063_n_6391), .c(g62431_sb), .o(n_6735) );
na02m02 g58284_u1 ( .a(g58284_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q), .o(g58284_da) );
na03f02 TIMEBOOST_cell_34982 ( .a(TIMEBOOST_net_9386), .b(FE_OFN1377_n_8567), .c(g57554_sb), .o(n_10302) );
in01f02 g53158_u1 ( .a(g53158_p), .o(n_16595) );
na03f02 TIMEBOOST_cell_73810 ( .a(TIMEBOOST_net_16548), .b(FE_OFN1775_n_13800), .c(FE_OFN1769_n_14054), .o(g53259_p) );
in01f02 g53159_u1 ( .a(g53159_p), .o(n_14478) );
na04s02 TIMEBOOST_cell_73083 ( .a(TIMEBOOST_net_10780), .b(g65826_sb), .c(g61891_sb), .d(g61891_db), .o(n_8047) );
na02s02 TIMEBOOST_cell_69747 ( .a(TIMEBOOST_net_22081), .b(FE_OFN1634_n_9531), .o(TIMEBOOST_net_16364) );
na02f01 TIMEBOOST_cell_71636 ( .a(FE_OFN1762_n_10780), .b(TIMEBOOST_net_13513), .o(TIMEBOOST_net_23026) );
in01f02 g53163_u1 ( .a(g53163_p), .o(n_14296) );
na03f02 TIMEBOOST_cell_73348 ( .a(n_4521), .b(g62820_sb), .c(TIMEBOOST_net_5739), .o(n_6115) );
na02m10 TIMEBOOST_cell_52671 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q), .o(TIMEBOOST_net_16553) );
na04f04 TIMEBOOST_cell_24328 ( .a(n_8559), .b(g58589_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q), .d(FE_OFN1403_n_8567), .o(n_8912) );
in01f02 g53167_u1 ( .a(g53167_p), .o(n_14475) );
na02s01 TIMEBOOST_cell_52377 ( .a(configuration_wb_err_data_574), .b(parchk_pci_ad_out_in_1171), .o(TIMEBOOST_net_16406) );
in01f02 g53170_u1 ( .a(g53170_p), .o(n_14292) );
in01f02 g53171_u1 ( .a(g53171_p), .o(n_14473) );
na02f02 TIMEBOOST_cell_51515 ( .a(n_16852), .b(n_3049), .o(TIMEBOOST_net_15975) );
na02s01 TIMEBOOST_cell_63226 ( .a(FE_OFN596_n_9694), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q), .o(TIMEBOOST_net_20560) );
in01f02 g53174_u1 ( .a(g53174_p), .o(n_14290) );
na04f04 TIMEBOOST_cell_24332 ( .a(n_9667), .b(g57264_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q), .d(FE_OFN1384_n_8567), .o(n_11489) );
in01f02 g53175_u1 ( .a(g53175_p), .o(n_14471) );
na04m02 TIMEBOOST_cell_67287 ( .a(n_3741), .b(g64888_sb), .c(g64888_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q), .o(TIMEBOOST_net_17002) );
in01f02 g53182_u1 ( .a(g53182_p), .o(n_14286) );
na02f01 TIMEBOOST_cell_70358 ( .a(TIMEBOOST_net_17293), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_22387) );
in01f02 g53183_u1 ( .a(g53183_p), .o(n_14468) );
na03f04 TIMEBOOST_cell_73492 ( .a(n_3290), .b(pciu_bar0_in_377), .c(n_3058), .o(TIMEBOOST_net_10014) );
na03m02 TIMEBOOST_cell_72379 ( .a(n_188), .b(n_5757), .c(n_3395), .o(TIMEBOOST_net_22037) );
in01f02 g53187_u1 ( .a(g53187_p), .o(n_16610) );
na04f04 TIMEBOOST_cell_24244 ( .a(n_9557), .b(g57378_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q), .d(FE_OFN1384_n_8567), .o(n_11370) );
na02m01 TIMEBOOST_cell_43675 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_124), .o(TIMEBOOST_net_12732) );
na03f02 TIMEBOOST_cell_66655 ( .a(TIMEBOOST_net_17410), .b(FE_OFN1270_n_4095), .c(g62965_sb), .o(n_5952) );
in01f02 g53199_u1 ( .a(g53199_p), .o(n_14275) );
na03f02 TIMEBOOST_cell_66852 ( .a(TIMEBOOST_net_20668), .b(n_14971), .c(g58652_sb), .o(n_9237) );
in01f02 g53203_u1 ( .a(g53203_p), .o(n_14460) );
na03m02 TIMEBOOST_cell_66851 ( .a(n_3226), .b(g60692_sb), .c(TIMEBOOST_net_5500), .o(n_7575) );
na02m02 TIMEBOOST_cell_53361 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_135), .o(TIMEBOOST_net_16898) );
in01f02 g53206_u1 ( .a(g53206_p), .o(n_14272) );
na03f10 TIMEBOOST_cell_34718 ( .a(FE_RN_500_0), .b(n_7712), .c(n_16167), .o(n_16299) );
in01f02 g53207_u1 ( .a(g53207_p), .o(n_14271) );
na03f02 TIMEBOOST_cell_73588 ( .a(TIMEBOOST_net_17317), .b(FE_OFN1116_g64577_p), .c(g63140_sb), .o(n_4968) );
na04m01 TIMEBOOST_cell_67130 ( .a(TIMEBOOST_net_14025), .b(g54205_sb), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_388), .d(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q), .o(TIMEBOOST_net_16799) );
na03f02 TIMEBOOST_cell_64635 ( .a(TIMEBOOST_net_14140), .b(g64169_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q), .o(TIMEBOOST_net_13059) );
in01f02 g53210_u1 ( .a(g53210_p), .o(n_14456) );
na02m01 TIMEBOOST_cell_42863 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_126), .o(TIMEBOOST_net_12326) );
in01f02 g53211_u1 ( .a(g53211_p), .o(n_14269) );
na04f04 TIMEBOOST_cell_24342 ( .a(n_9842), .b(g57085_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q), .d(FE_OFN1422_n_8567), .o(n_11657) );
in01f02 g53214_u1 ( .a(g53214_p), .o(n_14454) );
na04f10 TIMEBOOST_cell_47218 ( .a(FE_OCP_RBN2224_n_16322), .b(n_440), .c(n_46), .d(n_16322), .o(n_16547) );
na04f04 TIMEBOOST_cell_24248 ( .a(n_9554), .b(g57373_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q), .d(FE_OFN1419_n_8567), .o(n_11375) );
na04f04 TIMEBOOST_cell_24344 ( .a(n_9123), .b(g57083_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q), .d(FE_OFN1404_n_8567), .o(n_10493) );
na02s01 TIMEBOOST_cell_45821 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q), .o(TIMEBOOST_net_13805) );
na02f02 TIMEBOOST_cell_26341 ( .a(n_7622), .b(n_7725), .o(TIMEBOOST_net_7275) );
in01f02 g53226_u1 ( .a(g53226_p), .o(n_16622) );
na04f04 TIMEBOOST_cell_24348 ( .a(n_9854), .b(g57077_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q), .d(FE_OFN1408_n_8567), .o(n_11666) );
na02f08 TIMEBOOST_cell_25747 ( .a(n_3222), .b(n_2447), .o(TIMEBOOST_net_6978) );
in01f02 g53230_u1 ( .a(g53230_p), .o(n_16624) );
in01f02 g53231_u1 ( .a(g53231_p), .o(n_14446) );
na04f04 TIMEBOOST_cell_24350 ( .a(n_9859), .b(g57073_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q), .d(FE_OFN1415_n_8567), .o(n_11669) );
na03s01 TIMEBOOST_cell_72413 ( .a(wbs_dat_i_28_), .b(g61885_sb), .c(TIMEBOOST_net_9647), .o(TIMEBOOST_net_12831) );
in01f02 g53234_u1 ( .a(g53234_p), .o(n_14258) );
na02m08 TIMEBOOST_cell_43577 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q), .b(pci_target_unit_fifos_pciw_cbe_in), .o(TIMEBOOST_net_12683) );
in01f02 g53235_u1 ( .a(g53235_p), .o(n_14257) );
na02m08 TIMEBOOST_cell_69234 ( .a(FE_OFN643_n_4677), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q), .o(TIMEBOOST_net_21825) );
in01f02 g53238_u1 ( .a(g53238_p), .o(n_14255) );
na02f02 TIMEBOOST_cell_50168 ( .a(TIMEBOOST_net_15301), .b(g60620_sb), .o(n_4834) );
in01f02 g53239_u1 ( .a(g53239_p), .o(n_14442) );
na02m02 TIMEBOOST_cell_69236 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q), .b(FE_OFN644_n_4677), .o(TIMEBOOST_net_21826) );
na03m06 TIMEBOOST_cell_64634 ( .a(n_3774), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q), .c(FE_OFN667_n_4495), .o(TIMEBOOST_net_10567) );
in01f02 g53242_u1 ( .a(g53242_p), .o(n_14440) );
in01f02 g53243_u1 ( .a(g53243_p), .o(n_14253) );
na04f04 TIMEBOOST_cell_24250 ( .a(n_9561), .b(g57371_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q), .d(FE_OFN1423_n_8567), .o(n_11379) );
na03f02 TIMEBOOST_cell_47228 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_13518), .c(FE_OFN1584_n_12306), .o(n_12522) );
na03f02 TIMEBOOST_cell_73744 ( .a(TIMEBOOST_net_13667), .b(FE_OFN1755_n_12681), .c(FE_OCP_RBN1974_n_12381), .o(n_12767) );
na04f04 TIMEBOOST_cell_24352 ( .a(n_9861), .b(g57071_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q), .d(FE_OFN1425_n_8567), .o(n_11670) );
na04f02 TIMEBOOST_cell_34720 ( .a(n_1039), .b(n_9144), .c(wishbone_slave_unit_fifos_inGreyCount_reg_1__Q), .d(g57908_sb), .o(n_8920) );
in01f02 g53250_u1 ( .a(g53250_p), .o(n_14250) );
in01f02 g53251_u1 ( .a(g53251_p), .o(n_14435) );
na04f04 TIMEBOOST_cell_24252 ( .a(n_9050), .b(g57366_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q), .d(FE_OFN1396_n_8567), .o(n_10384) );
na02m08 TIMEBOOST_cell_52871 ( .a(wbs_dat_i_27_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q), .o(TIMEBOOST_net_16653) );
in01f02 g53254_u1 ( .a(g53254_p), .o(n_14515) );
na04m08 TIMEBOOST_cell_72719 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q), .b(FE_OFN1626_n_4438), .c(g64855_sb), .d(n_3739), .o(n_3721) );
in01f02 g53255_u1 ( .a(g53255_p), .o(n_14433) );
na03f04 TIMEBOOST_cell_73349 ( .a(TIMEBOOST_net_16686), .b(g54319_sb), .c(TIMEBOOST_net_387), .o(TIMEBOOST_net_11863) );
na02m10 TIMEBOOST_cell_45631 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_13710) );
in01f02 g53258_u1 ( .a(g53258_p), .o(n_14431) );
na02f04 TIMEBOOST_cell_26339 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q), .b(n_504), .o(TIMEBOOST_net_7274) );
in01f02 g53259_u1 ( .a(g53259_p), .o(n_14513) );
na04f02 TIMEBOOST_cell_67945 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q), .b(FE_OFN1115_g64577_p), .c(n_3844), .d(g63128_sb), .o(n_4996) );
na02m08 TIMEBOOST_cell_62618 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q), .b(pci_target_unit_fifos_pciw_addr_data_in), .o(TIMEBOOST_net_20256) );
in01f02 g53262_u1 ( .a(g53262_p), .o(n_14511) );
in01f02 g53263_u1 ( .a(g53263_p), .o(n_14429) );
na02m04 TIMEBOOST_cell_53363 ( .a(TIMEBOOST_net_12411), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q), .o(TIMEBOOST_net_16899) );
ao22f02 g53265_u0 ( .a(n_13555), .b(n_13447), .c(FE_OFN1618_n_1787), .d(conf_wb_err_bc_in), .o(n_13753) );
na02f02 TIMEBOOST_cell_69395 ( .a(TIMEBOOST_net_21905), .b(g64945_sb), .o(TIMEBOOST_net_20638) );
na02s06 TIMEBOOST_cell_43465 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q), .o(TIMEBOOST_net_12627) );
in01f02 g53267_u1 ( .a(g53267_p), .o(n_14427) );
na02f06 TIMEBOOST_cell_26301 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(TIMEBOOST_net_7255) );
in01f02 g53268_u1 ( .a(g53268_p), .o(n_14426) );
na02s01 TIMEBOOST_cell_43455 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q), .o(TIMEBOOST_net_12622) );
na02s01 TIMEBOOST_cell_43453 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q), .o(TIMEBOOST_net_12621) );
na02s01 TIMEBOOST_cell_43451 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q), .o(TIMEBOOST_net_12620) );
in01f02 g53275_u1 ( .a(g53275_p), .o(n_14421) );
na03f01 TIMEBOOST_cell_73022 ( .a(TIMEBOOST_net_22012), .b(FE_OFN1033_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q), .o(TIMEBOOST_net_23284) );
in01f02 g53276_u1 ( .a(g53276_p), .o(n_14420) );
na02f02 TIMEBOOST_cell_68357 ( .a(TIMEBOOST_net_21386), .b(g64087_sb), .o(TIMEBOOST_net_13103) );
na02f01 TIMEBOOST_cell_62805 ( .a(TIMEBOOST_net_20349), .b(FE_OFN1055_n_4727), .o(TIMEBOOST_net_16345) );
ao22f02 g53281_u0 ( .a(n_13554), .b(n_13447), .c(FE_OFN1618_n_1787), .d(conf_wb_err_bc_in_847), .o(n_13752) );
na02s01 TIMEBOOST_cell_43449 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_12619) );
na02m02 TIMEBOOST_cell_68928 ( .a(n_4465), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_21672) );
na04f04 TIMEBOOST_cell_24366 ( .a(n_9887), .b(g57043_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q), .d(FE_OFN1389_n_8567), .o(n_11691) );
na02m10 TIMEBOOST_cell_50015 ( .a(wishbone_slave_unit_pcim_sm_data_in_642), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q), .o(TIMEBOOST_net_15225) );
in01f02 g53288_u1 ( .a(g53288_p), .o(n_14413) );
na02m10 TIMEBOOST_cell_26321 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q), .b(n_13447), .o(TIMEBOOST_net_7265) );
in01f02 g53289_u1 ( .a(g53289_p), .o(n_16614) );
ao22f02 g53290_u0 ( .a(n_13553), .b(n_13447), .c(FE_OFN1618_n_1787), .d(conf_wb_err_bc_in_848), .o(n_13750) );
na04f04 TIMEBOOST_cell_36110 ( .a(parchk_pci_ad_out_in_1185), .b(g62088_sb), .c(configuration_wb_err_data_588), .d(FE_OFN1173_n_5592), .o(n_5619) );
na04f04 TIMEBOOST_cell_36111 ( .a(parchk_pci_ad_out_in_1181), .b(g62084_sb), .c(configuration_wb_err_data_584), .d(FE_OFN1165_n_5615), .o(n_5625) );
na02s01 TIMEBOOST_cell_45633 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q), .o(TIMEBOOST_net_13711) );
in01f02 g53298_u1 ( .a(g53298_p), .o(n_14499) );
na04f04 TIMEBOOST_cell_36112 ( .a(parchk_pci_ad_out_in_1179), .b(g62082_sb), .c(configuration_wb_err_data_582), .d(FE_OFN1173_n_5592), .o(n_5627) );
na02s01 TIMEBOOST_cell_31421 ( .a(FE_OFN211_n_9858), .b(g57965_sb), .o(TIMEBOOST_net_9815) );
na03f02 TIMEBOOST_cell_34984 ( .a(TIMEBOOST_net_9387), .b(FE_OFN1414_n_8567), .c(g57087_sb), .o(n_11655) );
in01f02 g53301_u1 ( .a(g53301_p), .o(n_14407) );
na03s02 TIMEBOOST_cell_73655 ( .a(FE_OFN533_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q), .c(TIMEBOOST_net_22916), .o(TIMEBOOST_net_21029) );
in01f02 g53302_u1 ( .a(g53302_p), .o(n_14497) );
na02s01 TIMEBOOST_cell_31422 ( .a(TIMEBOOST_net_9815), .b(g57950_db), .o(n_9859) );
in01f02 g53310_u1 ( .a(g53310_p), .o(n_14494) );
na02s01 TIMEBOOST_cell_49273 ( .a(FE_OFN552_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q), .o(TIMEBOOST_net_14854) );
na02m02 TIMEBOOST_cell_69226 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q), .b(FE_OFN643_n_4677), .o(TIMEBOOST_net_21821) );
in01f02 g53314_u1 ( .a(g53314_p), .o(n_16616) );
na02f01 TIMEBOOST_cell_52279 ( .a(TIMEBOOST_net_12704), .b(FE_OFN1051_n_16657), .o(TIMEBOOST_net_16357) );
in01s01 TIMEBOOST_cell_73966 ( .a(wbm_dat_i_3_), .o(TIMEBOOST_net_23531) );
na02f02 TIMEBOOST_cell_50152 ( .a(TIMEBOOST_net_15293), .b(g60665_sb), .o(n_5654) );
na02f02 TIMEBOOST_cell_70519 ( .a(TIMEBOOST_net_22467), .b(g63065_sb), .o(n_5120) );
na03m02 TIMEBOOST_cell_49123 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN2256_n_8060), .c(n_1919), .o(TIMEBOOST_net_14779) );
na04f04 TIMEBOOST_cell_24581 ( .a(n_9588), .b(g57340_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q), .d(FE_OFN1428_n_8567), .o(n_11411) );
na02s02 TIMEBOOST_cell_43758 ( .a(TIMEBOOST_net_12773), .b(g58243_sb), .o(TIMEBOOST_net_9339) );
na02s01 TIMEBOOST_cell_71420 ( .a(FE_OFN219_n_9853), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q), .o(TIMEBOOST_net_22918) );
na02m04 TIMEBOOST_cell_70756 ( .a(wbm_adr_o_26_), .b(g58636_sb), .o(TIMEBOOST_net_22586) );
na02m01 TIMEBOOST_cell_48889 ( .a(n_3780), .b(FE_OFN1645_n_4671), .o(TIMEBOOST_net_14662) );
na03m06 TIMEBOOST_cell_72614 ( .a(TIMEBOOST_net_23155), .b(FE_OFN1013_n_4734), .c(g64186_sb), .o(n_4735) );
na02f01 g53399_u0 ( .a(n_13901), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q), .o(n_14957) );
na02f02 g53400_u0 ( .a(FE_OCP_RBN1984_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q), .o(n_14956) );
na02s01 TIMEBOOST_cell_43671 ( .a(pci_target_unit_del_sync_addr_in_227), .b(parchk_pci_ad_reg_in_1228), .o(TIMEBOOST_net_12730) );
na02m02 TIMEBOOST_cell_3237 ( .a(TIMEBOOST_net_178), .b(g60688_sb), .o(n_3880) );
na02m06 TIMEBOOST_cell_42947 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_125), .o(TIMEBOOST_net_12368) );
na04f04 TIMEBOOST_cell_24329 ( .a(n_9717), .b(g57217_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q), .d(FE_OFN1423_n_8567), .o(n_11540) );
na03f02 TIMEBOOST_cell_73001 ( .a(TIMEBOOST_net_5401), .b(n_3453), .c(n_3423), .o(n_5723) );
na02f02 TIMEBOOST_cell_54734 ( .a(TIMEBOOST_net_17584), .b(FE_RN_702_0), .o(FE_RN_703_0) );
in01s01 TIMEBOOST_cell_63541 ( .a(TIMEBOOST_net_20721), .o(TIMEBOOST_net_20720) );
na04f04 TIMEBOOST_cell_24511 ( .a(n_9702), .b(g57243_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q), .d(FE_OFN1423_n_8567), .o(n_11515) );
na02f02 TIMEBOOST_cell_70531 ( .a(TIMEBOOST_net_22473), .b(g63114_sb), .o(n_5027) );
na03m01 TIMEBOOST_cell_67894 ( .a(TIMEBOOST_net_12620), .b(FE_OFN1043_n_2037), .c(g65831_sb), .o(n_1886) );
na02s02 TIMEBOOST_cell_53560 ( .a(TIMEBOOST_net_16997), .b(g57917_sb), .o(TIMEBOOST_net_9323) );
na04f04 TIMEBOOST_cell_24583 ( .a(n_8547), .b(g58609_sb), .c(n_393), .d(FE_OFN2185_n_8567), .o(n_8898) );
in01m03 TIMEBOOST_cell_62385 ( .a(TIMEBOOST_net_20138), .o(TIMEBOOST_net_20137) );
na02s02 TIMEBOOST_cell_44150 ( .a(TIMEBOOST_net_12969), .b(g57915_sb), .o(n_9894) );
na02m02 TIMEBOOST_cell_31431 ( .a(n_4444), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_9820) );
na03f02 TIMEBOOST_cell_66193 ( .a(TIMEBOOST_net_20982), .b(FE_OFN1200_n_4090), .c(g62610_sb), .o(n_7375) );
na02f02 g53427_u0 ( .a(FE_OFN1771_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q), .o(n_14055) );
na02f02 g53428_u0 ( .a(FE_OFN1774_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q), .o(n_14226) );
na02f02 g53429_u0 ( .a(n_13891), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q), .o(n_14961) );
na02f02 g53430_u0 ( .a(FE_OCP_RBN1961_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q), .o(n_14960) );
na02s01 TIMEBOOST_cell_63253 ( .a(TIMEBOOST_net_20573), .b(TIMEBOOST_net_11116), .o(TIMEBOOST_net_9437) );
na04f04 TIMEBOOST_cell_24239 ( .a(n_9550), .b(g57384_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q), .d(FE_OFN1419_n_8567), .o(n_11361) );
na04f04 TIMEBOOST_cell_24585 ( .a(n_8552), .b(g58596_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q), .d(FE_OFN2185_n_8567), .o(n_9191) );
na02f02 g53435_u0 ( .a(n_13891), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q), .o(n_14963) );
na04f04 TIMEBOOST_cell_24337 ( .a(n_9837), .b(g57089_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q), .d(FE_OFN1419_n_8567), .o(n_11652) );
na02s02 TIMEBOOST_cell_49124 ( .a(TIMEBOOST_net_14779), .b(g61763_sb), .o(n_8285) );
na03f02 TIMEBOOST_cell_66853 ( .a(TIMEBOOST_net_17176), .b(n_14971), .c(g58601_sb), .o(n_9241) );
na02f08 TIMEBOOST_cell_63421 ( .a(TIMEBOOST_net_20657), .b(n_16325), .o(n_16331) );
na03f02 TIMEBOOST_cell_65956 ( .a(TIMEBOOST_net_16407), .b(FE_OFN1163_n_5615), .c(g62079_sb), .o(n_5631) );
na02f02 TIMEBOOST_cell_70567 ( .a(TIMEBOOST_net_22491), .b(g63098_sb), .o(n_5058) );
na02f02 TIMEBOOST_cell_37977 ( .a(TIMEBOOST_net_10600), .b(g64164_sb), .o(n_4001) );
na02f02 TIMEBOOST_cell_70359 ( .a(TIMEBOOST_net_22387), .b(g63593_sb), .o(n_7171) );
na04f04 TIMEBOOST_cell_24321 ( .a(n_9659), .b(g57275_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q), .d(FE_OFN1423_n_8567), .o(n_11479) );
na04f04 TIMEBOOST_cell_24517 ( .a(n_9709), .b(g57228_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q), .d(FE_OFN1385_n_8567), .o(n_11528) );
na04f04 TIMEBOOST_cell_24343 ( .a(n_9843), .b(g57084_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q), .d(FE_OFN1424_n_8567), .o(n_11659) );
na02s02 TIMEBOOST_cell_38793 ( .a(TIMEBOOST_net_11008), .b(g65892_sb), .o(n_2569) );
na04f04 TIMEBOOST_cell_24545 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q), .b(FE_OFN2190_n_8567), .c(n_9670), .d(g57260_sb), .o(n_11493) );
na03f02 TIMEBOOST_cell_34983 ( .a(TIMEBOOST_net_9423), .b(FE_OFN1382_n_8567), .c(g57101_sb), .o(n_11645) );
na02f02 TIMEBOOST_cell_69813 ( .a(TIMEBOOST_net_22114), .b(g64831_sb), .o(TIMEBOOST_net_12821) );
na04f04 TIMEBOOST_cell_24577 ( .a(n_9565), .b(g57364_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q), .d(FE_OFN2170_n_8567), .o(n_11383) );
na04f04 TIMEBOOST_cell_24345 ( .a(n_9847), .b(g57082_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q), .d(FE_OFN1406_n_8567), .o(n_11660) );
na03f08 TIMEBOOST_cell_63420 ( .a(FE_RN_705_0), .b(FE_RN_592_0), .c(n_16330), .o(TIMEBOOST_net_20657) );
na02m20 TIMEBOOST_cell_43575 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_132), .o(TIMEBOOST_net_12682) );
na03m02 TIMEBOOST_cell_71930 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q), .b(FE_OFN624_n_4409), .c(g65046_sb), .o(TIMEBOOST_net_23173) );
na02s01 TIMEBOOST_cell_52619 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_16527) );
na02f02 g55321_u0 ( .a(FE_OFN1551_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q), .o(n_12372) );
na04f04 TIMEBOOST_cell_24349 ( .a(n_9857), .b(g57075_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q), .d(FE_OFN1405_n_8567), .o(n_11668) );
na02m10 TIMEBOOST_cell_53195 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58), .b(pci_target_unit_pcit_if_strd_addr_in_694), .o(TIMEBOOST_net_16815) );
na04m20 TIMEBOOST_cell_73023 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q), .c(FE_OFN1037_n_4732), .d(g64318_sb), .o(n_3858) );
na02s02 TIMEBOOST_cell_47752 ( .a(TIMEBOOST_net_14093), .b(g65686_sb), .o(n_2209) );
na04f04 TIMEBOOST_cell_24547 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q), .b(FE_OFN2182_n_8567), .c(n_9012), .d(g57510_sb), .o(n_10323) );
na03f02 TIMEBOOST_cell_73041 ( .a(n_1867), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q), .c(FE_OFN710_n_8232), .o(TIMEBOOST_net_14808) );
na02f02 g53481_u0 ( .a(FE_OFN1773_n_13800), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q), .o(n_14197) );
na03f01 TIMEBOOST_cell_69064 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q), .b(n_3774), .c(FE_OFN662_n_4392), .o(TIMEBOOST_net_21740) );
na02m02 TIMEBOOST_cell_43681 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN615_n_4501), .o(TIMEBOOST_net_12735) );
na02s02 TIMEBOOST_cell_54545 ( .a(g58124_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q), .o(TIMEBOOST_net_17490) );
na02s01 TIMEBOOST_cell_43667 ( .a(pci_target_unit_del_sync_addr_in_228), .b(parchk_pci_ad_reg_in_1229), .o(TIMEBOOST_net_12728) );
na02m02 TIMEBOOST_cell_72029 ( .a(TIMEBOOST_net_23222), .b(g64948_sb), .o(TIMEBOOST_net_17576) );
na03m06 TIMEBOOST_cell_73024 ( .a(TIMEBOOST_net_23226), .b(FE_OFN1031_n_4732), .c(g64320_sb), .o(n_3856) );
na02m10 TIMEBOOST_cell_53055 ( .a(configuration_pci_err_data_512), .b(wbm_dat_o_11_), .o(TIMEBOOST_net_16745) );
na04f04 TIMEBOOST_cell_24521 ( .a(n_9085), .b(g57223_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q), .d(FE_OFN1407_n_8567), .o(n_10436) );
na03m02 TIMEBOOST_cell_73117 ( .a(g64245_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q), .c(TIMEBOOST_net_12840), .o(TIMEBOOST_net_13058) );
na04f02 TIMEBOOST_cell_67647 ( .a(n_4466), .b(FE_OFN1223_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q), .d(g62426_sb), .o(n_6745) );
na02s01 TIMEBOOST_cell_71302 ( .a(FE_OFN1668_n_9477), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q), .o(TIMEBOOST_net_22859) );
na03m04 TIMEBOOST_cell_72829 ( .a(g65413_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q), .c(TIMEBOOST_net_14441), .o(TIMEBOOST_net_17469) );
na04f04 TIMEBOOST_cell_24523 ( .a(n_9716), .b(g57218_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q), .d(FE_OFN1389_n_8567), .o(n_11538) );
na03s02 TIMEBOOST_cell_73589 ( .a(FE_OFN268_n_9880), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q), .c(g58260_db), .o(TIMEBOOST_net_20609) );
na02f02 TIMEBOOST_cell_70319 ( .a(TIMEBOOST_net_22367), .b(g54147_sb), .o(n_13662) );
na02s01 TIMEBOOST_cell_63252 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q), .b(g58359_sb), .o(TIMEBOOST_net_20573) );
na04f04 TIMEBOOST_cell_24291 ( .a(n_9617), .b(g57312_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q), .d(FE_OFN1415_n_8567), .o(n_11438) );
na02m01 TIMEBOOST_cell_48587 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q), .b(n_3792), .o(TIMEBOOST_net_14511) );
na03f02 TIMEBOOST_cell_64998 ( .a(TIMEBOOST_net_14349), .b(g64359_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_9128) );
na03f04 TIMEBOOST_cell_66433 ( .a(TIMEBOOST_net_16784), .b(FE_OFN1311_n_6624), .c(g62663_sb), .o(n_6213) );
na04f04 TIMEBOOST_cell_24575 ( .a(n_9613), .b(g57316_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q), .d(FE_OFN2188_n_8567), .o(n_11435) );
na02s01 TIMEBOOST_cell_45635 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q), .o(TIMEBOOST_net_13712) );
na02m02 TIMEBOOST_cell_70361 ( .a(TIMEBOOST_net_22388), .b(g63610_sb), .o(n_7149) );
na04f04 TIMEBOOST_cell_36116 ( .a(parchk_pci_ad_out_in_1188), .b(g62092_sb), .c(configuration_wb_err_data_591), .d(FE_OFN1173_n_5592), .o(n_5614) );
na02f02 TIMEBOOST_cell_50892 ( .a(TIMEBOOST_net_15663), .b(g62418_sb), .o(n_6761) );
na02f01 TIMEBOOST_cell_62639 ( .a(TIMEBOOST_net_20266), .b(FE_OFN930_n_4730), .o(TIMEBOOST_net_14493) );
na04f04 TIMEBOOST_cell_36118 ( .a(parchk_pci_ad_out_in_1187), .b(g62091_sb), .c(configuration_wb_err_data_590), .d(FE_OFN1164_n_5615), .o(n_5616) );
na02f02 TIMEBOOST_cell_50272 ( .a(TIMEBOOST_net_15353), .b(g62386_sb), .o(n_6828) );
na02s02 TIMEBOOST_cell_48514 ( .a(TIMEBOOST_net_14474), .b(TIMEBOOST_net_10380), .o(TIMEBOOST_net_9368) );
na02m10 TIMEBOOST_cell_45629 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_13709) );
na02s01 TIMEBOOST_cell_31449 ( .a(g58039_sb), .b(FE_OFN207_n_9865), .o(TIMEBOOST_net_9829) );
na02f02 g53525_u0 ( .a(n_13891), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q), .o(n_13868) );
na02f04 g53526_u0 ( .a(FE_OCP_RBN1961_FE_OFN1591_n_13741), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q), .o(n_14022) );
in01s01 TIMEBOOST_cell_63540 ( .a(TIMEBOOST_net_20720), .o(wbs_adr_i_20_) );
na02s01 TIMEBOOST_cell_31450 ( .a(TIMEBOOST_net_9829), .b(g58039_db), .o(n_9750) );
na04f04 TIMEBOOST_cell_24579 ( .a(n_9054), .b(g57345_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q), .d(FE_OFN2180_n_8567), .o(n_10390) );
na04f04 TIMEBOOST_cell_24369 ( .a(n_9816), .b(g57110_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q), .d(FE_OFN1405_n_8567), .o(n_11637) );
na04f04 TIMEBOOST_cell_24257 ( .a(n_9569), .b(g57360_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q), .d(FE_OFN1384_n_8567), .o(n_11386) );
na04m02 TIMEBOOST_cell_67606 ( .a(TIMEBOOST_net_20932), .b(FE_OFN1655_n_9502), .c(g58323_sb), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q), .o(TIMEBOOST_net_9448) );
na04f04 TIMEBOOST_cell_67591 ( .a(TIMEBOOST_net_10054), .b(g62136_sb), .c(FE_OFN1170_n_5592), .d(configuration_wb_err_addr_537), .o(n_5557) );
na02m02 TIMEBOOST_cell_68773 ( .a(TIMEBOOST_net_21594), .b(g65759_sb), .o(n_1920) );
na04f04 TIMEBOOST_cell_36113 ( .a(parchk_pci_ad_out_in_1177), .b(g62080_sb), .c(configuration_wb_err_data_580), .d(FE_OFN1169_n_5592), .o(n_5630) );
na03s02 TIMEBOOST_cell_72666 ( .a(TIMEBOOST_net_12437), .b(FE_OFN1016_n_2053), .c(g65881_sb), .o(n_1865) );
na02m02 TIMEBOOST_cell_63225 ( .a(TIMEBOOST_net_20559), .b(g58086_sb), .o(n_9710) );
na04f04 TIMEBOOST_cell_24263 ( .a(n_9576), .b(g57352_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q), .d(FE_OFN1376_n_8567), .o(n_11396) );
na04f04 TIMEBOOST_cell_72471 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q), .b(FE_OFN906_n_4736), .c(pci_target_unit_fifos_pciw_addr_data_in_128), .d(g64201_sb), .o(n_3968) );
in01s01 TIMEBOOST_cell_73834 ( .a(n_11856), .o(TIMEBOOST_net_23399) );
na02m02 TIMEBOOST_cell_69390 ( .a(n_4323), .b(FE_OFN646_n_4497), .o(TIMEBOOST_net_21903) );
na02m10 TIMEBOOST_cell_52951 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q), .b(wishbone_slave_unit_pcim_sm_data_in), .o(TIMEBOOST_net_16693) );
na02f02 g53547_u0 ( .a(n_13790), .b(n_168), .o(n_14305) );
na02f01 g53548_u0 ( .a(n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q), .o(n_14163) );
na02f06 TIMEBOOST_cell_25748 ( .a(TIMEBOOST_net_6978), .b(n_4743), .o(n_8521) );
na02s02 TIMEBOOST_cell_54196 ( .a(TIMEBOOST_net_17315), .b(g58119_sb), .o(TIMEBOOST_net_9369) );
na02s02 TIMEBOOST_cell_68419 ( .a(TIMEBOOST_net_21417), .b(FE_OFN952_n_2055), .o(TIMEBOOST_net_20824) );
na02s01 TIMEBOOST_cell_43662 ( .a(TIMEBOOST_net_12725), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_11013) );
na03m02 TIMEBOOST_cell_72646 ( .a(TIMEBOOST_net_21488), .b(g64913_sb), .c(TIMEBOOST_net_21674), .o(TIMEBOOST_net_20977) );
na02s01 TIMEBOOST_cell_47514 ( .a(TIMEBOOST_net_13974), .b(g67042_sb), .o(n_1272) );
na02f02 g53556_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q), .o(n_14011) );
na02f02 g53557_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q), .o(n_13862) );
na02m10 TIMEBOOST_cell_53197 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53), .b(pci_target_unit_pcit_if_strd_addr_in_689), .o(TIMEBOOST_net_16816) );
na03f02 TIMEBOOST_cell_69964 ( .a(TIMEBOOST_net_16317), .b(FE_OFN1033_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_22190) );
na03f08 TIMEBOOST_cell_65978 ( .a(TIMEBOOST_net_20457), .b(FE_OCPN1909_n_16497), .c(g54321_sb), .o(n_13286) );
na03m04 TIMEBOOST_cell_72630 ( .a(g64916_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q), .c(TIMEBOOST_net_14248), .o(TIMEBOOST_net_17078) );
na04s02 TIMEBOOST_cell_73084 ( .a(TIMEBOOST_net_10782), .b(g65830_sb), .c(g61895_sb), .d(g61895_db), .o(n_8036) );
na02m02 TIMEBOOST_cell_52245 ( .a(n_3792), .b(FE_OFN644_n_4677), .o(TIMEBOOST_net_16340) );
na02s01 TIMEBOOST_cell_62638 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_149), .o(TIMEBOOST_net_20266) );
na04f04 TIMEBOOST_cell_24573 ( .a(n_9215), .b(g57469_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q), .d(FE_OFN2177_n_8567), .o(n_10820) );
in01s01 TIMEBOOST_cell_73868 ( .a(n_7879), .o(TIMEBOOST_net_23433) );
na03m02 TIMEBOOST_cell_73178 ( .a(TIMEBOOST_net_22182), .b(g64316_sb), .c(FE_OFN1134_g64577_p), .o(TIMEBOOST_net_15158) );
na02s02 TIMEBOOST_cell_44446 ( .a(TIMEBOOST_net_13117), .b(g58377_db), .o(n_9452) );
na02f01 g53572_u0 ( .a(n_13987), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q), .o(n_14000) );
na02f02 g53573_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q), .o(n_13999) );
na03f02 TIMEBOOST_cell_66277 ( .a(pci_target_unit_wishbone_master_bc_register_reg_2__Q), .b(g60638_sb), .c(TIMEBOOST_net_7600), .o(n_5694) );
na02s01 TIMEBOOST_cell_52379 ( .a(parchk_pci_ad_out_in), .b(configuration_wb_err_data), .o(TIMEBOOST_net_16407) );
na04f04 TIMEBOOST_cell_24331 ( .a(n_9747), .b(g57176_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q), .d(FE_OFN1408_n_8567), .o(n_11579) );
na03f02 TIMEBOOST_cell_73350 ( .a(TIMEBOOST_net_22416), .b(n_3591), .c(g63434_sb), .o(n_4930) );
na02s02 TIMEBOOST_cell_71371 ( .a(TIMEBOOST_net_22893), .b(g58050_sb), .o(TIMEBOOST_net_16942) );
na02f01 TIMEBOOST_cell_72198 ( .a(TIMEBOOST_net_12849), .b(FE_OFN2127_n_16497), .o(TIMEBOOST_net_23307) );
na02f02 g53582_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q), .o(n_13991) );
na02f02 g53583_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q), .o(n_13990) );
na02s01 TIMEBOOST_cell_37038 ( .a(pci_ad_i_14_), .b(parchk_pci_ad_reg_in_1218), .o(TIMEBOOST_net_10131) );
na02s02 TIMEBOOST_cell_48604 ( .a(TIMEBOOST_net_14519), .b(TIMEBOOST_net_10407), .o(TIMEBOOST_net_9535) );
na02m10 TIMEBOOST_cell_45283 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q), .o(TIMEBOOST_net_13536) );
na02f02 g53588_u0 ( .a(n_13987), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q), .o(n_13982) );
na02m06 TIMEBOOST_cell_68546 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_145), .o(TIMEBOOST_net_21481) );
na02f04 g53590_u0 ( .a(FE_OFN1606_n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q), .o(n_14144) );
na02f02 g53591_u0 ( .a(FE_OFN1600_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q), .o(n_14142) );
na02f02 g53592_u0 ( .a(FE_OCP_RBN1998_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q), .o(n_13980) );
na02f02 g53593_u0 ( .a(FE_OFN1587_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q), .o(n_13859) );
na02f02 TIMEBOOST_cell_70363 ( .a(TIMEBOOST_net_22389), .b(g63591_sb), .o(n_7180) );
na03f02 TIMEBOOST_cell_47313 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_13597), .c(FE_OCP_RBN1979_n_10273), .o(n_12760) );
na03f02 TIMEBOOST_cell_66279 ( .a(wbm_adr_o_6_), .b(g60632_sb), .c(TIMEBOOST_net_11654), .o(n_5704) );
na02s01 TIMEBOOST_cell_62637 ( .a(TIMEBOOST_net_20265), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_12734) );
na02s01 TIMEBOOST_cell_43666 ( .a(TIMEBOOST_net_12727), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_11015) );
na04m02 TIMEBOOST_cell_72921 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(FE_OFN1041_n_2037), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q), .d(g65890_sb), .o(n_1859) );
na03m02 TIMEBOOST_cell_66281 ( .a(wbm_adr_o_26_), .b(g60623_sb), .c(TIMEBOOST_net_7599), .o(n_4831) );
na02s01 TIMEBOOST_cell_37312 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q), .b(pci_target_unit_fifos_pcir_data_in_173), .o(TIMEBOOST_net_10268) );
na02f02 TIMEBOOST_cell_44664 ( .a(TIMEBOOST_net_13226), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_11599) );
na02s02 TIMEBOOST_cell_38096 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q), .b(g65818_sb), .o(TIMEBOOST_net_10660) );
na03f02 TIMEBOOST_cell_73590 ( .a(TIMEBOOST_net_17545), .b(FE_OFN1235_n_6391), .c(g62432_sb), .o(n_6733) );
na02s02 TIMEBOOST_cell_48164 ( .a(TIMEBOOST_net_14299), .b(g58230_sb), .o(TIMEBOOST_net_10528) );
na04s03 TIMEBOOST_cell_67367 ( .a(g61740_sb), .b(g61740_db), .c(TIMEBOOST_net_14172), .d(g65770_db), .o(n_8337) );
na04f04 TIMEBOOST_cell_24335 ( .a(n_9460), .b(g57504_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q), .d(FE_OFN1417_n_8567), .o(n_11234) );
na02f02 g53610_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q), .o(n_13972) );
na02f02 g53611_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q), .o(n_13857) );
na04m06 TIMEBOOST_cell_73031 ( .a(FE_OFN1810_n_4454), .b(TIMEBOOST_net_14542), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q), .d(g65045_sb), .o(TIMEBOOST_net_17073) );
na02f02 TIMEBOOST_cell_71105 ( .a(TIMEBOOST_net_22760), .b(g62380_sb), .o(n_6842) );
na02s01 TIMEBOOST_cell_53033 ( .a(wbm_adr_o_12_), .b(configuration_pci_err_addr_482), .o(TIMEBOOST_net_16734) );
na02s02 TIMEBOOST_cell_43668 ( .a(TIMEBOOST_net_12728), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_11016) );
na02m02 TIMEBOOST_cell_68547 ( .a(TIMEBOOST_net_21481), .b(FE_OFN1012_n_4734), .o(TIMEBOOST_net_20323) );
na02s02 TIMEBOOST_cell_48740 ( .a(TIMEBOOST_net_14587), .b(TIMEBOOST_net_10423), .o(TIMEBOOST_net_9481) );
na02f04 g53623_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q), .o(n_13856) );
na03f02 TIMEBOOST_cell_66435 ( .a(g62758_sb), .b(FE_OFN1320_n_6436), .c(TIMEBOOST_net_16777), .o(n_6123) );
na03f10 TIMEBOOST_cell_72381 ( .a(pci_cbe_i_2_), .b(g67070_sb), .c(parchk_pci_cbe_en_in), .o(TIMEBOOST_net_23125) );
na04f02 TIMEBOOST_cell_36860 ( .a(TIMEBOOST_net_8577), .b(n_10256), .c(g52618_sb), .d(TIMEBOOST_net_745), .o(n_11852) );
na03f04 TIMEBOOST_cell_72368 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .c(TIMEBOOST_net_23120), .o(n_1643) );
na02s01 TIMEBOOST_cell_43809 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q), .o(TIMEBOOST_net_12799) );
na04f02 TIMEBOOST_cell_72665 ( .a(TIMEBOOST_net_21518), .b(FE_OFN930_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q), .d(g64285_sb), .o(TIMEBOOST_net_13041) );
na03f02 TIMEBOOST_cell_47223 ( .a(FE_OFN1584_n_12306), .b(TIMEBOOST_net_13514), .c(FE_OFN1761_n_10780), .o(n_16596) );
na02m01 TIMEBOOST_cell_68492 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q), .b(g65272_sb), .o(TIMEBOOST_net_21454) );
na02s02 TIMEBOOST_cell_43672 ( .a(TIMEBOOST_net_12730), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_11018) );
na02s01 TIMEBOOST_cell_43734 ( .a(TIMEBOOST_net_12761), .b(g57913_sb), .o(n_9897) );
na02m02 TIMEBOOST_cell_68352 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(g65792_sb), .o(TIMEBOOST_net_21384) );
na02s01 TIMEBOOST_cell_43674 ( .a(TIMEBOOST_net_12731), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_11019) );
na02f02 TIMEBOOST_cell_69967 ( .a(TIMEBOOST_net_22191), .b(g52638_sb), .o(n_14750) );
na02s01 TIMEBOOST_cell_43736 ( .a(TIMEBOOST_net_12762), .b(g58012_sb), .o(n_9781) );
na02f04 g53643_u0 ( .a(FE_OFN1587_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q), .o(n_13854) );
na04f02 TIMEBOOST_cell_34719 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .b(n_9144), .c(wishbone_slave_unit_fifos_inGreyCount_reg_2__Q), .d(g58489_sb), .o(n_8919) );
na02f01 g53648_u0 ( .a(n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q), .o(n_14111) );
na02s01 TIMEBOOST_cell_45637 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q), .o(TIMEBOOST_net_13713) );
na02m10 TIMEBOOST_cell_62608 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q), .o(TIMEBOOST_net_20251) );
na03f10 TIMEBOOST_cell_64319 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q), .b(n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_405), .o(TIMEBOOST_net_17282) );
na02m04 TIMEBOOST_cell_69454 ( .a(g64844_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q), .o(TIMEBOOST_net_21935) );
na03f02 TIMEBOOST_cell_66924 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_16004), .c(FE_OFN1513_n_14987), .o(n_12629) );
na02m10 TIMEBOOST_cell_52621 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q), .o(TIMEBOOST_net_16528) );
na02s01 TIMEBOOST_cell_25321 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_99), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6765) );
na04f02 TIMEBOOST_cell_34721 ( .a(n_2051), .b(n_9144), .c(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .d(g57875_sb), .o(n_8921) );
na03m02 TIMEBOOST_cell_73025 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(FE_OFN1032_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q), .o(TIMEBOOST_net_23310) );
na03f02 TIMEBOOST_cell_73564 ( .a(TIMEBOOST_net_17071), .b(FE_OFN2064_n_6391), .c(g63042_sb), .o(n_5858) );
na03f02 TIMEBOOST_cell_66945 ( .a(TIMEBOOST_net_13612), .b(FE_OFN1572_n_11027), .c(FE_OFN1751_n_12086), .o(n_12606) );
na02s01 TIMEBOOST_cell_43744 ( .a(TIMEBOOST_net_12766), .b(g58057_db), .o(n_9732) );
na04f04 TIMEBOOST_cell_24355 ( .a(n_9867), .b(g57068_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q), .d(FE_OFN1423_n_8567), .o(n_11674) );
na02f02 TIMEBOOST_cell_47681 ( .a(g56934_sb), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_14058) );
na03s02 TIMEBOOST_cell_73003 ( .a(TIMEBOOST_net_21662), .b(TIMEBOOST_net_12497), .c(FE_OFN699_n_7845), .o(TIMEBOOST_net_22238) );
na02f02 TIMEBOOST_cell_30825 ( .a(n_9458), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q), .o(TIMEBOOST_net_9517) );
na03s02 TIMEBOOST_cell_73493 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q), .b(FE_OFN233_n_9876), .c(FE_OFN572_n_9502), .o(TIMEBOOST_net_12804) );
na04f04 TIMEBOOST_cell_73680 ( .a(n_2824), .b(n_2614), .c(n_2823), .d(n_3044), .o(n_4683) );
na02f02 g53674_u0 ( .a(FE_OFN1605_n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q), .o(n_13938) );
na02f02 g53675_u0 ( .a(FE_OFN1601_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q), .o(n_13937) );
na04f04 TIMEBOOST_cell_34713 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q), .b(FE_OFN1349_n_8567), .c(n_9882), .d(g57047_sb), .o(n_11687) );
na02s01 TIMEBOOST_cell_62636 ( .a(FE_OFN1651_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q), .o(TIMEBOOST_net_20265) );
na04m04 TIMEBOOST_cell_72732 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q), .b(FE_OFN660_n_4392), .c(g64940_sb), .d(n_4465), .o(n_4382) );
na02f01 g53680_u0 ( .a(n_13997), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q), .o(n_17021) );
na04f80 TIMEBOOST_cell_72541 ( .a(g58776_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q), .c(n_8884), .d(wbu_addr_in_267), .o(n_9851) );
na03f02 TIMEBOOST_cell_24019 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q), .b(g59113_sb), .c(TIMEBOOST_net_5529), .o(n_8703) );
na04f04 TIMEBOOST_cell_24367 ( .a(n_9888), .b(g57042_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q), .d(FE_OFN1423_n_8567), .o(n_11692) );
na02s01 TIMEBOOST_cell_38917 ( .a(TIMEBOOST_net_11070), .b(g52476_da), .o(TIMEBOOST_net_10018) );
na02f02 g53687_u0 ( .a(FE_OFN1602_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q), .o(n_14099) );
na02f02 g53688_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q), .o(n_13930) );
na02f02 g53689_u0 ( .a(FE_OFN1587_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q), .o(n_13849) );
na02s01 TIMEBOOST_cell_48513 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q), .b(FE_OFN525_n_9899), .o(TIMEBOOST_net_14474) );
na02m04 TIMEBOOST_cell_69077 ( .a(TIMEBOOST_net_21746), .b(g65422_sb), .o(n_4225) );
na02s01 TIMEBOOST_cell_53995 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q), .o(TIMEBOOST_net_17215) );
na02f01 TIMEBOOST_cell_68847 ( .a(TIMEBOOST_net_21631), .b(n_4488), .o(n_4261) );
na02f10 TIMEBOOST_cell_48660 ( .a(n_15014), .b(TIMEBOOST_net_14547), .o(n_15446) );
na03f02 TIMEBOOST_cell_72677 ( .a(TIMEBOOST_net_16586), .b(FE_OFN784_n_2678), .c(g65224_sb), .o(n_2663) );
na04f04 TIMEBOOST_cell_47191 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_782), .c(FE_OFN2088_n_13124), .d(g54346_sb), .o(n_12966) );
na02m01 TIMEBOOST_cell_43746 ( .a(TIMEBOOST_net_12767), .b(g57935_db), .o(n_9874) );
na03f02 TIMEBOOST_cell_66576 ( .a(TIMEBOOST_net_17536), .b(FE_OFN1268_n_4095), .c(g62487_sb), .o(n_6613) );
na02f04 g53701_u0 ( .a(FE_OFN1586_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q), .o(n_13847) );
na02f01 TIMEBOOST_cell_39117 ( .a(TIMEBOOST_net_11170), .b(g63020_sb), .o(n_5207) );
na02f02 g53706_u0 ( .a(FE_OCP_RBN1997_n_13971), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q), .o(n_13923) );
na02f02 g53707_u0 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q), .o(n_13846) );
no02f02 g53708_u0 ( .a(n_13710), .b(n_2629), .o(n_13749) );
no02f02 g53709_u0 ( .a(n_16456), .b(n_13921), .o(g53709_p) );
in01f02 g53709_u1 ( .a(g53709_p), .o(n_13922) );
ao12f04 g53710_u0 ( .a(n_13721), .b(n_13450), .c(n_1789), .o(n_13725) );
ao12f02 g53711_u0 ( .a(n_13721), .b(n_13448), .c(n_1785), .o(n_13722) );
ao12f02 g53712_u0 ( .a(n_13721), .b(n_13444), .c(n_1788), .o(n_13720) );
ao12f02 g53714_u0 ( .a(n_15347), .b(n_4795), .c(n_13813), .o(n_13844) );
na02f02 g53715_u0 ( .a(n_13681), .b(n_2630), .o(n_13748) );
ao22f06 g53716_u0 ( .a(n_1645), .b(n_7567), .c(n_1523), .d(n_15371), .o(n_7568) );
in01f02 g53718_u0 ( .a(n_13821), .o(n_13843) );
na02f02 TIMEBOOST_cell_18228 ( .a(TIMEBOOST_net_5477), .b(n_4664), .o(n_6984) );
ao22f02 g53720_u0 ( .a(n_2629), .b(n_13817), .c(n_13679), .d(n_13820), .o(n_13819) );
in01f02 g53721_u0 ( .a(n_13842), .o(n_13920) );
ao22f02 g53722_u0 ( .a(n_13625), .b(n_13820), .c(n_12167), .d(n_13817), .o(n_13842) );
in01f04 g53723_u0 ( .a(n_13715), .o(n_13716) );
no02f04 g53726_u0 ( .a(n_7093), .b(n_13335), .o(g53726_p) );
ao12f04 g53726_u1 ( .a(g53726_p), .b(n_13335), .c(n_7093), .o(n_13715) );
ao22f02 g53727_u0 ( .a(n_7531), .b(n_13679), .c(n_2764), .d(FE_OCPN1836_n_16798), .o(n_13919) );
no02f02 g53729_u0 ( .a(n_13679), .b(n_2629), .o(g53729_p) );
in01f02 g53729_u1 ( .a(g53729_p), .o(n_13681) );
na03f02 TIMEBOOST_cell_66631 ( .a(TIMEBOOST_net_8539), .b(FE_OCPN1847_n_14981), .c(g59090_sb), .o(n_8716) );
no02f02 g53731_u0 ( .a(n_13355), .b(n_13784), .o(n_13592) );
no02f02 g53732_u0 ( .a(n_13353), .b(n_13784), .o(n_13591) );
no02f02 g53734_u0 ( .a(n_13350), .b(n_13784), .o(n_13587) );
no02f02 g53735_u0 ( .a(n_13349), .b(n_13784), .o(n_13585) );
na02s01 TIMEBOOST_cell_54059 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_150), .o(TIMEBOOST_net_17247) );
no02f02 g53738_u0 ( .a(n_13416), .b(FE_OFN1709_n_4868), .o(n_13680) );
no02f02 g53739_u0 ( .a(n_13342), .b(FE_OFN1709_n_4868), .o(n_13582) );
ao12f02 g53740_u0 ( .a(FE_OFN969_n_13784), .b(n_13292), .c(n_7551), .o(n_13581) );
ao12f02 g53741_u0 ( .a(FE_OFN969_n_13784), .b(n_13291), .c(n_7550), .o(n_13579) );
ao12f02 g53742_u0 ( .a(FE_OFN969_n_13784), .b(n_13290), .c(n_7548), .o(n_13578) );
ao12f02 g53744_u0 ( .a(FE_OFN969_n_13784), .b(n_13287), .c(n_7547), .o(n_13576) );
no02f02 g53745_u0 ( .a(n_13339), .b(FE_OFN1946_n_13784), .o(n_13575) );
no02f02 g53746_u0 ( .a(n_13338), .b(FE_OFN1946_n_13784), .o(n_13574) );
no02f02 g53747_u0 ( .a(n_13337), .b(n_13784), .o(n_13573) );
na02s01 TIMEBOOST_cell_42723 ( .a(pci_ad_i_0_), .b(parchk_pci_ad_reg_in), .o(TIMEBOOST_net_12256) );
in01f02 g53750_u0 ( .a(n_13710), .o(n_13711) );
na02f04 g53751_u0 ( .a(n_15611), .b(n_13679), .o(n_13710) );
na02f02 g53752_u0 ( .a(n_13814), .b(n_13813), .o(g53752_p) );
in01f02 g53752_u1 ( .a(g53752_p), .o(n_13921) );
na02m02 TIMEBOOST_cell_72011 ( .a(TIMEBOOST_net_23213), .b(TIMEBOOST_net_10702), .o(TIMEBOOST_net_17025) );
no02f02 g53754_u0 ( .a(n_13784), .b(n_13346), .o(n_13569) );
na03f02 TIMEBOOST_cell_34986 ( .a(TIMEBOOST_net_9392), .b(FE_OFN1412_n_8567), .c(g57538_sb), .o(n_10311) );
na03f02 TIMEBOOST_cell_72570 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .b(n_6986), .c(n_4662), .o(TIMEBOOST_net_22446) );
na03m02 TIMEBOOST_cell_68746 ( .a(FE_OFN661_n_4392), .b(g64928_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q), .o(TIMEBOOST_net_21581) );
no02f02 g53759_u0 ( .a(n_13417), .b(n_13784), .o(n_13678) );
ao12f02 g53760_u0 ( .a(n_13784), .b(n_13295), .c(n_7307), .o(n_13564) );
in01f06 g53762_u0 ( .a(n_13743), .o(n_13903) );
in01f04 g53764_u0 ( .a(n_13743), .o(n_13891) );
in01f02 g53765_u0 ( .a(n_13743), .o(n_13873) );
in01f02 g53769_u0 ( .a(n_13807), .o(n_13987) );
in01f08 g53772_u0 ( .a(n_13807), .o(n_13971) );
in01f02 g53773_u0 ( .a(n_13807), .o(n_13993) );
na02m01 TIMEBOOST_cell_26565 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q), .b(n_12595), .o(TIMEBOOST_net_7387) );
in01f04 g53787_u0 ( .a(n_13674), .o(n_13741) );
na02m01 TIMEBOOST_cell_71988 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q), .o(TIMEBOOST_net_23202) );
na02s01 TIMEBOOST_cell_68186 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q), .b(pci_target_unit_fifos_pcir_data_in_185), .o(TIMEBOOST_net_21301) );
ao12f02 g53817_u0 ( .a(n_3333), .b(n_13273), .c(n_13447), .o(n_13563) );
na02m02 TIMEBOOST_cell_49102 ( .a(TIMEBOOST_net_14768), .b(g61995_sb), .o(n_7905) );
na02f08 TIMEBOOST_cell_37339 ( .a(TIMEBOOST_net_10281), .b(n_2982), .o(n_2983) );
na02f02 TIMEBOOST_cell_70521 ( .a(TIMEBOOST_net_22468), .b(g62828_sb), .o(n_5320) );
na02f04 g53823_u0 ( .a(n_13361), .b(n_2108), .o(n_13561) );
na02f04 g53824_u0 ( .a(n_13495), .b(n_2106), .o(n_13704) );
na02m01 TIMEBOOST_cell_68513 ( .a(TIMEBOOST_net_21464), .b(g66401_db), .o(n_2540) );
na02m04 TIMEBOOST_cell_38612 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q), .b(g65357_sb), .o(TIMEBOOST_net_10918) );
na02f01 TIMEBOOST_cell_70688 ( .a(TIMEBOOST_net_13047), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_22552) );
na03f02 TIMEBOOST_cell_72716 ( .a(g64893_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q), .c(TIMEBOOST_net_16253), .o(TIMEBOOST_net_17151) );
in01f06 g53839_u0 ( .a(n_13703), .o(n_13997) );
in01f04 g53848_u0 ( .a(n_13701), .o(n_13995) );
in01f04 g53856_u0 ( .a(n_16206), .o(n_13736) );
na02s02 TIMEBOOST_cell_53068 ( .a(TIMEBOOST_net_16751), .b(g58283_db), .o(n_9519) );
na03f02 TIMEBOOST_cell_67994 ( .a(TIMEBOOST_net_17409), .b(FE_OFN1204_n_4090), .c(g62915_sb), .o(n_6049) );
na02m01 TIMEBOOST_cell_25284 ( .a(TIMEBOOST_net_6746), .b(n_574), .o(TIMEBOOST_net_538) );
na02f02 g53863_u0 ( .a(n_13441), .b(n_4692), .o(n_13654) );
na02s01 TIMEBOOST_cell_43446 ( .a(TIMEBOOST_net_12617), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_10780) );
na02s01 TIMEBOOST_cell_25286 ( .a(TIMEBOOST_net_6747), .b(n_574), .o(TIMEBOOST_net_539) );
na02s01 TIMEBOOST_cell_47907 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q), .o(TIMEBOOST_net_14171) );
na03m02 TIMEBOOST_cell_72040 ( .a(n_3752), .b(FE_OFN1642_n_4671), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q), .o(TIMEBOOST_net_23228) );
na02s01 TIMEBOOST_cell_25288 ( .a(TIMEBOOST_net_6748), .b(n_574), .o(TIMEBOOST_net_5357) );
oa12f02 g53870_u0 ( .a(n_13434), .b(n_4712), .c(FE_OFN2072_n_15978), .o(n_13648) );
oa12f02 g53871_u0 ( .a(n_13432), .b(n_4200), .c(FE_OFN2072_n_15978), .o(n_13647) );
oa12f02 g53872_u0 ( .a(n_13431), .b(n_4161), .c(FE_OFN1000_n_15978), .o(n_13646) );
oa12f02 g53873_u0 ( .a(n_13430), .b(n_3474), .c(FE_OFN2072_n_15978), .o(n_13645) );
oa12f02 g53874_u0 ( .a(n_13359), .b(n_4206), .c(FE_OFN1000_n_15978), .o(n_13559) );
oa12f02 g53875_u0 ( .a(n_13429), .b(n_4714), .c(FE_OFN2072_n_15978), .o(n_13643) );
oa12f02 g53876_u0 ( .a(n_13428), .b(n_4668), .c(FE_OFN1000_n_15978), .o(n_13642) );
oa12f02 g53877_u0 ( .a(n_13427), .b(n_4201), .c(FE_OFN1000_n_15978), .o(n_13641) );
oa12f02 g53878_u0 ( .a(n_13358), .b(n_4886), .c(FE_OFN1000_n_15978), .o(n_13558) );
oa12f02 g53879_u0 ( .a(n_13490), .b(n_5753), .c(FE_OFN2072_n_15978), .o(n_13695) );
oa12f02 g53880_u0 ( .a(n_13426), .b(n_4862), .c(FE_OFN1000_n_15978), .o(n_13640) );
oa12f02 g53881_u0 ( .a(n_13425), .b(n_4700), .c(FE_OFN2072_n_15978), .o(n_13638) );
oa12f02 g53882_u0 ( .a(n_13424), .b(n_7341), .c(FE_OFN1000_n_15978), .o(n_13636) );
oa12f02 g53883_u0 ( .a(n_13357), .b(n_7362), .c(FE_OFN1000_n_15978), .o(n_13557) );
oa12f02 g53884_u0 ( .a(n_13423), .b(n_5731), .c(FE_OFN1001_n_15978), .o(n_13635) );
oa12f02 g53885_u0 ( .a(n_13422), .b(n_4158), .c(FE_OFN1001_n_15978), .o(n_13634) );
oa12f02 g53886_u0 ( .a(n_13421), .b(n_3477), .c(FE_OFN1001_n_15978), .o(n_13632) );
oa12f02 g53887_u0 ( .a(n_13420), .b(n_3484), .c(FE_OFN1001_n_15978), .o(n_13631) );
oa12f02 g53888_u0 ( .a(n_13419), .b(n_4157), .c(FE_OFN1001_n_15978), .o(n_13629) );
oa12f02 g53889_u0 ( .a(n_13418), .b(n_3479), .c(FE_OFN1000_n_15978), .o(n_13628) );
na03f04 TIMEBOOST_cell_66808 ( .a(TIMEBOOST_net_16849), .b(FE_OFN1344_n_8567), .c(g57395_sb), .o(n_11347) );
na02s01 TIMEBOOST_cell_45589 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q), .o(TIMEBOOST_net_13689) );
na02s02 TIMEBOOST_cell_28238 ( .a(TIMEBOOST_net_8223), .b(g65734_sb), .o(n_1909) );
na02m04 g53891_u2 ( .a(n_13548), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(g53891_db) );
na02f04 g53891_u3 ( .a(g53891_da), .b(g53891_db), .o(n_13555) );
in01f08 g53892_u0 ( .a(n_692), .o(g53892_sb) );
na03m01 TIMEBOOST_cell_41946 ( .a(g58173_sb), .b(FE_OFN211_n_9858), .c(g58173_db), .o(n_9617) );
na02m06 g53893_u2 ( .a(n_13541), .b(n_692), .o(g53893_db) );
na02f04 g53893_u3 ( .a(g53893_da), .b(g53893_db), .o(n_13553) );
ao12f01 g53894_u0 ( .a(n_13494), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q), .c(n_1041), .o(n_13692) );
ao12f01 g53895_u0 ( .a(n_13493), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q), .c(n_1041), .o(n_13691) );
ao12f01 g53896_u0 ( .a(n_13491), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q), .c(n_1041), .o(n_13689) );
in01f04 g53897_u0 ( .a(FE_OFN2072_n_15978), .o(g53897_sb) );
na02f20 TIMEBOOST_cell_62878 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_781), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q), .o(TIMEBOOST_net_20386) );
na02m01 TIMEBOOST_cell_68676 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q), .b(FE_OFN661_n_4392), .o(TIMEBOOST_net_21546) );
in01f02 g53898_u0 ( .a(FE_OFN1330_n_13547), .o(g53898_sb) );
na02m02 TIMEBOOST_cell_69402 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q), .b(FE_OFN646_n_4497), .o(TIMEBOOST_net_21909) );
na02s01 TIMEBOOST_cell_52331 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q), .b(g58352_sb), .o(TIMEBOOST_net_16383) );
na03f02 TIMEBOOST_cell_73709 ( .a(TIMEBOOST_net_13536), .b(FE_OCPN1825_n_12030), .c(FE_OFN1565_n_12502), .o(n_12518) );
in01f02 g53899_u0 ( .a(FE_OFN1330_n_13547), .o(g53899_sb) );
na02s01 TIMEBOOST_cell_63057 ( .a(TIMEBOOST_net_20475), .b(TIMEBOOST_net_202), .o(TIMEBOOST_net_9329) );
na03m02 TIMEBOOST_cell_65893 ( .a(n_4598), .b(g61956_sb), .c(g61956_db), .o(n_6961) );
in01f02 g53900_u0 ( .a(FE_OFN1330_n_13547), .o(g53900_sb) );
na03m02 TIMEBOOST_cell_73204 ( .a(TIMEBOOST_net_7130), .b(g65874_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q), .o(TIMEBOOST_net_22324) );
na03f02 TIMEBOOST_cell_73533 ( .a(TIMEBOOST_net_17500), .b(FE_OFN1236_n_6391), .c(g63144_sb), .o(n_5852) );
na02s01 TIMEBOOST_cell_52332 ( .a(TIMEBOOST_net_16383), .b(g58352_db), .o(n_9469) );
in01f02 g53901_u0 ( .a(FE_OFN1333_n_13547), .o(g53901_sb) );
no02m06 TIMEBOOST_cell_27629 ( .a(FE_RN_396_0), .b(n_13784), .o(TIMEBOOST_net_7919) );
na03f02 TIMEBOOST_cell_68032 ( .a(TIMEBOOST_net_17580), .b(FE_OFN1212_n_4151), .c(g62659_sb), .o(n_6226) );
in01f01 g53902_u0 ( .a(FE_OFN1331_n_13547), .o(g53902_sb) );
na02s01 TIMEBOOST_cell_48862 ( .a(TIMEBOOST_net_14648), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_9471) );
na02f02 TIMEBOOST_cell_71066 ( .a(TIMEBOOST_net_20529), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_22741) );
na02s01 TIMEBOOST_cell_3906 ( .a(n_16818), .b(n_1323), .o(TIMEBOOST_net_513) );
in01f02 g53903_u0 ( .a(FE_OFN1326_n_13547), .o(g53903_sb) );
na03s02 TIMEBOOST_cell_70216 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q), .b(FE_OFN2257_n_8060), .c(n_4516), .o(TIMEBOOST_net_22316) );
na03f02 TIMEBOOST_cell_65930 ( .a(TIMEBOOST_net_16667), .b(FE_OFN1164_n_5615), .c(g62103_sb), .o(n_5598) );
in01f02 g53904_u0 ( .a(FE_OFN1330_n_13547), .o(g53904_sb) );
na03m02 TIMEBOOST_cell_72977 ( .a(TIMEBOOST_net_16610), .b(FE_OFN1056_n_4727), .c(g64342_sb), .o(TIMEBOOST_net_13056) );
na02s03 TIMEBOOST_cell_3910 ( .a(pci_target_unit_del_sync_comp_done_reg_main), .b(n_1816), .o(TIMEBOOST_net_515) );
in01f02 g53905_u0 ( .a(FE_OFN1332_n_13547), .o(g53905_sb) );
na02m06 TIMEBOOST_cell_3911 ( .a(TIMEBOOST_net_515), .b(n_1817), .o(n_2468) );
in01s01 TIMEBOOST_cell_45998 ( .a(TIMEBOOST_net_13959), .o(TIMEBOOST_net_13958) );
in01f01 g53906_u0 ( .a(FE_OFN1331_n_13547), .o(g53906_sb) );
na03f02 TIMEBOOST_cell_34796 ( .a(TIMEBOOST_net_9424), .b(FE_OFN1392_n_8567), .c(g57385_sb), .o(n_11359) );
in01s01 TIMEBOOST_cell_45999 ( .a(TIMEBOOST_net_13960), .o(TIMEBOOST_net_13899) );
na02s01 TIMEBOOST_cell_3914 ( .a(n_8486), .b(n_653), .o(TIMEBOOST_net_517) );
in01f02 g53907_u0 ( .a(FE_OFN1331_n_13547), .o(g53907_sb) );
na04f02 TIMEBOOST_cell_67947 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q), .b(FE_OFN1115_g64577_p), .c(n_3861), .d(g63107_sb), .o(n_5040) );
na02s01 TIMEBOOST_cell_3915 ( .a(TIMEBOOST_net_517), .b(n_177), .o(TIMEBOOST_net_392) );
na02s02 TIMEBOOST_cell_51913 ( .a(g58262_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q), .o(TIMEBOOST_net_16174) );
in01f02 g53908_u0 ( .a(FE_OFN1331_n_13547), .o(g53908_sb) );
na03s01 TIMEBOOST_cell_72454 ( .a(pci_target_unit_del_sync_addr_in_213), .b(FE_OFN2094_n_2520), .c(g66414_db), .o(n_2519) );
na02s02 TIMEBOOST_cell_51914 ( .a(TIMEBOOST_net_16174), .b(TIMEBOOST_net_10350), .o(TIMEBOOST_net_9386) );
in01f02 g53909_u0 ( .a(FE_OFN1326_n_13547), .o(g53909_sb) );
na02f02 TIMEBOOST_cell_71215 ( .a(TIMEBOOST_net_22815), .b(g62447_sb), .o(n_7385) );
na02f02 TIMEBOOST_cell_52306 ( .a(TIMEBOOST_net_16370), .b(g61784_sb), .o(n_8236) );
in01f02 g53910_u0 ( .a(FE_OFN1332_n_13547), .o(g53910_sb) );
na04f04 TIMEBOOST_cell_42461 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q), .b(n_13184), .c(FE_OFN1326_n_13547), .d(g53903_sb), .o(n_13538) );
na02s02 TIMEBOOST_cell_49410 ( .a(TIMEBOOST_net_14922), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_12970) );
na03f02 TIMEBOOST_cell_73351 ( .a(TIMEBOOST_net_22417), .b(n_3995), .c(g62822_sb), .o(n_5335) );
in01f02 g53911_u0 ( .a(FE_OFN1327_n_13547), .o(g53911_sb) );
na02m04 TIMEBOOST_cell_26219 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q), .b(g64239_sb), .o(TIMEBOOST_net_7214) );
na02m04 TIMEBOOST_cell_18214 ( .a(TIMEBOOST_net_5470), .b(n_14839), .o(g52400_db) );
in01f02 g53912_u0 ( .a(FE_OFN1333_n_13547), .o(g53912_sb) );
na03f02 TIMEBOOST_cell_41754 ( .a(TIMEBOOST_net_10569), .b(g64150_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_8336) );
na02m02 TIMEBOOST_cell_54730 ( .a(TIMEBOOST_net_17582), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_15439) );
in01f02 g53913_u0 ( .a(FE_OFN1331_n_13547), .o(g53913_sb) );
na02m08 TIMEBOOST_cell_52797 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_142), .o(TIMEBOOST_net_16616) );
in01f02 g53914_u0 ( .a(FE_OFN1330_n_13547), .o(g53914_sb) );
na02m02 TIMEBOOST_cell_71918 ( .a(FE_OFN1623_n_4438), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q), .o(TIMEBOOST_net_23167) );
na02f01 TIMEBOOST_cell_70248 ( .a(TIMEBOOST_net_17284), .b(FE_OFN1095_g64577_p), .o(TIMEBOOST_net_22332) );
in01f01 g53915_u0 ( .a(FE_OFN1331_n_13547), .o(g53915_sb) );
na03f02 TIMEBOOST_cell_73042 ( .a(n_3887), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q), .c(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_15188) );
na02s01 TIMEBOOST_cell_68515 ( .a(TIMEBOOST_net_21465), .b(g66400_db), .o(n_2542) );
na02m01 TIMEBOOST_cell_43039 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q), .b(pci_target_unit_fifos_pciw_cbe_in_152), .o(TIMEBOOST_net_12414) );
in01f02 g53916_u0 ( .a(FE_OFN1326_n_13547), .o(g53916_sb) );
na02m02 TIMEBOOST_cell_26229 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q), .b(g64310_sb), .o(TIMEBOOST_net_7219) );
na02s03 TIMEBOOST_cell_52673 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q), .o(TIMEBOOST_net_16554) );
in01f02 g53917_u0 ( .a(FE_OFN1327_n_13547), .o(g53917_sb) );
na03f02 TIMEBOOST_cell_73767 ( .a(TIMEBOOST_net_13709), .b(FE_OFN1774_n_13800), .c(FE_OFN1771_n_14054), .o(g74886_p) );
na03f01 TIMEBOOST_cell_65063 ( .a(n_3774), .b(FE_OFN686_n_4417), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q), .o(TIMEBOOST_net_16259) );
na02f02 TIMEBOOST_cell_44662 ( .a(TIMEBOOST_net_13225), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_11577) );
in01f02 g53918_u0 ( .a(FE_OFN1327_n_13547), .o(g53918_sb) );
na02s02 TIMEBOOST_cell_48790 ( .a(TIMEBOOST_net_14612), .b(TIMEBOOST_net_11294), .o(TIMEBOOST_net_9355) );
in01f02 g53919_u0 ( .a(FE_OFN1330_n_13547), .o(g53919_sb) );
na03f02 TIMEBOOST_cell_66169 ( .a(TIMEBOOST_net_15239), .b(FE_OFN1181_n_3476), .c(g60627_sb), .o(n_5710) );
na02f02 TIMEBOOST_cell_68211 ( .a(TIMEBOOST_net_21313), .b(n_973), .o(TIMEBOOST_net_20664) );
na02f01 TIMEBOOST_cell_3940 ( .a(n_7044), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(TIMEBOOST_net_530) );
in01f02 g53920_u0 ( .a(FE_OFN1332_n_13547), .o(g53920_sb) );
na02m04 TIMEBOOST_cell_72098 ( .a(TIMEBOOST_net_12923), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q), .o(TIMEBOOST_net_23257) );
na02f02 TIMEBOOST_cell_3941 ( .a(TIMEBOOST_net_530), .b(n_243), .o(TIMEBOOST_net_77) );
na02m02 TIMEBOOST_cell_43055 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q), .b(FE_OFN629_n_4454), .o(TIMEBOOST_net_12422) );
in01f01 g53921_u0 ( .a(FE_OFN1331_n_13547), .o(g53921_sb) );
na02m02 TIMEBOOST_cell_3943 ( .a(TIMEBOOST_net_531), .b(g67057_sb), .o(n_1677) );
in01f01 g53922_u0 ( .a(FE_OFN1331_n_13547), .o(g53922_sb) );
na03f04 TIMEBOOST_cell_73480 ( .a(wbm_adr_o_21_), .b(g59382_sb), .c(g52401_sb), .o(TIMEBOOST_net_16456) );
na02s01 TIMEBOOST_cell_45367 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q), .o(TIMEBOOST_net_13578) );
in01f02 g53923_u0 ( .a(FE_OFN1327_n_13547), .o(g53923_sb) );
na04m06 TIMEBOOST_cell_72994 ( .a(TIMEBOOST_net_16619), .b(FE_OFN1051_n_16657), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q), .d(g64195_sb), .o(TIMEBOOST_net_16975) );
na02m02 TIMEBOOST_cell_3948 ( .a(FE_OCPN1839_n_1238), .b(n_15856), .o(TIMEBOOST_net_534) );
in01f02 g53924_u0 ( .a(FE_OFN1326_n_13547), .o(g53924_sb) );
na03m02 TIMEBOOST_cell_73085 ( .a(g65359_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q), .c(TIMEBOOST_net_20366), .o(TIMEBOOST_net_17417) );
in01f02 g53925_u0 ( .a(FE_OFN1331_n_13547), .o(g53925_sb) );
na02f02 TIMEBOOST_cell_3951 ( .a(TIMEBOOST_net_535), .b(g67040_sb), .o(n_1641) );
na03f02 TIMEBOOST_cell_34991 ( .a(TIMEBOOST_net_10013), .b(g57200_sb), .c(FE_OFN2170_n_8567), .o(n_10834) );
in01f02 g53926_u0 ( .a(FE_OFN1327_n_13547), .o(g53926_sb) );
na03f02 TIMEBOOST_cell_65968 ( .a(n_4610), .b(g61840_sb), .c(g61840_db), .o(n_6971) );
na02f01 TIMEBOOST_cell_3953 ( .a(TIMEBOOST_net_536), .b(g67051_sb), .o(n_1497) );
na03f02 TIMEBOOST_cell_66636 ( .a(TIMEBOOST_net_17097), .b(FE_OFN1316_n_6624), .c(g62416_sb), .o(n_6766) );
in01f02 g53927_u0 ( .a(FE_OFN1327_n_13547), .o(g53927_sb) );
na03m02 TIMEBOOST_cell_72704 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q), .b(g64824_sb), .c(TIMEBOOST_net_14290), .o(TIMEBOOST_net_16775) );
na03m02 TIMEBOOST_cell_72727 ( .a(g65672_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q), .c(TIMEBOOST_net_14314), .o(TIMEBOOST_net_17032) );
na03f02 TIMEBOOST_cell_34988 ( .a(TIMEBOOST_net_9419), .b(FE_OFN1407_n_8567), .c(g57048_sb), .o(n_10511) );
in01f01 g53928_u0 ( .a(FE_OFN1331_n_13547), .o(g53928_sb) );
na04f04 TIMEBOOST_cell_65970 ( .a(wbm_adr_o_14_), .b(g52402_sb), .c(g58843_sb), .d(g52445_db), .o(TIMEBOOST_net_15708) );
na02f02 TIMEBOOST_cell_3957 ( .a(TIMEBOOST_net_538), .b(g67040_sb), .o(n_1501) );
in01f02 g53929_u0 ( .a(FE_OFN1333_n_13547), .o(g53929_sb) );
na02f01 TIMEBOOST_cell_3959 ( .a(TIMEBOOST_net_539), .b(g67040_sb), .o(n_1704) );
na02m10 TIMEBOOST_cell_52675 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_16555) );
in01f02 g53930_u0 ( .a(FE_OFN1327_n_13547), .o(g53930_sb) );
na02f02 TIMEBOOST_cell_70775 ( .a(TIMEBOOST_net_22595), .b(g59801_sb), .o(TIMEBOOST_net_20554) );
in01s01 TIMEBOOST_cell_67752 ( .a(TIMEBOOST_net_21178), .o(TIMEBOOST_net_21179) );
na03f02 TIMEBOOST_cell_34763 ( .a(TIMEBOOST_net_9359), .b(FE_OFN1401_n_8567), .c(g57431_sb), .o(n_11303) );
in01f01 g53931_u0 ( .a(FE_OFN1331_n_13547), .o(g53931_sb) );
na03f02 TIMEBOOST_cell_72957 ( .a(TIMEBOOST_net_21785), .b(g64275_sb), .c(FE_OFN2104_g64577_p), .o(TIMEBOOST_net_22545) );
na02s01 TIMEBOOST_cell_49529 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_14982) );
in01f02 g53932_u0 ( .a(FE_OFN1326_n_13547), .o(g53932_sb) );
na02s01 TIMEBOOST_cell_43663 ( .a(pci_target_unit_del_sync_addr_in_213), .b(parchk_pci_ad_reg_in_1214), .o(TIMEBOOST_net_12726) );
na02s01 TIMEBOOST_cell_3967 ( .a(TIMEBOOST_net_543), .b(n_14070), .o(TIMEBOOST_net_412) );
ao22f02 g53934_u0 ( .a(pci_target_unit_wishbone_master_retried), .b(wbm_cyc_o_1378), .c(wbm_ack_i), .d(wbm_stb_o), .o(n_13790) );
na02s01 TIMEBOOST_cell_3638 ( .a(n_2353), .b(n_8498), .o(TIMEBOOST_net_379) );
na02f02 g53935_u3 ( .a(g53935_da), .b(g53935_db), .o(n_13512) );
na02s01 TIMEBOOST_cell_39773 ( .a(TIMEBOOST_net_11498), .b(g58095_db), .o(n_9081) );
in01s01 TIMEBOOST_cell_73914 ( .a(n_2521), .o(TIMEBOOST_net_23479) );
in01f02 g53937_u0 ( .a(FE_OFN2072_n_15978), .o(g53937_sb) );
na02s01 TIMEBOOST_cell_4018 ( .a(parchk_pci_ad_reg_in_1220), .b(g65858_sb), .o(TIMEBOOST_net_569) );
na03f02 TIMEBOOST_cell_25000 ( .a(FE_RN_92_0), .b(n_10977), .c(n_12586), .o(n_12848) );
na02s02 TIMEBOOST_cell_25979 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q), .b(FE_OFN952_n_2055), .o(TIMEBOOST_net_7094) );
na02f02 TIMEBOOST_cell_3619 ( .a(TIMEBOOST_net_369), .b(n_7739), .o(n_14491) );
na02f02 TIMEBOOST_cell_70174 ( .a(TIMEBOOST_net_12927), .b(g64205_sb), .o(TIMEBOOST_net_22295) );
na02m10 TIMEBOOST_cell_3620 ( .a(n_2415), .b(n_1615), .o(TIMEBOOST_net_370) );
in01f06 g53939_u0 ( .a(FE_OFN1001_n_15978), .o(g53939_sb) );
na02s01 TIMEBOOST_cell_38218 ( .a(n_3030), .b(g65216_sb), .o(TIMEBOOST_net_10721) );
na02s03 TIMEBOOST_cell_68420 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q), .b(TIMEBOOST_net_13907), .o(TIMEBOOST_net_21418) );
in01f01 g53940_u0 ( .a(FE_OFN1001_n_15978), .o(g53940_sb) );
na02m08 TIMEBOOST_cell_52953 ( .a(wishbone_slave_unit_pcim_sm_data_in_654), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q), .o(TIMEBOOST_net_16694) );
na03f04 TIMEBOOST_cell_73481 ( .a(wbm_adr_o_24_), .b(g60681_sb), .c(g52398_sb), .o(TIMEBOOST_net_8552) );
na02s01 TIMEBOOST_cell_45369 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q), .o(TIMEBOOST_net_13579) );
na02f01 g62450_u2 ( .a(n_3791), .b(FE_OFN1222_n_6391), .o(g62450_db) );
na02m01 TIMEBOOST_cell_68906 ( .a(n_4465), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q), .o(TIMEBOOST_net_21661) );
na02s02 TIMEBOOST_cell_28173 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q), .b(g65867_sb), .o(TIMEBOOST_net_8191) );
in01s01 TIMEBOOST_cell_46000 ( .a(TIMEBOOST_net_13961), .o(TIMEBOOST_net_13960) );
na04m10 TIMEBOOST_cell_73004 ( .a(FE_OFN1046_n_16657), .b(TIMEBOOST_net_16615), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q), .d(g64108_sb), .o(TIMEBOOST_net_9916) );
na03f02 TIMEBOOST_cell_73768 ( .a(TIMEBOOST_net_13700), .b(FE_OFN1774_n_13800), .c(FE_OFN1770_n_14054), .o(g53171_p) );
na03f02 TIMEBOOST_cell_66228 ( .a(TIMEBOOST_net_13232), .b(FE_OFN1295_n_4098), .c(g62341_sb), .o(n_6917) );
no03f06 TIMEBOOST_cell_184 ( .a(n_15142), .b(g74749_p), .c(FE_RN_9_0), .o(n_15457) );
na03m02 TIMEBOOST_cell_72755 ( .a(n_4488), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q), .c(TIMEBOOST_net_20288), .o(TIMEBOOST_net_17005) );
na02m04 g53945_u1 ( .a(conf_wb_err_bc_in), .b(g53939_sb), .o(g53945_da) );
na04f04 TIMEBOOST_cell_25002 ( .a(n_10599), .b(n_10596), .c(n_10010), .d(n_10014), .o(n_12141) );
na04f04 TIMEBOOST_cell_67543 ( .a(g61875_sb), .b(FE_OFN706_n_8119), .c(n_1896), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q), .o(n_8082) );
in01m01 g53946_u0 ( .a(FE_OFN2072_n_15978), .o(g53946_sb) );
na02m02 g53946_u1 ( .a(wishbone_slave_unit_pci_initiator_if_current_byte_address), .b(g53946_sb), .o(g53946_da) );
na03m02 TIMEBOOST_cell_73005 ( .a(TIMEBOOST_net_16600), .b(TIMEBOOST_net_7092), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q), .o(TIMEBOOST_net_22130) );
na03f02 TIMEBOOST_cell_66521 ( .a(TIMEBOOST_net_21041), .b(FE_OFN1330_n_13547), .c(g53900_sb), .o(n_13543) );
na03f02 TIMEBOOST_cell_66855 ( .a(TIMEBOOST_net_20667), .b(n_14971), .c(g58653_sb), .o(n_9236) );
na03s01 TIMEBOOST_cell_42002 ( .a(FE_OFN252_n_9868), .b(g58258_sb), .c(g58258_db), .o(n_9539) );
na02f02 TIMEBOOST_cell_71065 ( .a(TIMEBOOST_net_22740), .b(g63180_sb), .o(n_5790) );
na02m10 TIMEBOOST_cell_62606 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q), .b(pci_target_unit_fifos_pciw_cbe_in_154), .o(TIMEBOOST_net_20250) );
na02m02 TIMEBOOST_cell_69125 ( .a(TIMEBOOST_net_21770), .b(TIMEBOOST_net_20242), .o(TIMEBOOST_net_17100) );
na03s02 TIMEBOOST_cell_46547 ( .a(TIMEBOOST_net_12975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q), .c(g58282_sb), .o(TIMEBOOST_net_9552) );
na03f02 TIMEBOOST_cell_66028 ( .a(n_14681), .b(n_14839), .c(TIMEBOOST_net_20942), .o(TIMEBOOST_net_15556) );
na03f02 TIMEBOOST_cell_34893 ( .a(TIMEBOOST_net_9328), .b(FE_OFN1396_n_8567), .c(g57571_sb), .o(n_11180) );
na02s02 TIMEBOOST_cell_68133 ( .a(TIMEBOOST_net_21274), .b(TIMEBOOST_net_6804), .o(TIMEBOOST_net_16803) );
na02s01 TIMEBOOST_cell_37040 ( .a(pci_ad_i_9_), .b(parchk_pci_ad_reg_in_1213), .o(TIMEBOOST_net_10132) );
na02f02 TIMEBOOST_cell_69815 ( .a(TIMEBOOST_net_22115), .b(n_4450), .o(TIMEBOOST_net_17431) );
na02m02 TIMEBOOST_cell_68735 ( .a(TIMEBOOST_net_21575), .b(TIMEBOOST_net_10455), .o(TIMEBOOST_net_20588) );
na02s02 TIMEBOOST_cell_53561 ( .a(g57905_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q), .o(TIMEBOOST_net_16998) );
na02f02 TIMEBOOST_cell_50484 ( .a(TIMEBOOST_net_15459), .b(g62585_sb), .o(n_6382) );
na02f01 g62805_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN1134_g64577_p), .o(g62805_db) );
na02f01 g62757_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q), .b(FE_OFN1125_g64577_p), .o(g62757_db) );
in01f08 g53980_u0 ( .a(n_13679), .o(n_13625) );
na03f02 TIMEBOOST_cell_73791 ( .a(TIMEBOOST_net_16543), .b(FE_OFN1600_n_13995), .c(FE_OCPN2218_n_13997), .o(g53163_p) );
na02f02 g58800_u2 ( .a(n_3485), .b(FE_OFN1697_n_5751), .o(g58800_db) );
na03m02 TIMEBOOST_cell_72850 ( .a(g64756_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q), .c(TIMEBOOST_net_16237), .o(TIMEBOOST_net_17146) );
na03s02 TIMEBOOST_cell_41948 ( .a(FE_OFN221_n_9846), .b(g57926_sb), .c(g57926_db), .o(n_9883) );
no02f06 g53988_u0 ( .a(n_15370), .b(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .o(n_1645) );
na02f02 g53990_u0 ( .a(n_1684), .b(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .o(g53990_p) );
in01f02 g53990_u1 ( .a(g53990_p), .o(n_1979) );
no02f01 g53991_u0 ( .a(n_13329), .b(n_1041), .o(n_13494) );
no02f01 g53992_u0 ( .a(n_13328), .b(n_1041), .o(n_13493) );
no02f01 g53993_u0 ( .a(n_13327), .b(n_1041), .o(n_13491) );
na03s02 TIMEBOOST_cell_72302 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q), .b(FE_OFN268_n_9880), .c(FE_OFN592_n_9694), .o(TIMEBOOST_net_23359) );
na02m08 TIMEBOOST_cell_42951 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q), .o(TIMEBOOST_net_12370) );
na02m02 TIMEBOOST_cell_62829 ( .a(TIMEBOOST_net_20361), .b(FE_OFN1037_n_4732), .o(TIMEBOOST_net_14752) );
na02f01 TIMEBOOST_cell_62455 ( .a(TIMEBOOST_net_20174), .b(FE_OFN905_n_4736), .o(TIMEBOOST_net_14139) );
in01f40 g53_u0 ( .a(n_15929), .o(n_4743) );
na04f04 TIMEBOOST_cell_25004 ( .a(n_9315), .b(n_10188), .c(n_10183), .d(n_9319), .o(n_12161) );
na04s02 TIMEBOOST_cell_67487 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q), .b(FE_OFN588_n_9692), .c(TIMEBOOST_net_20377), .d(g58188_sb), .o(TIMEBOOST_net_9542) );
na02s01 TIMEBOOST_cell_48015 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_143), .o(TIMEBOOST_net_14225) );
na02s02 TIMEBOOST_cell_71305 ( .a(TIMEBOOST_net_22860), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_14927) );
na02f02 TIMEBOOST_cell_70169 ( .a(TIMEBOOST_net_22292), .b(g64088_sb), .o(n_4067) );
na02m01 TIMEBOOST_cell_25290 ( .a(TIMEBOOST_net_6749), .b(n_574), .o(TIMEBOOST_net_5356) );
na02m02 TIMEBOOST_cell_69689 ( .a(TIMEBOOST_net_22052), .b(g65384_sb), .o(TIMEBOOST_net_12756) );
na03s02 TIMEBOOST_cell_73352 ( .a(FE_OFN528_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q), .c(g58031_sb), .o(TIMEBOOST_net_14636) );
na02s01 TIMEBOOST_cell_62438 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q), .b(g65865_sb), .o(TIMEBOOST_net_20166) );
in01m04 TIMEBOOST_cell_67745 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .o(TIMEBOOST_net_21172) );
ao12f02 g54015_u0 ( .a(n_7084), .b(n_13027), .c(n_13354), .o(n_13355) );
ao12f02 g54016_u0 ( .a(n_7083), .b(n_13026), .c(n_7822), .o(n_13353) );
ao12f02 g54018_u0 ( .a(n_7082), .b(n_13022), .c(n_13354), .o(n_13350) );
ao12f02 g54019_u0 ( .a(n_7081), .b(n_13020), .c(n_13354), .o(n_13349) );
ao12f02 g54020_u0 ( .a(n_7080), .b(n_13018), .c(n_13354), .o(n_13348) );
na02s02 g54022_u0 ( .a(n_2027), .b(wbm_cyc_o), .o(n_13789) );
ao12f02 g54023_u0 ( .a(n_7320), .b(n_12985), .c(n_7822), .o(n_13346) );
in01f01 g54024_u0 ( .a(n_13813), .o(n_13732) );
no02f02 g54025_u0 ( .a(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .b(wishbone_slave_unit_wbs_sm_wbr_control_in), .o(n_13813) );
ao12f02 g54029_u0 ( .a(n_7707), .b(n_13098), .c(n_13354), .o(n_13417) );
in01f01 g54030_u0 ( .a(n_12595), .o(g54030_sb) );
na03m02 TIMEBOOST_cell_72561 ( .a(TIMEBOOST_net_21441), .b(FE_OFN684_n_4417), .c(TIMEBOOST_net_21600), .o(TIMEBOOST_net_17520) );
na02s01 TIMEBOOST_cell_63625 ( .a(TIMEBOOST_net_20798), .b(g54207_da), .o(TIMEBOOST_net_13450) );
na03f02 TIMEBOOST_cell_47314 ( .a(FE_OFN1553_n_12104), .b(TIMEBOOST_net_13598), .c(FE_OCP_RBN1977_n_10273), .o(n_12520) );
ao22f02 g54031_u0 ( .a(n_7338), .b(n_13415), .c(n_13102), .d(n_13341), .o(n_13416) );
ao22f02 g54032_u0 ( .a(n_7504), .b(n_13415), .c(n_13012), .d(n_13341), .o(n_13342) );
ao22f02 g54033_u0 ( .a(n_12986), .b(n_13341), .c(n_8488), .d(n_13415), .o(n_13340) );
ao12f02 g54034_u0 ( .a(n_7046), .b(n_12998), .c(n_13354), .o(n_13339) );
ao12f02 g54035_u0 ( .a(n_7045), .b(n_12994), .c(n_13354), .o(n_13338) );
ao12f02 g54036_u0 ( .a(n_7075), .b(n_12992), .c(n_13354), .o(n_13337) );
in01m20 g54038_u0 ( .a(parchk_pci_par_en_in), .o(g54038_sb) );
na02m02 TIMEBOOST_cell_50036 ( .a(TIMEBOOST_net_15235), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_13316) );
na02m40 g54038_u2 ( .a(pci_par_i), .b(parchk_pci_par_en_in), .o(g54038_db) );
na02m10 TIMEBOOST_cell_52993 ( .a(wishbone_slave_unit_pcim_sm_data_in_637), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q), .o(TIMEBOOST_net_16714) );
in01f02 g54039_u0 ( .a(n_12595), .o(g54039_sb) );
in01f04 g54040_u0 ( .a(n_7822), .o(g54040_sb) );
na02f04 TIMEBOOST_cell_63798 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_411), .b(n_1793), .o(TIMEBOOST_net_20885) );
na02s01 TIMEBOOST_cell_53529 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q), .o(TIMEBOOST_net_16982) );
in01s01 g54044_u0 ( .a(wbm_cyc_o_1378), .o(wbm_cyc_o) );
na02s01 TIMEBOOST_cell_49530 ( .a(TIMEBOOST_net_14982), .b(FE_OFN555_n_9864), .o(TIMEBOOST_net_12966) );
na02s02 TIMEBOOST_cell_49727 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q), .b(g58286_sb), .o(TIMEBOOST_net_15081) );
na02s01 TIMEBOOST_cell_42967 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_137), .o(TIMEBOOST_net_12378) );
na02s01 TIMEBOOST_cell_47517 ( .a(parchk_pci_ad_reg_in_1210), .b(g67042_db), .o(TIMEBOOST_net_13976) );
na02s01 TIMEBOOST_cell_62479 ( .a(TIMEBOOST_net_20186), .b(wishbone_slave_unit_delayed_write_data_comp_wdata_out_81), .o(TIMEBOOST_net_14101) );
na02s01 TIMEBOOST_cell_47516 ( .a(TIMEBOOST_net_13975), .b(g67049_sb), .o(n_1274) );
in01m01 g54125_u0 ( .a(n_13332), .o(n_13333) );
ao12f02 g54127_u0 ( .a(n_13306), .b(n_13486), .c(wbm_sel_o_0_), .o(n_13488) );
ao12f02 g54128_u0 ( .a(n_13305), .b(n_13486), .c(wbm_sel_o_1_), .o(n_13487) );
ao12f02 g54129_u0 ( .a(n_13303), .b(n_13486), .c(wbm_sel_o_2_), .o(n_13485) );
ao12f02 g54130_u0 ( .a(n_13302), .b(n_13486), .c(wbm_sel_o_3_), .o(n_13484) );
in01f06 g54131_u0 ( .a(FE_OFN2125_n_16497), .o(g54131_sb) );
na02f08 g54131_u1 ( .a(n_13145), .b(g54131_sb), .o(g54131_da) );
na03f02 TIMEBOOST_cell_24838 ( .a(n_14895), .b(n_13485), .c(n_14830), .o(n_14896) );
na02m02 TIMEBOOST_cell_68792 ( .a(g65086_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q), .o(TIMEBOOST_net_21604) );
in01f02 g54132_u0 ( .a(FE_OFN1150_n_13249), .o(g54132_sb) );
na02s01 TIMEBOOST_cell_45285 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q), .o(TIMEBOOST_net_13537) );
in01f04 g54133_u0 ( .a(FE_OFN1150_n_13249), .o(g54133_sb) );
na04f04 TIMEBOOST_cell_36866 ( .a(TIMEBOOST_net_9618), .b(FE_OFN2200_n_10256), .c(g52602_sb), .d(TIMEBOOST_net_711), .o(n_11869) );
na02f02 TIMEBOOST_cell_70365 ( .a(TIMEBOOST_net_22390), .b(g63621_sb), .o(n_7174) );
in01f02 g54134_u0 ( .a(FE_OFN1151_n_13249), .o(g54134_sb) );
na02f02 TIMEBOOST_cell_70844 ( .a(TIMEBOOST_net_16695), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_22630) );
na02s01 TIMEBOOST_cell_70460 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q), .b(FE_OFN1649_n_9428), .o(TIMEBOOST_net_22438) );
na03f02 TIMEBOOST_cell_73591 ( .a(TIMEBOOST_net_17325), .b(FE_OFN1135_g64577_p), .c(g63053_sb), .o(n_5143) );
in01f02 g54135_u0 ( .a(FE_OFN1149_n_13249), .o(g54135_sb) );
na02s02 TIMEBOOST_cell_64037 ( .a(TIMEBOOST_net_21004), .b(g57914_sb), .o(TIMEBOOST_net_9490) );
na02s01 TIMEBOOST_cell_28971 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_), .o(TIMEBOOST_net_8590) );
na02f01 TIMEBOOST_cell_37300 ( .a(n_12179), .b(n_2315), .o(TIMEBOOST_net_10262) );
in01f04 g54137_u0 ( .a(FE_OFN1148_n_13249), .o(g54137_sb) );
na03s02 TIMEBOOST_cell_70064 ( .a(n_1936), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q), .c(FE_OFN2257_n_8060), .o(TIMEBOOST_net_22240) );
na04f06 TIMEBOOST_cell_64382 ( .a(FE_RN_313_0), .b(FE_RN_323_0), .c(FE_RN_354_0), .d(FE_RN_333_0), .o(FE_RN_355_0) );
na02s02 TIMEBOOST_cell_53562 ( .a(TIMEBOOST_net_16998), .b(TIMEBOOST_net_10316), .o(TIMEBOOST_net_9322) );
in01f02 g54138_u0 ( .a(FE_OFN1149_n_13249), .o(g54138_sb) );
na03s02 TIMEBOOST_cell_21308 ( .a(FE_OFN217_n_9889), .b(g58113_sb), .c(g58113_db), .o(n_9682) );
na02f02 g54139_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_404), .b(FE_OCPN1910_FE_OFN1152_n_13249), .o(g54139_da) );
na02f01 TIMEBOOST_cell_68900 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q), .b(FE_OFN1643_n_4671), .o(TIMEBOOST_net_21658) );
na02f02 TIMEBOOST_cell_71067 ( .a(TIMEBOOST_net_22741), .b(g62643_sb), .o(n_7371) );
in01f02 g54140_u0 ( .a(FE_OFN1150_n_13249), .o(g54140_sb) );
na02m02 TIMEBOOST_cell_68981 ( .a(TIMEBOOST_net_21698), .b(g65294_sb), .o(TIMEBOOST_net_12592) );
na03f02 TIMEBOOST_cell_73592 ( .a(TIMEBOOST_net_17415), .b(FE_OFN1253_n_4143), .c(g62499_sb), .o(n_6585) );
in01f04 g54141_u0 ( .a(FE_OFN1151_n_13249), .o(g54141_sb) );
na03f02 TIMEBOOST_cell_66090 ( .a(TIMEBOOST_net_20934), .b(FE_OFN1688_n_9528), .c(g58274_sb), .o(n_9035) );
na04f04 TIMEBOOST_cell_65711 ( .a(TIMEBOOST_net_7209), .b(FE_OFN1144_n_15261), .c(TIMEBOOST_net_658), .d(g54202_da), .o(TIMEBOOST_net_16463) );
in01f02 g54143_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54143_sb) );
na02s01 TIMEBOOST_cell_37310 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q), .b(pci_target_unit_fifos_pcir_data_in_165), .o(TIMEBOOST_net_10267) );
na03m02 TIMEBOOST_cell_72486 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q), .b(n_3752), .c(TIMEBOOST_net_21581), .o(TIMEBOOST_net_17523) );
in01f02 g54144_u0 ( .a(FE_OFN1147_n_13249), .o(g54144_sb) );
na03f02 TIMEBOOST_cell_67926 ( .a(n_3894), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q), .c(FE_OFN882_g64577_p), .o(TIMEBOOST_net_13188) );
na03f02 TIMEBOOST_cell_34895 ( .a(TIMEBOOST_net_9326), .b(FE_OFN1414_n_8567), .c(g57412_sb), .o(n_11330) );
in01f02 g54145_u0 ( .a(FE_OFN1149_n_13249), .o(g54145_sb) );
na02m01 TIMEBOOST_cell_53427 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_142), .o(TIMEBOOST_net_16931) );
na03m02 TIMEBOOST_cell_65807 ( .a(g58363_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q), .c(TIMEBOOST_net_15024), .o(TIMEBOOST_net_9483) );
in01f02 g54146_u0 ( .a(FE_OFN1150_n_13249), .o(g54146_sb) );
na02m10 TIMEBOOST_cell_52677 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_16556) );
na02s01 TIMEBOOST_cell_68189 ( .a(TIMEBOOST_net_21302), .b(FE_OFN936_n_2292), .o(TIMEBOOST_net_14093) );
in01f02 g54147_u0 ( .a(FE_OFN1149_n_13249), .o(g54147_sb) );
na02s02 TIMEBOOST_cell_42826 ( .a(TIMEBOOST_net_12307), .b(n_539), .o(n_9830) );
in01s01 TIMEBOOST_cell_45884 ( .a(TIMEBOOST_net_13844), .o(TIMEBOOST_net_13845) );
in01f02 g54148_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54148_sb) );
no04f06 TIMEBOOST_cell_20809 ( .a(n_2818), .b(n_231), .c(FE_RN_669_0), .d(FE_RN_674_0), .o(TIMEBOOST_net_119) );
na03f02 TIMEBOOST_cell_34852 ( .a(TIMEBOOST_net_9446), .b(FE_OFN1389_n_8567), .c(g57463_sb), .o(n_11270) );
na04f02 TIMEBOOST_cell_72480 ( .a(TIMEBOOST_net_12330), .b(FE_OFN906_n_4736), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q), .d(g64148_sb), .o(TIMEBOOST_net_13098) );
in01f02 g54149_u0 ( .a(FE_OFN1151_n_13249), .o(g54149_sb) );
na02s01 TIMEBOOST_cell_42787 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q), .o(TIMEBOOST_net_12288) );
na02s01 TIMEBOOST_cell_45651 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q), .o(TIMEBOOST_net_13720) );
in01f02 g54150_u0 ( .a(FE_OFN1150_n_13249), .o(g54150_sb) );
na02m01 TIMEBOOST_cell_70126 ( .a(n_4470), .b(n_18), .o(TIMEBOOST_net_22271) );
na04f04 TIMEBOOST_cell_25006 ( .a(n_10066), .b(n_9271), .c(n_10641), .d(n_9272), .o(n_12147) );
in01f02 g54151_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54151_sb) );
na03f02 TIMEBOOST_cell_66857 ( .a(TIMEBOOST_net_20665), .b(n_14971), .c(g58600_sb), .o(n_9239) );
na03m02 TIMEBOOST_cell_72562 ( .a(TIMEBOOST_net_23133), .b(FE_OFN630_n_4454), .c(TIMEBOOST_net_21509), .o(TIMEBOOST_net_17110) );
in01f04 g54152_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54152_sb) );
na02f02 TIMEBOOST_cell_64014 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_del_addr_hit), .o(TIMEBOOST_net_20993) );
na03s02 TIMEBOOST_cell_72910 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q), .b(g65976_sb), .c(TIMEBOOST_net_23236), .o(n_1838) );
na03s02 TIMEBOOST_cell_72902 ( .a(n_1583), .b(g61932_sb), .c(g61932_db), .o(n_7959) );
in01f02 g54153_u0 ( .a(FE_OFN1148_n_13249), .o(g54153_sb) );
na02m01 TIMEBOOST_cell_53415 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN612_n_4501), .o(TIMEBOOST_net_16925) );
na03m02 TIMEBOOST_cell_72689 ( .a(TIMEBOOST_net_23137), .b(g65962_db), .c(TIMEBOOST_net_22777), .o(n_7895) );
in01m02 g54154_u0 ( .a(FE_OFN1148_n_13249), .o(g54154_sb) );
na03f02 TIMEBOOST_cell_66668 ( .a(TIMEBOOST_net_17427), .b(FE_OFN1218_n_6886), .c(g62603_sb), .o(n_6345) );
na03f02 TIMEBOOST_cell_73043 ( .a(TIMEBOOST_net_22041), .b(FE_OFN717_n_8176), .c(g61759_sb), .o(n_8295) );
na02f01 g62789_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN1124_g64577_p), .o(g62789_db) );
in01f06 g54155_u0 ( .a(FE_OFN1151_n_13249), .o(g54155_sb) );
na02f10 TIMEBOOST_cell_42773 ( .a(n_15417), .b(n_16854), .o(TIMEBOOST_net_12281) );
in01s01 TIMEBOOST_cell_67747 ( .a(pci_target_unit_fifos_pcir_data_in_180), .o(TIMEBOOST_net_21174) );
na02m02 TIMEBOOST_cell_71989 ( .a(TIMEBOOST_net_23202), .b(FE_OFN640_n_4669), .o(TIMEBOOST_net_16251) );
in01f01 g54157_u0 ( .a(FE_OFN1151_n_13249), .o(g54157_sb) );
na02f20 TIMEBOOST_cell_53439 ( .a(configuration_pci_err_data_509), .b(pciu_am1_in), .o(TIMEBOOST_net_16937) );
na02s02 TIMEBOOST_cell_63668 ( .a(g57971_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q), .o(TIMEBOOST_net_20820) );
in01f06 g54158_u0 ( .a(FE_OFN1147_n_13249), .o(g54158_sb) );
in01s01 TIMEBOOST_cell_63588 ( .a(TIMEBOOST_net_20768), .o(TIMEBOOST_net_20743) );
na03f02 TIMEBOOST_cell_67054 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_16541), .c(FE_OFN1600_n_13995), .o(FE_RN_890_0) );
in01f01 g54159_u0 ( .a(n_13548), .o(n_13329) );
in01m40 g54160_u0 ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .o(g54160_sb) );
in01s01 TIMEBOOST_cell_73869 ( .a(TIMEBOOST_net_23433), .o(TIMEBOOST_net_23434) );
na03f02 TIMEBOOST_cell_34992 ( .a(TIMEBOOST_net_9568), .b(g57112_sb), .c(FE_OFN2187_n_8567), .o(n_11634) );
na03f02 TIMEBOOST_cell_34994 ( .a(TIMEBOOST_net_9570), .b(g57568_sb), .c(FE_OFN1376_n_8567), .o(n_11184) );
in01f06 g54161_u0 ( .a(FE_OFN1147_n_13249), .o(g54161_sb) );
na02m02 TIMEBOOST_cell_44905 ( .a(TIMEBOOST_net_9942), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_13347) );
na02s01 TIMEBOOST_cell_71306 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q), .b(FE_OFN556_n_9864), .o(TIMEBOOST_net_22861) );
na03f02 TIMEBOOST_cell_66836 ( .a(TIMEBOOST_net_16844), .b(FE_OFN1345_n_8567), .c(g57117_sb), .o(n_10477) );
in01f01 g54162_u0 ( .a(n_13544), .o(n_13328) );
na02f40 g54163_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_cbe_in_416), .b(FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54163_da) );
in01s02 TIMEBOOST_cell_31890 ( .a(TIMEBOOST_net_10053), .o(TIMEBOOST_net_10054) );
in01f08 g54164_u0 ( .a(FE_OFN1147_n_13249), .o(g54164_sb) );
na02s01 TIMEBOOST_cell_42958 ( .a(TIMEBOOST_net_12373), .b(FE_OFN950_n_2055), .o(TIMEBOOST_net_10531) );
na03f02 TIMEBOOST_cell_34973 ( .a(TIMEBOOST_net_9479), .b(FE_OFN1412_n_8567), .c(g57065_sb), .o(n_10499) );
in01f01 g54165_u0 ( .a(n_13541), .o(n_13327) );
in01s01 TIMEBOOST_cell_73870 ( .a(n_7857), .o(TIMEBOOST_net_23435) );
in01s01 TIMEBOOST_cell_31891 ( .a(TIMEBOOST_net_10055), .o(wbs_dat_i_20_) );
na02s02 TIMEBOOST_cell_30597 ( .a(n_9418), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q), .o(TIMEBOOST_net_9403) );
in01s02 g54167_u0 ( .a(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54167_sb) );
na03f02 TIMEBOOST_cell_66317 ( .a(TIMEBOOST_net_17144), .b(n_6319), .c(g62619_sb), .o(n_6321) );
na02s01 g54167_u2 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_88), .b(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54167_db) );
na02s01 TIMEBOOST_cell_51585 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q), .o(TIMEBOOST_net_16010) );
in01f02 g54168_u0 ( .a(FE_OFN1083_n_13221), .o(g54168_sb) );
na03f03 TIMEBOOST_cell_73745 ( .a(TIMEBOOST_net_13670), .b(FE_OFN1757_n_12681), .c(FE_OCP_RBN1976_n_12381), .o(n_17029) );
na03f02 TIMEBOOST_cell_66319 ( .a(TIMEBOOST_net_17052), .b(n_6287), .c(g62368_sb), .o(n_6867) );
in01f02 g54169_u0 ( .a(FE_OFN1083_n_13221), .o(g54169_sb) );
na03s01 TIMEBOOST_cell_20811 ( .a(wishbone_slave_unit_wishbone_slave_pref_en_reg_Q), .b(TIMEBOOST_net_513), .c(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q), .o(n_1721) );
na02f10 g74951_u0 ( .a(n_16565), .b(FE_OCPN1823_n_16560), .o(n_16322) );
na02m01 TIMEBOOST_cell_62635 ( .a(TIMEBOOST_net_20264), .b(FE_OFN930_n_4730), .o(TIMEBOOST_net_16290) );
in01f02 g54170_u0 ( .a(FE_OFN1083_n_13221), .o(g54170_sb) );
na03s02 TIMEBOOST_cell_68414 ( .a(TIMEBOOST_net_8191), .b(g65867_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q), .o(TIMEBOOST_net_21415) );
na02s02 TIMEBOOST_cell_49613 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q), .b(g58363_sb), .o(TIMEBOOST_net_15024) );
na04f04 TIMEBOOST_cell_25008 ( .a(n_10944), .b(n_9290), .c(n_9293), .d(n_10102), .o(n_12153) );
in01m08 g54171_u0 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54171_sb) );
na04s02 TIMEBOOST_cell_33414 ( .a(FE_OFN268_n_9880), .b(g58153_sb), .c(g58153_db), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q), .o(TIMEBOOST_net_9569) );
na03s02 TIMEBOOST_cell_41735 ( .a(g58318_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q), .c(g58318_db), .o(n_9494) );
in01m01 g54172_u0 ( .a(FE_OFN1082_n_13221), .o(g54172_sb) );
na02f06 FE_RC_500_0 ( .a(FE_RN_302_0), .b(n_15458), .o(n_16976) );
na02s01 TIMEBOOST_cell_25301 ( .a(pci_ad_i_13_), .b(parchk_pci_ad_reg_in_1217), .o(TIMEBOOST_net_6755) );
in01m01 g54173_u0 ( .a(FE_OFN1082_n_13221), .o(g54173_sb) );
na02f02 g54314_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q), .b(FE_OFN2126_n_16497), .o(g54314_db) );
in01f01 g54174_u0 ( .a(n_13221), .o(g54174_sb) );
na02m01 TIMEBOOST_cell_69440 ( .a(n_4645), .b(n_4312), .o(TIMEBOOST_net_21928) );
na02f02 g54174_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_2__Q), .b(n_13221), .o(g54174_db) );
na02f02 TIMEBOOST_cell_72260 ( .a(TIMEBOOST_net_17018), .b(FE_OFN1226_n_6391), .o(TIMEBOOST_net_23338) );
in01f01 g54175_u0 ( .a(n_13221), .o(g54175_sb) );
na02f02 g54175_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_395), .b(g54175_sb), .o(g54175_da) );
na02s02 TIMEBOOST_cell_52471 ( .a(g58215_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_16453) );
na04m08 TIMEBOOST_cell_73086 ( .a(n_3785), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q), .c(FE_OFN1806_n_4501), .d(g64763_sb), .o(n_3786) );
in01f04 g54176_u0 ( .a(FE_OFN1085_n_13221), .o(g54176_sb) );
na03s02 TIMEBOOST_cell_73656 ( .a(FE_OFN532_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q), .c(TIMEBOOST_net_22922), .o(TIMEBOOST_net_21067) );
na02f02 TIMEBOOST_cell_50242 ( .a(TIMEBOOST_net_15338), .b(g62438_sb), .o(n_6720) );
in01f02 g54177_u0 ( .a(FE_OFN1082_n_13221), .o(g54177_sb) );
na02f02 TIMEBOOST_cell_53646 ( .a(TIMEBOOST_net_17040), .b(g62923_sb), .o(n_6035) );
in01f02 g54178_u0 ( .a(FE_OFN1082_n_13221), .o(g54178_sb) );
na02f04 g54178_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_398), .b(g54178_sb), .o(g54178_da) );
na02f02 TIMEBOOST_cell_70367 ( .a(TIMEBOOST_net_22391), .b(g63617_sb), .o(n_7157) );
in01f02 g54179_u0 ( .a(FE_OFN1084_n_13221), .o(g54179_sb) );
na02m06 TIMEBOOST_cell_54117 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_132), .o(TIMEBOOST_net_17276) );
na02m04 TIMEBOOST_cell_52695 ( .a(n_3007), .b(n_2281), .o(TIMEBOOST_net_16565) );
na02s02 TIMEBOOST_cell_47863 ( .a(TIMEBOOST_net_21151), .b(g65795_sb), .o(TIMEBOOST_net_14149) );
in01f02 g54180_u0 ( .a(n_13221), .o(g54180_sb) );
na02f02 g54180_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_17__Q), .b(n_13221), .o(g54180_db) );
in01f04 g54181_u0 ( .a(FE_OFN1084_n_13221), .o(g54181_sb) );
na02f06 g54181_u1 ( .a(g54181_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_401), .o(g54181_da) );
na02m02 TIMEBOOST_cell_69416 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q), .o(TIMEBOOST_net_21916) );
na02s01 TIMEBOOST_cell_25305 ( .a(pci_ad_i_17_), .b(parchk_pci_ad_reg_in_1221), .o(TIMEBOOST_net_6757) );
in01m01 g54182_u0 ( .a(n_13221), .o(g54182_sb) );
na03f04 TIMEBOOST_cell_67006 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_16519), .c(FE_OFN1587_n_13736), .o(g53288_p) );
na02m02 g54182_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_19__Q), .b(n_13221), .o(g54182_db) );
na02f04 TIMEBOOST_cell_49996 ( .a(TIMEBOOST_net_15215), .b(g54237_sb), .o(n_13651) );
in01f02 g54183_u0 ( .a(FE_OFN1084_n_13221), .o(g54183_sb) );
na03s02 TIMEBOOST_cell_41953 ( .a(FE_OFN215_n_9856), .b(g58175_sb), .c(g58175_db), .o(n_9615) );
na03m02 TIMEBOOST_cell_73205 ( .a(TIMEBOOST_net_22063), .b(FE_OFN699_n_7845), .c(g61890_sb), .o(n_8049) );
na02f02 TIMEBOOST_cell_28004 ( .a(n_13901), .b(TIMEBOOST_net_8106), .o(TIMEBOOST_net_759) );
in01m01 g54184_u0 ( .a(n_13221), .o(g54184_sb) );
na02m06 TIMEBOOST_cell_69691 ( .a(TIMEBOOST_net_22053), .b(g65396_sb), .o(TIMEBOOST_net_12758) );
na02m01 g54184_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_21__Q), .b(n_13221), .o(g54184_db) );
na02s01 TIMEBOOST_cell_47835 ( .a(TIMEBOOST_net_13831), .b(g65717_sb), .o(TIMEBOOST_net_14135) );
in01f02 g54185_u0 ( .a(n_13221), .o(g54185_sb) );
na02f02 g54185_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_3__Q), .b(n_13221), .o(g54185_db) );
na02f02 TIMEBOOST_cell_72307 ( .a(TIMEBOOST_net_23361), .b(TIMEBOOST_net_14929), .o(TIMEBOOST_net_9513) );
in01m01 g54186_u0 ( .a(FE_OFN1084_n_13221), .o(g54186_sb) );
na02s01 TIMEBOOST_cell_28005 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q), .o(TIMEBOOST_net_8107) );
in01m02 g54187_u0 ( .a(FE_OFN1085_n_13221), .o(g54187_sb) );
na03s01 TIMEBOOST_cell_41920 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q), .b(g58356_sb), .c(g58356_db), .o(n_9466) );
na02s01 TIMEBOOST_cell_43445 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q), .o(TIMEBOOST_net_12617) );
in01m01 g54188_u0 ( .a(n_13221), .o(g54188_sb) );
na02m02 g54188_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_24__Q), .b(n_13221), .o(g54188_db) );
na02m10 TIMEBOOST_cell_52955 ( .a(wishbone_slave_unit_pcim_sm_data_in_648), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q), .o(TIMEBOOST_net_16695) );
in01m01 g54189_u0 ( .a(n_13221), .o(g54189_sb) );
na02m02 g54189_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_25__Q), .b(n_13221), .o(g54189_db) );
in01s01 TIMEBOOST_cell_67749 ( .a(pci_target_unit_fifos_pcir_data_in_163), .o(TIMEBOOST_net_21176) );
in01f02 g54190_u0 ( .a(FE_OFN1085_n_13221), .o(g54190_sb) );
na02m01 TIMEBOOST_cell_42889 ( .a(n_2284), .b(n_657), .o(TIMEBOOST_net_12339) );
na03s02 TIMEBOOST_cell_65525 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q), .b(g58285_sb), .c(TIMEBOOST_net_11114), .o(TIMEBOOST_net_9519) );
na02s02 TIMEBOOST_cell_44447 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q), .b(g58317_sb), .o(TIMEBOOST_net_13118) );
in01f02 g54191_u0 ( .a(FE_OFN1085_n_13221), .o(g54191_sb) );
na03m02 TIMEBOOST_cell_69222 ( .a(n_4476), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q), .c(FE_OFN642_n_4677), .o(TIMEBOOST_net_21819) );
in01m02 g54192_u0 ( .a(FE_OFN1082_n_13221), .o(g54192_sb) );
na02s01 TIMEBOOST_cell_38826 ( .a(FE_OFN1025_n_11877), .b(wbu_addr_in_257), .o(TIMEBOOST_net_11025) );
na02m02 TIMEBOOST_cell_40023 ( .a(TIMEBOOST_net_11623), .b(g63183_sb), .o(n_5786) );
na03s02 TIMEBOOST_cell_65196 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q), .b(g65954_sb), .c(TIMEBOOST_net_20378), .o(TIMEBOOST_net_10838) );
in01m02 g54193_u0 ( .a(FE_OFN1084_n_13221), .o(g54193_sb) );
na03f02 TIMEBOOST_cell_73449 ( .a(TIMEBOOST_net_20544), .b(FE_OFN1269_n_4095), .c(g62333_sb), .o(n_6934) );
in01m01 g54194_u0 ( .a(n_13221), .o(g54194_sb) );
na02f02 TIMEBOOST_cell_70369 ( .a(TIMEBOOST_net_22392), .b(g63604_sb), .o(n_7168) );
na02m01 TIMEBOOST_cell_25292 ( .a(TIMEBOOST_net_6750), .b(n_574), .o(TIMEBOOST_net_5359) );
in01m02 g54195_u0 ( .a(FE_OFN1082_n_13221), .o(g54195_sb) );
na03f02 TIMEBOOST_cell_34886 ( .a(TIMEBOOST_net_9331), .b(FE_OFN1370_n_8567), .c(g57519_sb), .o(n_10317) );
in01f08 TIMEBOOST_cell_35474 ( .a(TIMEBOOST_net_10065), .o(n_3157) );
na02m02 TIMEBOOST_cell_44448 ( .a(TIMEBOOST_net_13118), .b(TIMEBOOST_net_11171), .o(TIMEBOOST_net_9528) );
in01f01 g54196_u0 ( .a(n_13221), .o(g54196_sb) );
na02s01 TIMEBOOST_cell_63838 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q), .o(TIMEBOOST_net_20905) );
no02f01 TIMEBOOST_cell_47771 ( .a(n_1014), .b(FE_OCPN1832_n_16949), .o(TIMEBOOST_net_14103) );
in01f02 g54197_u0 ( .a(FE_OFN1082_n_13221), .o(g54197_sb) );
na02m02 TIMEBOOST_cell_69664 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q), .b(FE_OFN702_n_7845), .o(TIMEBOOST_net_22040) );
na02s01 TIMEBOOST_cell_47994 ( .a(TIMEBOOST_net_14214), .b(TIMEBOOST_net_10353), .o(TIMEBOOST_net_9327) );
na04m06 TIMEBOOST_cell_72628 ( .a(g64903_sb), .b(n_3792), .c(n_3691), .d(g64903_db), .o(TIMEBOOST_net_17518) );
in01m01 g54198_u0 ( .a(n_13221), .o(g54198_sb) );
na03f10 TIMEBOOST_cell_41276 ( .a(n_15330), .b(n_2092), .c(n_16936), .o(n_3395) );
in01m01 g54199_u0 ( .a(n_13221), .o(g54199_sb) );
na03f08 TIMEBOOST_cell_46050 ( .a(FE_RN_83_0), .b(n_2380), .c(n_7092), .o(n_16325) );
na03m02 TIMEBOOST_cell_72474 ( .a(TIMEBOOST_net_12326), .b(FE_OFN902_n_4736), .c(g64122_sb), .o(TIMEBOOST_net_14971) );
na02s01 TIMEBOOST_cell_45371 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_13580) );
in01f02 g54200_u0 ( .a(FE_OFN1082_n_13221), .o(g54200_sb) );
na03f02 TIMEBOOST_cell_34888 ( .a(TIMEBOOST_net_9389), .b(FE_OFN1392_n_8567), .c(g57081_sb), .o(n_11661) );
na02f04 TIMEBOOST_cell_71328 ( .a(wishbone_slave_unit_pcim_if_wbw_cbe_in), .b(g54168_sb), .o(TIMEBOOST_net_22872) );
in01m01 g54201_u0 ( .a(n_13221), .o(g54201_sb) );
na02m04 TIMEBOOST_cell_68710 ( .a(FE_OFN684_n_4417), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q), .o(TIMEBOOST_net_21563) );
na03f02 TIMEBOOST_cell_73798 ( .a(TIMEBOOST_net_12144), .b(n_13997), .c(FE_OFN1602_n_13995), .o(g53199_p) );
na03f02 TIMEBOOST_cell_68037 ( .a(FE_OFN1774_n_13800), .b(TIMEBOOST_net_13710), .c(FE_OFN1770_n_14054), .o(n_14447) );
in01f04 g54202_u0 ( .a(FE_OFN1084_n_13221), .o(g54202_sb) );
na03f01 TIMEBOOST_cell_64619 ( .a(n_12595), .b(FE_RN_578_0), .c(g54030_sb), .o(TIMEBOOST_net_17184) );
na03f02 TIMEBOOST_cell_72859 ( .a(TIMEBOOST_net_21744), .b(g64925_sb), .c(TIMEBOOST_net_21927), .o(TIMEBOOST_net_20959) );
in01f02 g54203_u0 ( .a(n_13221), .o(g54203_sb) );
na02s02 TIMEBOOST_cell_48767 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q), .b(g58357_sb), .o(TIMEBOOST_net_14601) );
na02s01 TIMEBOOST_cell_48901 ( .a(FE_OFN1648_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q), .o(TIMEBOOST_net_14668) );
na02f08 g74397_u0 ( .a(FE_OFN1069_n_15729), .b(configuration_wb_err_data_582), .o(n_15731) );
in01s01 TIMEBOOST_cell_63599 ( .a(TIMEBOOST_net_20779), .o(TIMEBOOST_net_20778) );
na03f02 TIMEBOOST_cell_65836 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(g64083_sb), .c(g64083_db), .o(n_4072) );
na02m06 TIMEBOOST_cell_69061 ( .a(TIMEBOOST_net_21738), .b(g64877_sb), .o(TIMEBOOST_net_12547) );
in01s02 g54205_u0 ( .a(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54205_sb) );
na03f08 TIMEBOOST_cell_33367 ( .a(n_7038), .b(n_4814), .c(n_16914), .o(TIMEBOOST_net_338) );
na02s02 TIMEBOOST_cell_53268 ( .a(TIMEBOOST_net_16851), .b(TIMEBOOST_net_11198), .o(TIMEBOOST_net_9578) );
na02s01 TIMEBOOST_cell_48739 ( .a(FE_OFN531_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q), .o(TIMEBOOST_net_14587) );
na02m02 TIMEBOOST_cell_43199 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q), .b(FE_OFN659_n_4392), .o(TIMEBOOST_net_12494) );
in01s02 g54207_u0 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54207_sb) );
na04f04 TIMEBOOST_cell_73494 ( .a(FE_OFN252_n_9868), .b(FE_OFN1670_n_9477), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q), .d(g58373_sb), .o(n_9456) );
na03f02 TIMEBOOST_cell_34797 ( .a(TIMEBOOST_net_9547), .b(FE_OFN1407_n_8567), .c(g57319_sb), .o(n_11432) );
na03m04 TIMEBOOST_cell_72762 ( .a(n_4452), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q), .c(TIMEBOOST_net_12758), .o(TIMEBOOST_net_20582) );
na03f02 TIMEBOOST_cell_73279 ( .a(TIMEBOOST_net_23317), .b(FE_OFN1166_n_5615), .c(g62140_sb), .o(n_5553) );
na03m02 TIMEBOOST_cell_69632 ( .a(FE_OFN640_n_4669), .b(n_4447), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q), .o(TIMEBOOST_net_22024) );
na03s02 TIMEBOOST_cell_41811 ( .a(n_1938), .b(g61797_sb), .c(g61797_db), .o(n_8203) );
in01s04 g54209_u0 ( .a(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54209_sb) );
na03f02 TIMEBOOST_cell_34907 ( .a(TIMEBOOST_net_9450), .b(FE_OFN1398_n_8567), .c(g57344_sb), .o(n_10391) );
na03f04 TIMEBOOST_cell_67068 ( .a(FE_OFN1768_n_14054), .b(TIMEBOOST_net_16550), .c(FE_OFN1775_n_13800), .o(n_14507) );
na02s01 TIMEBOOST_cell_51915 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q), .o(TIMEBOOST_net_16175) );
in01s01 TIMEBOOST_cell_31892 ( .a(TIMEBOOST_net_10056), .o(TIMEBOOST_net_10055) );
na03m02 TIMEBOOST_cell_42133 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q), .b(g58348_sb), .c(g58348_db), .o(n_9473) );
na02s01 TIMEBOOST_cell_39369 ( .a(TIMEBOOST_net_11296), .b(g58369_db), .o(n_9012) );
na03f02 TIMEBOOST_cell_65896 ( .a(TIMEBOOST_net_14912), .b(g63569_da), .c(g61961_sb), .o(TIMEBOOST_net_13028) );
na02m01 TIMEBOOST_cell_52381 ( .a(configuration_wb_err_cs_bit_568), .b(parchk_pci_cbe_out_in_1202), .o(TIMEBOOST_net_16408) );
na02f02 TIMEBOOST_cell_71118 ( .a(FE_OFN1265_n_4095), .b(TIMEBOOST_net_17419), .o(TIMEBOOST_net_22767) );
na02m02 TIMEBOOST_cell_47854 ( .a(TIMEBOOST_net_14144), .b(g57890_sb), .o(TIMEBOOST_net_10321) );
na04f04 TIMEBOOST_cell_34733 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q), .b(FE_OFN1373_n_8567), .c(n_9214), .d(g57470_sb), .o(n_10819) );
na02f01 TIMEBOOST_cell_47765 ( .a(pci_ad_i_16_), .b(FE_OFN989_n_574), .o(TIMEBOOST_net_14100) );
na02s01 TIMEBOOST_cell_50037 ( .a(wbm_adr_o_4_), .b(configuration_pci_err_addr_474), .o(TIMEBOOST_net_15236) );
na03f02 TIMEBOOST_cell_34478 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q), .b(g59796_sb), .c(g59796_db), .o(n_7621) );
na02s01 TIMEBOOST_cell_51916 ( .a(TIMEBOOST_net_16175), .b(FE_OFN1651_n_9428), .o(TIMEBOOST_net_10923) );
na02m02 TIMEBOOST_cell_39931 ( .a(TIMEBOOST_net_11577), .b(g62371_sb), .o(n_6861) );
in01s02 g54216_u0 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54216_sb) );
na02s01 g54216_u1 ( .a(g54216_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_404), .o(g54216_da) );
in01s01 TIMEBOOST_cell_31893 ( .a(TIMEBOOST_net_10057), .o(wbs_dat_i_9_) );
no02f10 TIMEBOOST_cell_68085 ( .a(TIMEBOOST_net_21250), .b(n_15210), .o(n_15729) );
na02m02 TIMEBOOST_cell_53060 ( .a(TIMEBOOST_net_16747), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_16447) );
in01s01 TIMEBOOST_cell_31894 ( .a(TIMEBOOST_net_10058), .o(TIMEBOOST_net_10057) );
in01s01 TIMEBOOST_cell_31895 ( .a(TIMEBOOST_net_10059), .o(wbs_dat_i_1_) );
in01s06 g54219_u0 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(g54219_sb) );
na02m02 TIMEBOOST_cell_52862 ( .a(TIMEBOOST_net_16648), .b(g58091_sb), .o(n_9706) );
na02f01 TIMEBOOST_cell_39410 ( .a(TIMEBOOST_net_8336), .b(FE_OFN2104_g64577_p), .o(TIMEBOOST_net_11317) );
na02m02 TIMEBOOST_cell_50038 ( .a(TIMEBOOST_net_15236), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_13317) );
na02s02 TIMEBOOST_cell_49728 ( .a(TIMEBOOST_net_15081), .b(g58286_db), .o(n_9517) );
na02m02 TIMEBOOST_cell_72041 ( .a(TIMEBOOST_net_23228), .b(TIMEBOOST_net_10646), .o(TIMEBOOST_net_17391) );
na03f01 TIMEBOOST_cell_72422 ( .a(TIMEBOOST_net_12285), .b(FE_OFN989_n_574), .c(g63590_sb), .o(n_1411) );
na03m02 TIMEBOOST_cell_69086 ( .a(g65058_sb), .b(n_4493), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q), .o(TIMEBOOST_net_21751) );
na02f02 TIMEBOOST_cell_70585 ( .a(TIMEBOOST_net_22500), .b(g63079_sb), .o(n_5094) );
na04m02 TIMEBOOST_cell_67852 ( .a(TIMEBOOST_net_14215), .b(FE_OFN654_n_4508), .c(g65327_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q), .o(TIMEBOOST_net_17364) );
na03f02 TIMEBOOST_cell_73667 ( .a(TIMEBOOST_net_20920), .b(FE_OFN1137_g64577_p), .c(g62767_sb), .o(n_5461) );
na03m02 TIMEBOOST_cell_65762 ( .a(TIMEBOOST_net_10921), .b(TIMEBOOST_net_8776), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q), .o(TIMEBOOST_net_17452) );
in01s01 TIMEBOOST_cell_31896 ( .a(TIMEBOOST_net_10060), .o(TIMEBOOST_net_10059) );
na02f01 TIMEBOOST_cell_68135 ( .a(TIMEBOOST_net_21275), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_393), .o(TIMEBOOST_net_16798) );
na02s01 TIMEBOOST_cell_64087 ( .a(TIMEBOOST_net_21029), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9366) );
na02s02 TIMEBOOST_cell_54735 ( .a(g58115_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_17585) );
na02s02 TIMEBOOST_cell_48158 ( .a(TIMEBOOST_net_14296), .b(g57949_sb), .o(TIMEBOOST_net_10516) );
na02s02 TIMEBOOST_cell_53472 ( .a(TIMEBOOST_net_16953), .b(g61800_sb), .o(n_8196) );
na02m10 TIMEBOOST_cell_45619 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q), .o(TIMEBOOST_net_13704) );
na03f02 TIMEBOOST_cell_35059 ( .a(TIMEBOOST_net_9592), .b(FE_OFN1441_n_9372), .c(g58463_sb), .o(n_9389) );
na02f02 TIMEBOOST_cell_72180 ( .a(TIMEBOOST_net_14886), .b(g64220_sb), .o(TIMEBOOST_net_23298) );
na03m02 TIMEBOOST_cell_65750 ( .a(TIMEBOOST_net_20365), .b(n_4517), .c(g61947_sb), .o(n_7931) );
na03m02 TIMEBOOST_cell_72895 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q), .b(g64292_sb), .c(TIMEBOOST_net_22096), .o(TIMEBOOST_net_13038) );
na02s01 TIMEBOOST_cell_50730 ( .a(TIMEBOOST_net_15582), .b(TIMEBOOST_net_10583), .o(TIMEBOOST_net_9440) );
na04f04 TIMEBOOST_cell_24203 ( .a(n_9011), .b(g57511_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q), .d(FE_OFN1405_n_8567), .o(n_10321) );
na04m06 TIMEBOOST_cell_72757 ( .a(g64926_sb), .b(n_4447), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q), .d(g64926_db), .o(TIMEBOOST_net_17543) );
in01s01 TIMEBOOST_cell_31897 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .o(TIMEBOOST_net_10061) );
na02m01 TIMEBOOST_cell_47655 ( .a(FE_OFN2054_n_8831), .b(wbu_addr_in), .o(TIMEBOOST_net_14045) );
na02m01 TIMEBOOST_cell_37950 ( .a(FE_OFN1663_n_4490), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_10587) );
na03m02 TIMEBOOST_cell_65954 ( .a(TIMEBOOST_net_20435), .b(FE_OFN1166_n_5615), .c(g62135_sb), .o(n_5558) );
na04m02 TIMEBOOST_cell_72758 ( .a(FE_OFN653_n_4508), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q), .c(n_4645), .d(g65430_sb), .o(n_4222) );
na02m02 TIMEBOOST_cell_71981 ( .a(TIMEBOOST_net_23198), .b(TIMEBOOST_net_16273), .o(TIMEBOOST_net_17566) );
na02f02 TIMEBOOST_cell_49870 ( .a(TIMEBOOST_net_15152), .b(g62849_sb), .o(n_5272) );
na03f02 TIMEBOOST_cell_73746 ( .a(FE_OFN1756_n_12681), .b(TIMEBOOST_net_13671), .c(FE_OCP_RBN1976_n_12381), .o(n_12638) );
in01f02 g54234_u0 ( .a(FE_OFN1148_n_13249), .o(g54234_sb) );
na03m02 TIMEBOOST_cell_65394 ( .a(wbs_sel_i_3_), .b(g63586_sb), .c(g63587_db), .o(n_4101) );
na02m01 TIMEBOOST_cell_62828 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_132), .o(TIMEBOOST_net_20361) );
in01f02 g54235_u0 ( .a(FE_OFN1150_n_13249), .o(g54235_sb) );
in01s01 TIMEBOOST_cell_73835 ( .a(TIMEBOOST_net_23399), .o(TIMEBOOST_net_23400) );
na02s04 TIMEBOOST_cell_52623 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q), .o(TIMEBOOST_net_16529) );
na02f02 g59231_u2 ( .a(n_3478), .b(FE_OFN1697_n_5751), .o(g59231_db) );
in01f02 g54236_u0 ( .a(FE_OFN1151_n_13249), .o(g54236_sb) );
na04f04 TIMEBOOST_cell_34996 ( .a(n_9059), .b(g57325_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q), .d(FE_OFN1380_n_8567), .o(n_10399) );
na02f01 TIMEBOOST_cell_69774 ( .a(pci_target_unit_del_sync_bc_in_202), .b(g65940_sb), .o(TIMEBOOST_net_22095) );
in01f04 g54237_u0 ( .a(FE_OCPN1911_FE_OFN1152_n_13249), .o(g54237_sb) );
na02f01 TIMEBOOST_cell_26069 ( .a(pci_target_unit_pcit_if_strd_addr_in_715), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_7139) );
na02s02 TIMEBOOST_cell_47867 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q), .b(g65878_sb), .o(TIMEBOOST_net_14151) );
na02f02 TIMEBOOST_cell_54275 ( .a(n_2486), .b(FE_OFN1698_n_5751), .o(TIMEBOOST_net_17355) );
in01f02 g54238_u0 ( .a(FE_OFN1149_n_13249), .o(g54238_sb) );
na02m01 TIMEBOOST_cell_69742 ( .a(n_4444), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q), .o(TIMEBOOST_net_22079) );
in01f02 g54239_u0 ( .a(FE_OFN1150_n_13249), .o(g54239_sb) );
na02s01 TIMEBOOST_cell_68215 ( .a(TIMEBOOST_net_21315), .b(g66427_db), .o(n_3000) );
na02s01 TIMEBOOST_cell_48919 ( .a(FE_OFN1649_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q), .o(TIMEBOOST_net_14677) );
in01f02 g54244_u0 ( .a(FE_OFN1306_n_13124), .o(g54244_sb) );
na03s02 TIMEBOOST_cell_41722 ( .a(g58320_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q), .c(g58320_db), .o(n_9024) );
na03f02 TIMEBOOST_cell_68039 ( .a(FE_OFN1774_n_13800), .b(TIMEBOOST_net_13705), .c(FE_OFN1771_n_14054), .o(n_14477) );
na03f02 TIMEBOOST_cell_65950 ( .a(TIMEBOOST_net_20439), .b(FE_OFN1170_n_5592), .c(g62125_sb), .o(n_5571) );
na02f02 g54265_u0 ( .a(n_13410), .b(wbm_cti_o_0_), .o(n_13412) );
na02f02 g54266_u0 ( .a(n_13410), .b(wbm_cti_o_2_), .o(n_13411) );
no02f04 g54267_u0 ( .a(n_13486), .b(n_8757), .o(n_13624) );
na02f02 g54269_u0 ( .a(n_13317), .b(n_13068), .o(n_13409) );
na02f02 g54271_u0 ( .a(n_13315), .b(n_12963), .o(n_13407) );
na02f02 g54273_u0 ( .a(n_13063), .b(n_13314), .o(n_13406) );
na02f02 g54274_u0 ( .a(n_13313), .b(n_13066), .o(n_13405) );
na02f02 g54283_u0 ( .a(n_16413), .b(n_13056), .o(n_13404) );
na02f02 g54289_u0 ( .a(n_13311), .b(n_12958), .o(n_13403) );
na02f02 g54290_u0 ( .a(n_13310), .b(n_13052), .o(n_13402) );
oa12f02 g54294_u0 ( .a(n_13620), .b(n_13621), .c(pci_target_unit_fifos_pciw_outTransactionCount_1_), .o(n_13623) );
oa12f02 g54295_u0 ( .a(n_13620), .b(n_13621), .c(pci_target_unit_fifos_outGreyCount_0_), .o(n_13622) );
na02f02 g54297_u0 ( .a(n_13309), .b(n_13048), .o(n_13401) );
na02f02 g54298_u0 ( .a(n_13308), .b(n_13047), .o(n_13400) );
na02f02 g54303_u0 ( .a(n_16401), .b(n_13042), .o(n_13399) );
in01f04 g54304_u0 ( .a(FE_OFN2128_n_16497), .o(g54304_sb) );
in01s01 TIMEBOOST_cell_63581 ( .a(TIMEBOOST_net_20760), .o(TIMEBOOST_net_20761) );
na02f01 TIMEBOOST_cell_29021 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q), .o(TIMEBOOST_net_8615) );
in01f02 g54305_u0 ( .a(FE_OFN2128_n_16497), .o(g54305_sb) );
na03m02 TIMEBOOST_cell_72778 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q), .c(TIMEBOOST_net_16327), .o(TIMEBOOST_net_17582) );
na02s01 TIMEBOOST_cell_42799 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q), .o(TIMEBOOST_net_12294) );
in01f02 g54306_u0 ( .a(FE_OFN2128_n_16497), .o(g54306_sb) );
na02f02 TIMEBOOST_cell_28209 ( .a(FE_RN_602_0), .b(FE_RN_593_0), .o(TIMEBOOST_net_8209) );
na02s02 TIMEBOOST_cell_63015 ( .a(TIMEBOOST_net_20454), .b(g58219_db), .o(TIMEBOOST_net_9332) );
na02f02 TIMEBOOST_cell_28210 ( .a(TIMEBOOST_net_8209), .b(FE_RN_606_0), .o(TIMEBOOST_net_319) );
ao12f02 g54308_u0 ( .a(n_13073), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q), .c(FE_OCPN1909_n_16497), .o(n_13127) );
in01f01 g54309_u0 ( .a(FE_OFN2128_n_16497), .o(g54309_sb) );
na03f02 TIMEBOOST_cell_66523 ( .a(g53916_sb), .b(FE_OFN1326_n_13547), .c(TIMEBOOST_net_16803), .o(n_13526) );
in01f02 g54310_u0 ( .a(FE_OFN2128_n_16497), .o(g54310_sb) );
na02s02 TIMEBOOST_cell_70035 ( .a(TIMEBOOST_net_22225), .b(g61830_sb), .o(n_8125) );
in01f04 g54311_u0 ( .a(FE_OFN2126_n_16497), .o(g54311_sb) );
na02f02 g54311_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q), .b(FE_OFN2126_n_16497), .o(g54311_db) );
na03f02 TIMEBOOST_cell_34924 ( .a(TIMEBOOST_net_9494), .b(FE_OFN1401_n_8567), .c(g57197_sb), .o(n_11556) );
in01f01 g54312_u0 ( .a(FE_OFN2127_n_16497), .o(g54312_sb) );
na03f01 TIMEBOOST_cell_47370 ( .a(FE_OFN1579_n_12306), .b(TIMEBOOST_net_13680), .c(FE_OFN1760_n_10780), .o(n_12667) );
na02s01 TIMEBOOST_cell_49729 ( .a(FE_OFN1793_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q), .o(TIMEBOOST_net_15082) );
in01f01 g54314_u0 ( .a(FE_OFN2126_n_16497), .o(g54314_sb) );
na03f04 TIMEBOOST_cell_73482 ( .a(wbm_adr_o_17_), .b(g59230_sb), .c(g52393_sb), .o(TIMEBOOST_net_15659) );
na02m10 TIMEBOOST_cell_52957 ( .a(wishbone_slave_unit_pcim_sm_data_in_644), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q), .o(TIMEBOOST_net_16696) );
in01f01 g54315_u0 ( .a(FE_OFN2126_n_16497), .o(g54315_sb) );
na02m20 TIMEBOOST_cell_42713 ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .b(g54160_sb), .o(TIMEBOOST_net_12251) );
na02f02 g54315_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q), .b(FE_OFN2125_n_16497), .o(g54315_db) );
na02m04 TIMEBOOST_cell_62604 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q), .b(n_3755), .o(TIMEBOOST_net_20249) );
in01f01 g54316_u0 ( .a(FE_OCPN1909_n_16497), .o(g54316_sb) );
na02m01 TIMEBOOST_cell_68642 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q), .b(FE_OFN667_n_4495), .o(TIMEBOOST_net_21529) );
in01f01 g54317_u0 ( .a(FE_OFN2127_n_16497), .o(g54317_sb) );
na04f04 TIMEBOOST_cell_34998 ( .a(n_9071), .b(g57272_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q), .d(FE_OFN1412_n_8567), .o(n_10414) );
na02s01 TIMEBOOST_cell_37624 ( .a(FE_OFN217_n_9889), .b(g57984_sb), .o(TIMEBOOST_net_10424) );
na02m02 TIMEBOOST_cell_54559 ( .a(n_1852), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q), .o(TIMEBOOST_net_17497) );
in01f01 g54318_u0 ( .a(FE_OFN2127_n_16497), .o(g54318_sb) );
na02f08 TIMEBOOST_cell_47716 ( .a(TIMEBOOST_net_14075), .b(n_1619), .o(TIMEBOOST_net_363) );
in01s01 TIMEBOOST_cell_45966 ( .a(TIMEBOOST_net_13926), .o(TIMEBOOST_net_13927) );
na02s02 TIMEBOOST_cell_48783 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q), .b(g58372_sb), .o(TIMEBOOST_net_14609) );
in01f01 g54319_u0 ( .a(FE_OCPN1909_n_16497), .o(g54319_sb) );
na03m04 TIMEBOOST_cell_73206 ( .a(TIMEBOOST_net_23231), .b(g65836_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q), .o(TIMEBOOST_net_22373) );
na02s01 TIMEBOOST_cell_47518 ( .a(TIMEBOOST_net_13976), .b(g67042_sb), .o(n_1276) );
in01f01 g54320_u0 ( .a(FE_OCPN1909_n_16497), .o(g54320_sb) );
na02m06 TIMEBOOST_cell_43489 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q), .o(TIMEBOOST_net_12639) );
na02s01 TIMEBOOST_cell_47519 ( .a(parchk_pci_ad_reg_in_1215), .b(g67075_db), .o(TIMEBOOST_net_13977) );
in01f04 g54321_u0 ( .a(FE_OCPN1909_n_16497), .o(g54321_sb) );
in01s02 TIMEBOOST_cell_45968 ( .a(TIMEBOOST_net_13928), .o(TIMEBOOST_net_13929) );
na02m02 TIMEBOOST_cell_69693 ( .a(TIMEBOOST_net_22054), .b(g65383_sb), .o(TIMEBOOST_net_16327) );
in01f02 g54322_u0 ( .a(FE_OCPN1909_n_16497), .o(g54322_sb) );
na02f02 TIMEBOOST_cell_71002 ( .a(TIMEBOOST_net_13248), .b(FE_OFN1226_n_6391), .o(TIMEBOOST_net_22709) );
in01s01 TIMEBOOST_cell_45970 ( .a(TIMEBOOST_net_13930), .o(TIMEBOOST_net_13931) );
no02f10 FE_RC_830_0 ( .a(FE_RN_538_0), .b(FE_RN_539_0), .o(FE_RN_540_0) );
in01f01 g54323_u0 ( .a(FE_OFN2127_n_16497), .o(g54323_sb) );
na04f04 TIMEBOOST_cell_24650 ( .a(n_9705), .b(g57232_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q), .d(FE_OFN2174_n_8567), .o(n_11523) );
na04f04 TIMEBOOST_cell_73044 ( .a(n_1595), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q), .c(FE_OFN714_n_8140), .d(g61806_sb), .o(n_8182) );
in01f02 g54324_u0 ( .a(FE_OCPN1909_n_16497), .o(g54324_sb) );
na02m02 TIMEBOOST_cell_68716 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q), .b(n_3747), .o(TIMEBOOST_net_21566) );
in01s01 TIMEBOOST_cell_45972 ( .a(TIMEBOOST_net_13932), .o(TIMEBOOST_net_13933) );
in01f01 g54325_u0 ( .a(FE_OFN2125_n_16497), .o(g54325_sb) );
na03f02 TIMEBOOST_cell_65952 ( .a(TIMEBOOST_net_17309), .b(FE_OFN1171_n_5592), .c(g62128_sb), .o(n_5568) );
na02s01 TIMEBOOST_cell_45373 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q), .o(TIMEBOOST_net_13581) );
in01f01 g54326_u0 ( .a(FE_OFN2127_n_16497), .o(g54326_sb) );
na02m01 TIMEBOOST_cell_68553 ( .a(TIMEBOOST_net_21484), .b(FE_OFN2071_n_15978), .o(TIMEBOOST_net_20612) );
na04f04 TIMEBOOST_cell_24652 ( .a(n_9708), .b(g57229_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q), .d(FE_OFN2177_n_8567), .o(n_11526) );
na03f02 TIMEBOOST_cell_73593 ( .a(TIMEBOOST_net_17530), .b(FE_OFN2064_n_6391), .c(g62441_sb), .o(n_6714) );
in01f02 g54328_u0 ( .a(FE_OFN2126_n_16497), .o(g54328_sb) );
na04f04 TIMEBOOST_cell_24840 ( .a(wbs_dat_o_13_), .b(g52507_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_112), .d(FE_OFN2243_g52675_p), .o(n_13719) );
na02m04 TIMEBOOST_cell_71890 ( .a(n_3739), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q), .o(TIMEBOOST_net_23153) );
no02f02 g54329_u0 ( .a(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q), .b(n_13621), .o(g54329_p) );
ao12f01 g54329_u1 ( .a(g54329_p), .b(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q), .c(n_13621), .o(n_13483) );
in01f02 g54330_u0 ( .a(FE_OCPN1909_n_16497), .o(g54330_sb) );
no04f08 TIMEBOOST_cell_21033 ( .a(FE_RN_647_0), .b(FE_RN_659_0), .c(FE_RN_665_0), .d(FE_RN_653_0), .o(FE_RN_666_0) );
na02m02 TIMEBOOST_cell_68398 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(g64190_sb), .o(TIMEBOOST_net_21407) );
na03f02 TIMEBOOST_cell_66947 ( .a(FE_OFN1751_n_12086), .b(FE_OFN1572_n_11027), .c(TIMEBOOST_net_13610), .o(n_12670) );
in01f02 g54331_u0 ( .a(FE_OFN2126_n_16497), .o(g54331_sb) );
no02f10 TIMEBOOST_cell_42695 ( .a(conf_wb_err_bc_in), .b(conf_wb_err_bc_in_846), .o(TIMEBOOST_net_12242) );
na02s01 TIMEBOOST_cell_42721 ( .a(pci_ad_i_22_), .b(parchk_pci_ad_reg_in_1226), .o(TIMEBOOST_net_12255) );
in01f02 g54332_u0 ( .a(FE_OFN2128_n_16497), .o(g54332_sb) );
na03f02 TIMEBOOST_cell_66527 ( .a(g53911_sb), .b(FE_OFN1327_n_13547), .c(TIMEBOOST_net_16793), .o(n_13530) );
na02m02 TIMEBOOST_cell_69568 ( .a(TIMEBOOST_net_14204), .b(FE_OFN917_n_4725), .o(TIMEBOOST_net_21992) );
in01f06 g54333_u0 ( .a(FE_OFN2128_n_16497), .o(g54333_sb) );
na02f02 TIMEBOOST_cell_71033 ( .a(TIMEBOOST_net_22724), .b(g62545_sb), .o(n_6477) );
na04f02 TIMEBOOST_cell_67949 ( .a(n_4722), .b(n_384), .c(FE_OFN1127_g64577_p), .d(g63044_sb), .o(n_7123) );
na02m04 TIMEBOOST_cell_68580 ( .a(FE_OFN629_n_4454), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q), .o(TIMEBOOST_net_21498) );
in01f01 g54334_u0 ( .a(FE_OFN2128_n_16497), .o(g54334_sb) );
na02s01 TIMEBOOST_cell_47520 ( .a(TIMEBOOST_net_13977), .b(g67049_sb), .o(n_1429) );
na02f01 TIMEBOOST_cell_48612 ( .a(TIMEBOOST_net_14523), .b(g65249_sb), .o(n_2633) );
na03f02 TIMEBOOST_cell_66949 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_16500), .c(FE_OFN2210_n_11027), .o(n_12717) );
in01f02 g54335_u0 ( .a(FE_OFN2126_n_16497), .o(g54335_sb) );
na03f02 TIMEBOOST_cell_34854 ( .a(TIMEBOOST_net_9422), .b(FE_OFN1385_n_8567), .c(g57359_sb), .o(n_11388) );
in01f01 g54336_u0 ( .a(FE_OFN2128_n_16497), .o(g54336_sb) );
na02m02 TIMEBOOST_cell_72328 ( .a(g64766_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q), .o(TIMEBOOST_net_23372) );
na02m10 TIMEBOOST_cell_52959 ( .a(wishbone_slave_unit_pcim_sm_data_in_658), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q), .o(TIMEBOOST_net_16697) );
in01f02 g54337_u0 ( .a(n_13621), .o(g54337_sb) );
na02m10 TIMEBOOST_cell_45639 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q), .o(TIMEBOOST_net_13714) );
in01f02 g54338_u0 ( .a(FE_OFN1305_n_13124), .o(g54338_sb) );
na04m02 TIMEBOOST_cell_72542 ( .a(TIMEBOOST_net_14170), .b(FE_OFN916_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q), .d(g64356_sb), .o(TIMEBOOST_net_20472) );
na02m02 TIMEBOOST_cell_69127 ( .a(TIMEBOOST_net_21771), .b(g65326_sb), .o(TIMEBOOST_net_12543) );
in01f02 g54339_u0 ( .a(FE_OFN2136_n_13124), .o(g54339_sb) );
in01s01 TIMEBOOST_cell_73836 ( .a(n_11855), .o(TIMEBOOST_net_23401) );
na03m04 TIMEBOOST_cell_72478 ( .a(TIMEBOOST_net_20176), .b(FE_OFN905_n_4736), .c(g64102_sb), .o(TIMEBOOST_net_9945) );
na02s01 g61989_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61989_db) );
in01f02 g54340_u0 ( .a(FE_OFN2134_n_13124), .o(g54340_sb) );
na02f02 TIMEBOOST_cell_72305 ( .a(TIMEBOOST_net_23360), .b(TIMEBOOST_net_14977), .o(TIMEBOOST_net_9382) );
na02m02 TIMEBOOST_cell_43089 ( .a(n_3739), .b(n_4669), .o(TIMEBOOST_net_12439) );
in01s01 TIMEBOOST_cell_31898 ( .a(TIMEBOOST_net_10061), .o(TIMEBOOST_net_10062) );
in01f02 g54341_u0 ( .a(FE_OFN2134_n_13124), .o(g54341_sb) );
na03m04 TIMEBOOST_cell_72978 ( .a(g64942_sb), .b(n_3672), .c(TIMEBOOST_net_14559), .o(TIMEBOOST_net_13362) );
na04f02 TIMEBOOST_cell_36823 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q), .b(FE_OFN1394_n_8567), .c(n_8562), .d(g58586_sb), .o(n_8959) );
in01f02 g54342_u0 ( .a(FE_OFN2134_n_13124), .o(g54342_sb) );
na04m04 TIMEBOOST_cell_73045 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q), .b(FE_OFN704_n_8069), .c(n_2200), .d(g61719_sb), .o(n_8387) );
in01s01 TIMEBOOST_cell_31899 ( .a(TIMEBOOST_net_10063), .o(wbs_adr_i_0_) );
in01f02 g54343_u0 ( .a(FE_OFN2136_n_13124), .o(g54343_sb) );
na04f02 TIMEBOOST_cell_72546 ( .a(g58768_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q), .c(n_8884), .d(wbu_addr_in_259), .o(n_9862) );
na02m08 TIMEBOOST_cell_52873 ( .a(wbs_dat_i_30_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q), .o(TIMEBOOST_net_16654) );
in01f02 g54344_u0 ( .a(FE_OFN2134_n_13124), .o(g54344_sb) );
na02m10 TIMEBOOST_cell_72030 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_23223) );
na02s02 TIMEBOOST_cell_28242 ( .a(TIMEBOOST_net_8225), .b(g65761_sb), .o(n_1919) );
na02s01 TIMEBOOST_cell_4086 ( .a(g61880_sb), .b(g61983_db), .o(TIMEBOOST_net_603) );
in01f02 g54345_u0 ( .a(FE_OFN2134_n_13124), .o(g54345_sb) );
na02m08 TIMEBOOST_cell_72032 ( .a(g65404_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q), .o(TIMEBOOST_net_23224) );
na02f02 TIMEBOOST_cell_50514 ( .a(TIMEBOOST_net_15474), .b(g62524_sb), .o(n_6528) );
na02m20 TIMEBOOST_cell_52837 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69), .b(pci_target_unit_pcit_if_strd_addr_in_705), .o(TIMEBOOST_net_16636) );
in01f02 g54346_u0 ( .a(FE_OFN2134_n_13124), .o(g54346_sb) );
na02f02 TIMEBOOST_cell_70028 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q), .b(FE_OFN2256_n_8060), .o(TIMEBOOST_net_22222) );
in01f02 g54347_u0 ( .a(FE_OFN2134_n_13124), .o(g54347_sb) );
na02s01 TIMEBOOST_cell_28246 ( .a(TIMEBOOST_net_8227), .b(g58033_db), .o(n_9098) );
na03s02 TIMEBOOST_cell_72903 ( .a(n_1657), .b(g61934_sb), .c(g61934_db), .o(n_7955) );
in01f02 g54348_u0 ( .a(FE_OFN2135_n_13124), .o(g54348_sb) );
na04m02 TIMEBOOST_cell_73046 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q), .b(FE_OFN702_n_7845), .c(n_2186), .d(g62002_sb), .o(n_7891) );
na04m04 TIMEBOOST_cell_65104 ( .a(g65388_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q), .c(FE_OFN639_n_4669), .d(n_4442), .o(TIMEBOOST_net_7548) );
na02s01 g61962_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61962_db) );
in01f02 g54349_u0 ( .a(FE_OFN1306_n_13124), .o(g54349_sb) );
na03f02 TIMEBOOST_cell_73534 ( .a(TIMEBOOST_net_17503), .b(FE_OFN1230_n_6391), .c(g62379_sb), .o(n_6845) );
na04f04 TIMEBOOST_cell_73280 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q), .b(FE_OFN1106_g64577_p), .c(n_3930), .d(g62835_sb), .o(n_5196) );
in01f02 g54350_u0 ( .a(FE_OFN2134_n_13124), .o(g54350_sb) );
na04f02 TIMEBOOST_cell_36859 ( .a(TIMEBOOST_net_10023), .b(g52621_sb), .c(n_2257), .d(n_10256), .o(n_11848) );
na02f02 TIMEBOOST_cell_70457 ( .a(TIMEBOOST_net_22436), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_11420) );
na02s01 TIMEBOOST_cell_62423 ( .a(TIMEBOOST_net_20158), .b(g58042_sb), .o(TIMEBOOST_net_14259) );
in01f02 g54351_u0 ( .a(FE_OFN2134_n_13124), .o(g54351_sb) );
na04f04 TIMEBOOST_cell_36855 ( .a(n_2924), .b(n_2868), .c(n_3054), .d(n_2867), .o(n_4171) );
na02f02 TIMEBOOST_cell_54650 ( .a(TIMEBOOST_net_17542), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_15487) );
na02f01 TIMEBOOST_cell_4096 ( .a(n_6986), .b(g59226_da), .o(TIMEBOOST_net_608) );
in01f02 g54352_u0 ( .a(FE_OFN2135_n_13124), .o(g54352_sb) );
na03m02 TIMEBOOST_cell_72881 ( .a(g61864_sb), .b(g61864_db), .c(n_1845), .o(n_8109) );
na02f02 TIMEBOOST_cell_4097 ( .a(TIMEBOOST_net_608), .b(n_4202), .o(n_5748) );
na02f02 TIMEBOOST_cell_4098 ( .a(n_7622), .b(n_16914), .o(TIMEBOOST_net_609) );
in01f02 g54353_u0 ( .a(FE_OFN1305_n_13124), .o(g54353_sb) );
na02s02 TIMEBOOST_cell_72056 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(FE_OFN1017_n_2053), .o(TIMEBOOST_net_23236) );
na02s01 TIMEBOOST_cell_37625 ( .a(TIMEBOOST_net_10424), .b(g57984_db), .o(n_9814) );
na02f02 TIMEBOOST_cell_54671 ( .a(n_4480), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q), .o(TIMEBOOST_net_17553) );
in01f02 g54354_u0 ( .a(FE_OFN1305_n_13124), .o(g54354_sb) );
na02f01 TIMEBOOST_cell_44406 ( .a(TIMEBOOST_net_13097), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_11298) );
in01f02 g54355_u0 ( .a(FE_OFN2136_n_13124), .o(g54355_sb) );
na02s01 TIMEBOOST_cell_42893 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q), .o(TIMEBOOST_net_12341) );
na03f02 TIMEBOOST_cell_69398 ( .a(n_4479), .b(g64952_db), .c(n_74), .o(TIMEBOOST_net_21907) );
na02f01 TIMEBOOST_cell_69309 ( .a(TIMEBOOST_net_21862), .b(FE_OFN1810_n_4454), .o(TIMEBOOST_net_14680) );
in01f02 g54356_u0 ( .a(FE_OFN2136_n_13124), .o(g54356_sb) );
na02m01 TIMEBOOST_cell_42871 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q), .b(pci_target_unit_fifos_pciw_cbe_in_152), .o(TIMEBOOST_net_12330) );
na02f02 TIMEBOOST_cell_70777 ( .a(TIMEBOOST_net_22596), .b(g63576_sb), .o(TIMEBOOST_net_20992) );
in01f02 g54357_u0 ( .a(FE_OFN1306_n_13124), .o(g54357_sb) );
na03f02 TIMEBOOST_cell_66951 ( .a(FE_OFN1753_n_12086), .b(FE_OFN1568_n_11027), .c(TIMEBOOST_net_13620), .o(n_12641) );
na04m04 TIMEBOOST_cell_67188 ( .a(g65038_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q), .c(n_4479), .d(FE_OFN633_n_4454), .o(n_4330) );
in01f02 g54358_u0 ( .a(FE_OFN1305_n_13124), .o(g54358_sb) );
na02m02 TIMEBOOST_cell_72064 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q), .o(TIMEBOOST_net_23240) );
na03m02 TIMEBOOST_cell_73148 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(g64133_sb), .c(TIMEBOOST_net_7320), .o(n_4029) );
in01f02 g54359_u0 ( .a(FE_OFN1306_n_13124), .o(g54359_sb) );
na03m02 TIMEBOOST_cell_72786 ( .a(n_4498), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q), .c(TIMEBOOST_net_12685), .o(TIMEBOOST_net_17374) );
in01f02 g54360_u0 ( .a(FE_OFN1306_n_13124), .o(g54360_sb) );
na03m02 TIMEBOOST_cell_72058 ( .a(n_4482), .b(FE_OFN1642_n_4671), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q), .o(TIMEBOOST_net_23237) );
na02s02 TIMEBOOST_cell_37685 ( .a(TIMEBOOST_net_10454), .b(g65767_sb), .o(n_1915) );
na02m02 TIMEBOOST_cell_44255 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q), .b(g58271_sb), .o(TIMEBOOST_net_13022) );
in01f02 g54361_u0 ( .a(FE_OFN1306_n_13124), .o(g54361_sb) );
in01f02 g54362_u0 ( .a(FE_OFN1305_n_13124), .o(g54362_sb) );
na02m04 TIMEBOOST_cell_69734 ( .a(FE_OFN1678_n_4655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q), .o(TIMEBOOST_net_22075) );
na02s01 TIMEBOOST_cell_70256 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_22336) );
in01f02 g54363_u0 ( .a(FE_OFN1306_n_13124), .o(g54363_sb) );
na03m06 TIMEBOOST_cell_72072 ( .a(TIMEBOOST_net_16934), .b(FE_OFN1055_n_4727), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q), .o(TIMEBOOST_net_23244) );
na02f02 TIMEBOOST_cell_70617 ( .a(TIMEBOOST_net_22516), .b(g63083_sb), .o(n_5088) );
na02s02 TIMEBOOST_cell_4044 ( .a(n_1798), .b(n_3341), .o(TIMEBOOST_net_582) );
in01f01 g54364_u0 ( .a(FE_OFN1305_n_13124), .o(g54364_sb) );
na04f04 TIMEBOOST_cell_35000 ( .a(n_9001), .b(g57548_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q), .d(FE_OFN1412_n_8567), .o(n_10304) );
na02s01 TIMEBOOST_cell_52625 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_16530) );
in01f02 g54365_u0 ( .a(FE_OFN1306_n_13124), .o(g54365_sb) );
na02s01 TIMEBOOST_cell_45433 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_13611) );
na04f04 TIMEBOOST_cell_24649 ( .a(n_9221), .b(g57234_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q), .d(FE_OFN2178_n_8567), .o(n_10833) );
in01f02 g54366_u0 ( .a(FE_OFN1305_n_13124), .o(g54366_sb) );
na03m02 TIMEBOOST_cell_71346 ( .a(n_2054), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q), .c(FE_OFN701_n_7845), .o(TIMEBOOST_net_22881) );
no02f06 TIMEBOOST_cell_4046 ( .a(FE_RN_159_0), .b(FE_RN_160_0), .o(TIMEBOOST_net_583) );
in01f02 g54367_u0 ( .a(FE_OFN1305_n_13124), .o(g54367_sb) );
na04f04 TIMEBOOST_cell_73070 ( .a(n_1590), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q), .c(FE_OFN714_n_8140), .d(g61803_sb), .o(n_8189) );
na03f02 TIMEBOOST_cell_34856 ( .a(TIMEBOOST_net_9471), .b(FE_OFN1382_n_8567), .c(g57368_sb), .o(n_10381) );
na02s01 TIMEBOOST_cell_4050 ( .a(FE_OCPN1875_n_14526), .b(n_16451), .o(TIMEBOOST_net_585) );
in01f02 g54368_u0 ( .a(FE_OFN2135_n_13124), .o(g54368_sb) );
na02m02 TIMEBOOST_cell_68655 ( .a(TIMEBOOST_net_21535), .b(g65671_db), .o(TIMEBOOST_net_16764) );
na03f02 TIMEBOOST_cell_66878 ( .a(FE_OFN1564_n_12502), .b(TIMEBOOST_net_15983), .c(n_12313), .o(n_12648) );
in01f02 g54369_u0 ( .a(FE_OFN2135_n_13124), .o(g54369_sb) );
na02m01 TIMEBOOST_cell_69046 ( .a(n_95), .b(FE_OFN620_n_4490), .o(TIMEBOOST_net_21731) );
na02s01 TIMEBOOST_cell_47768 ( .a(TIMEBOOST_net_14101), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_394), .o(n_13184) );
na03s02 TIMEBOOST_cell_72548 ( .a(FE_OFN551_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q), .c(TIMEBOOST_net_20820), .o(TIMEBOOST_net_14972) );
no02f02 g54408_u0 ( .a(n_13041), .b(n_12759), .o(n_13317) );
no02f02 g54410_u0 ( .a(n_17028), .b(n_17029), .o(n_13315) );
no02f02 g54411_u0 ( .a(n_16600), .b(n_16601), .o(n_13314) );
no02f02 g54412_u0 ( .a(n_16602), .b(n_16603), .o(n_13313) );
no02f02 g54414_u0 ( .a(n_15440), .b(n_15441), .o(n_13311) );
no02f02 g54415_u0 ( .a(n_16588), .b(n_16589), .o(n_13310) );
no02f02 g54416_u0 ( .a(n_15438), .b(n_15439), .o(n_13309) );
no02f02 g54417_u0 ( .a(n_16591), .b(n_16592), .o(n_13308) );
na02f06 g54419_u0 ( .a(n_998), .b(n_13621), .o(n_13620) );
na02f02 g54420_u0 ( .a(FE_OFN2163_n_16301), .b(wbm_dat_o_0_), .o(n_13398) );
na02f02 g54422_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_11_), .o(n_13395) );
na02f02 g54423_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_12_), .o(n_13394) );
na02f02 g54424_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_13_), .o(n_13393) );
na02f02 g54425_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_14_), .o(n_13392) );
na02f02 g54426_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_15_), .o(n_13391) );
na02f02 g54427_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_16_), .o(n_13390) );
na02f02 g54428_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_17_), .o(n_13389) );
na02f02 g54429_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_18_), .o(n_13388) );
na02f02 g54430_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_19_), .o(n_13387) );
na02f02 g54431_u0 ( .a(FE_OFN2163_n_16301), .b(wbm_dat_o_1_), .o(n_13386) );
na02f02 g54432_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_20_), .o(n_13384) );
na02f02 g54433_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_21_), .o(n_13383) );
na02f02 g54435_u0 ( .a(FE_OFN2165_n_16301), .b(wbm_dat_o_23_), .o(n_13381) );
na02f02 g54436_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_24_), .o(n_13380) );
na02f02 g54437_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_25_), .o(n_13379) );
na02f02 g54438_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_26_), .o(n_13378) );
na02f02 g54439_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_27_), .o(n_13377) );
na02f02 g54440_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_28_), .o(n_13376) );
na02f02 g54441_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_29_), .o(n_13375) );
na02f02 g54442_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_2_), .o(n_13374) );
na02f02 g54443_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_30_), .o(n_13373) );
na02f02 g54444_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_31_), .o(n_13372) );
na02f02 g54445_u0 ( .a(FE_OFN2163_n_16301), .b(wbm_dat_o_3_), .o(n_13371) );
na02f02 g54446_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_4_), .o(n_13370) );
na02f02 g54447_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_5_), .o(n_13369) );
na02f02 g54448_u0 ( .a(FE_OFN2162_n_16301), .b(wbm_dat_o_6_), .o(n_13368) );
na02f02 g54449_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_7_), .o(n_13367) );
na02f02 g54450_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_8_), .o(n_13366) );
na02f02 g54451_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_9_), .o(n_13365) );
no02f02 g54452_u0 ( .a(n_12952), .b(FE_OCPN1909_n_16497), .o(n_13073) );
na02f02 g54453_u0 ( .a(n_16495), .b(pci_target_unit_pcit_if_pcir_fifo_control_in_637), .o(g54453_p) );
in01f02 g54453_u1 ( .a(g54453_p), .o(n_13145) );
in01f03 g54454_u0 ( .a(n_13410), .o(n_14518) );
no02f02 g54456_u0 ( .a(n_16299), .b(n_13122), .o(g54456_p) );
in01f02 g54456_u1 ( .a(g54456_p), .o(n_14898) );
no02f06 g54457_u0 ( .a(FE_OFN1705_n_4868), .b(n_13721), .o(n_13754) );
na02f02 g54458_u0 ( .a(n_16299), .b(n_12956), .o(g54458_p) );
in01f04 g54458_u1 ( .a(g54458_p), .o(n_13486) );
no02f02 g54459_u0 ( .a(n_13304), .b(pci_target_unit_del_sync_be_out_reg_0__Q), .o(n_13306) );
na02f02 g54460_u0 ( .a(n_14967), .b(n_13122), .o(n_14895) );
no02f02 g54461_u0 ( .a(n_13304), .b(pci_target_unit_del_sync_be_out_reg_1__Q), .o(n_13305) );
no02f02 g54462_u0 ( .a(n_13304), .b(pci_target_unit_del_sync_be_out_reg_2__Q), .o(n_13303) );
no02f02 g54463_u0 ( .a(n_13304), .b(pci_target_unit_del_sync_be_out_reg_3__Q), .o(n_13302) );
no02f01 g54464_u0 ( .a(FE_OFN969_n_13784), .b(n_12595), .o(TIMEBOOST_net_13971) );
na02f02 g54465_u0 ( .a(n_12776), .b(n_12595), .o(g54465_p) );
in01f04 g54465_u1 ( .a(g54465_p), .o(n_13341) );
no02f02 g54466_u0 ( .a(FE_OFN2165_n_16301), .b(n_8757), .o(n_13481) );
na03f02 TIMEBOOST_cell_73565 ( .a(TIMEBOOST_net_20580), .b(FE_OFN1232_n_6391), .c(g62697_sb), .o(n_6160) );
in01s01 g54468_u0 ( .a(n_12855), .o(n_12954) );
no02s01 g54470_u0 ( .a(n_13721), .b(n_14905), .o(n_12855) );
in01f02 g54471_u0 ( .a(n_13617), .o(g54471_sb) );
na04f04 TIMEBOOST_cell_24607 ( .a(n_9002), .b(g57547_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q), .d(FE_OFN2167_n_8567), .o(n_10306) );
na03f02 TIMEBOOST_cell_72530 ( .a(TIMEBOOST_net_21380), .b(g64177_sb), .c(FE_OFN877_g64577_p), .o(TIMEBOOST_net_22639) );
na04f06 TIMEBOOST_cell_73207 ( .a(TIMEBOOST_net_14856), .b(FE_OFN1149_n_13249), .c(n_1782), .d(g54141_sb), .o(n_13666) );
in01f02 g54472_u0 ( .a(n_13617), .o(g54472_sb) );
na04f04 TIMEBOOST_cell_24591 ( .a(n_9491), .b(g57461_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q), .d(FE_OFN2187_n_8567), .o(n_11273) );
na03m02 TIMEBOOST_cell_65656 ( .a(TIMEBOOST_net_12714), .b(TIMEBOOST_net_9860), .c(n_6), .o(TIMEBOOST_net_20966) );
in01f02 g54474_u0 ( .a(n_16967), .o(n_13479) );
in01f02 g54480_u0 ( .a(n_16205), .o(n_13475) );
in01f02 g54484_u0 ( .a(n_13617), .o(g54484_sb) );
na04f04 TIMEBOOST_cell_24593 ( .a(n_9025), .b(g57449_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q), .d(FE_OFN2168_n_8567), .o(n_10348) );
in01f02 g54485_u0 ( .a(n_13617), .o(g54485_sb) );
na04f04 TIMEBOOST_cell_24595 ( .a(n_8563), .b(g58587_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q), .d(FE_OFN2185_n_8567), .o(n_8916) );
na03f01 TIMEBOOST_cell_67157 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q), .b(n_3755), .c(FE_OFN682_n_4460), .o(TIMEBOOST_net_10520) );
na03m06 TIMEBOOST_cell_68822 ( .a(g64816_db), .b(g64816_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_21619) );
in01f02 g54486_u0 ( .a(n_13617), .o(g54486_sb) );
na04f04 TIMEBOOST_cell_24597 ( .a(n_9411), .b(g57588_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q), .d(FE_OFN2184_n_8567), .o(n_11164) );
na04f04 TIMEBOOST_cell_24565 ( .a(n_9226), .b(g57130_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q), .d(FE_OFN1417_n_8567), .o(n_10839) );
na03f02 TIMEBOOST_cell_73118 ( .a(g64232_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q), .c(TIMEBOOST_net_23308), .o(TIMEBOOST_net_9983) );
in01f02 g54487_u0 ( .a(n_13617), .o(g54487_sb) );
na04f04 TIMEBOOST_cell_24605 ( .a(n_9202), .b(g57559_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q), .d(FE_OFN2175_n_8567), .o(n_10802) );
na02s01 TIMEBOOST_cell_45675 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q), .o(TIMEBOOST_net_13732) );
na02f02 TIMEBOOST_cell_70569 ( .a(TIMEBOOST_net_22492), .b(g63120_sb), .o(n_5016) );
in01f02 g54488_u0 ( .a(n_13617), .o(g54488_sb) );
na04f04 TIMEBOOST_cell_24599 ( .a(n_9414), .b(g57581_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q), .d(FE_OFN2177_n_8567), .o(n_11169) );
na02s02 TIMEBOOST_cell_49416 ( .a(TIMEBOOST_net_14925), .b(FE_OFN569_n_9528), .o(TIMEBOOST_net_12975) );
na03s02 TIMEBOOST_cell_73353 ( .a(TIMEBOOST_net_12431), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q), .c(FE_OFN587_n_9692), .o(TIMEBOOST_net_15217) );
in01f02 g54489_u0 ( .a(n_13617), .o(g54489_sb) );
na02m10 TIMEBOOST_cell_45711 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q), .o(TIMEBOOST_net_13750) );
na02f01 TIMEBOOST_cell_26618 ( .a(TIMEBOOST_net_7413), .b(g62720_sb), .o(n_5543) );
in01f02 g54490_u0 ( .a(n_13617), .o(g54490_sb) );
na04f04 TIMEBOOST_cell_24601 ( .a(n_8997), .b(g57566_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q), .d(FE_OFN2168_n_8567), .o(n_10296) );
in01s01 TIMEBOOST_cell_45992 ( .a(TIMEBOOST_net_13952), .o(TIMEBOOST_net_13953) );
in01f02 g54491_u0 ( .a(n_13617), .o(g54491_sb) );
na04f04 TIMEBOOST_cell_24603 ( .a(n_9427), .b(g57562_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q), .d(FE_OFN2180_n_8567), .o(n_11190) );
no04f08 TIMEBOOST_cell_72461 ( .a(TIMEBOOST_net_21290), .b(n_300), .c(FE_RN_638_0), .d(FE_RN_636_0), .o(FE_RN_641_0) );
na02s01 TIMEBOOST_cell_42891 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q), .o(TIMEBOOST_net_12340) );
in01f02 g54492_u0 ( .a(n_13617), .o(g54492_sb) );
na04f04 TIMEBOOST_cell_24623 ( .a(n_9814), .b(g57111_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q), .d(FE_OFN2182_n_8567), .o(n_11635) );
na02s01 TIMEBOOST_cell_48491 ( .a(FE_OFN1648_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q), .o(TIMEBOOST_net_14463) );
na02s01 TIMEBOOST_cell_37042 ( .a(pci_ad_i_24_), .b(parchk_pci_ad_reg_in_1228), .o(TIMEBOOST_net_10133) );
in01f02 g54493_u0 ( .a(n_13617), .o(g54493_sb) );
na04f04 TIMEBOOST_cell_24625 ( .a(n_9231), .b(g57094_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q), .d(FE_OFN2184_n_8567), .o(n_10845) );
na03f02 TIMEBOOST_cell_24957 ( .a(FE_RN_146_0), .b(n_10912), .c(n_12571), .o(n_12833) );
na02f02 TIMEBOOST_cell_27243 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_7726) );
in01f02 g54494_u0 ( .a(n_13617), .o(g54494_sb) );
na04f04 TIMEBOOST_cell_24571 ( .a(n_9020), .b(g57475_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q), .d(FE_OFN2167_n_8567), .o(n_10338) );
na02s01 TIMEBOOST_cell_37044 ( .a(pci_ad_i_26_), .b(parchk_pci_ad_reg_in_1230), .o(TIMEBOOST_net_10134) );
in01f02 g54495_u0 ( .a(n_13617), .o(g54495_sb) );
na03f02 TIMEBOOST_cell_66314 ( .a(TIMEBOOST_net_13364), .b(n_6232), .c(g62491_sb), .o(n_6603) );
oa12f01 g54496_u0 ( .a(n_13474), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .c(n_13617), .o(n_13682) );
in01f20 g54504_u0 ( .a(n_13784), .o(TIMEBOOST_net_5253) );
in01f10 g54510_u0 ( .a(n_12776), .o(n_13763) );
in01f08 g54511_u0 ( .a(n_12776), .o(n_13781) );
in01f20 g54512_u0 ( .a(FE_OFN969_n_13784), .o(n_12776) );
in01s01 g54519_u0 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_766), .o(n_12952) );
na02f02 g54549_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .b(n_13617), .o(n_13474) );
no02f02 g54567_u0 ( .a(n_12764), .b(n_12819), .o(n_12964) );
na02f02 g54568_u0 ( .a(n_12946), .b(n_12756), .o(g54568_p) );
in01f02 g54568_u1 ( .a(g54568_p), .o(n_13068) );
na02f02 g54569_u0 ( .a(n_12943), .b(n_12528), .o(g54569_p) );
in01f02 g54569_u1 ( .a(g54569_p), .o(n_13067) );
no02f02 g54570_u0 ( .a(n_12818), .b(n_12806), .o(n_12963) );
no02f02 g54571_u0 ( .a(n_12817), .b(n_12741), .o(n_12962) );
na02f02 g54572_u0 ( .a(n_12936), .b(n_12736), .o(g54572_p) );
in01f02 g54572_u1 ( .a(g54572_p), .o(n_13063) );
na02f02 g54573_u0 ( .a(n_12731), .b(n_12933), .o(g54573_p) );
in01f02 g54573_u1 ( .a(g54573_p), .o(n_13066) );
na02f02 g54574_u0 ( .a(n_12930), .b(n_12725), .o(g54574_p) );
in01f02 g54574_u1 ( .a(g54574_p), .o(n_13065) );
in01f02 g54575_u0 ( .a(n_13064), .o(n_13120) );
na02f02 g54576_u0 ( .a(n_12519), .b(n_12927), .o(n_13064) );
na02f02 g54579_u0 ( .a(n_12921), .b(n_12709), .o(g54579_p) );
in01f02 g54579_u1 ( .a(g54579_p), .o(n_13059) );
na02f02 g54580_u0 ( .a(n_12705), .b(n_12919), .o(g54580_p) );
in01f02 g54580_u1 ( .a(g54580_p), .o(n_13061) );
na02f02 g54581_u0 ( .a(n_12916), .b(n_12699), .o(g54581_p) );
in01f02 g54581_u1 ( .a(g54581_p), .o(n_13060) );
in01f02 g54582_u0 ( .a(n_12961), .o(n_13058) );
na02f02 g54583_u0 ( .a(n_12693), .b(n_12815), .o(n_12961) );
in01f02 g54584_u0 ( .a(n_13057), .o(n_13118) );
na02f02 g54585_u0 ( .a(n_12688), .b(n_12911), .o(n_13057) );
na02f02 g54586_u0 ( .a(n_12682), .b(n_12908), .o(g54586_p) );
in01f02 g54586_u1 ( .a(g54586_p), .o(n_13056) );
na02f02 g54587_u0 ( .a(n_12905), .b(n_12503), .o(g54587_p) );
in01f02 g54587_u1 ( .a(g54587_p), .o(n_13055) );
no02f02 g54588_u0 ( .a(n_12813), .b(n_12676), .o(n_12960) );
no02f02 g54589_u0 ( .a(n_12672), .b(n_12901), .o(n_13054) );
no02f02 g54590_u0 ( .a(n_12898), .b(n_12667), .o(n_13053) );
na02f02 g54591_u0 ( .a(n_12812), .b(n_12662), .o(g54591_p) );
in01f02 g54591_u1 ( .a(g54591_p), .o(n_12959) );
no02f02 g54592_u0 ( .a(n_12811), .b(n_12788), .o(n_12958) );
na02f02 g54593_u0 ( .a(n_12891), .b(n_12495), .o(g54593_p) );
in01f02 g54593_u1 ( .a(g54593_p), .o(n_13052) );
na02f02 g54594_u0 ( .a(n_12888), .b(n_12647), .o(g54594_p) );
in01f02 g54594_u1 ( .a(g54594_p), .o(n_13051) );
na02f02 g54595_u0 ( .a(n_12885), .b(n_12642), .o(g54595_p) );
in01f02 g54595_u1 ( .a(g54595_p), .o(n_13050) );
na02f02 g54596_u0 ( .a(n_12882), .b(n_12636), .o(g54596_p) );
in01f02 g54596_u1 ( .a(g54596_p), .o(n_13049) );
na02f06 g54597_u0 ( .a(n_13116), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in), .o(g54597_p) );
in01f06 g54597_u1 ( .a(g54597_p), .o(n_13621) );
no02f02 g54598_u0 ( .a(n_12810), .b(n_12784), .o(n_12957) );
no02f02 g54599_u0 ( .a(n_12877), .b(n_12783), .o(n_13048) );
no02f02 g54600_u0 ( .a(n_12623), .b(n_12874), .o(n_13047) );
na02f02 g54601_u0 ( .a(n_12871), .b(n_12619), .o(g54601_p) );
in01f02 g54601_u1 ( .a(g54601_p), .o(n_13046) );
no02f02 g54602_u0 ( .a(n_12868), .b(n_12614), .o(n_13045) );
na02f02 g54603_u0 ( .a(n_12865), .b(n_12484), .o(g54603_p) );
in01f02 g54603_u1 ( .a(g54603_p), .o(n_13044) );
in01f02 g54604_u0 ( .a(n_13043), .o(n_13117) );
na02f02 g54605_u0 ( .a(n_12602), .b(n_12862), .o(n_13043) );
na02f02 g54606_u0 ( .a(n_12859), .b(n_12480), .o(g54606_p) );
in01f02 g54606_u1 ( .a(g54606_p), .o(n_13042) );
in01f20 g54610_u0 ( .a(n_13363), .o(n_14725) );
in01f06 g54616_u0 ( .a(n_13363), .o(n_14800) );
na03m02 TIMEBOOST_cell_70072 ( .a(n_2207), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q), .c(FE_OFN2257_n_8060), .o(TIMEBOOST_net_22244) );
na02s01 TIMEBOOST_cell_52627 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_16531) );
in01f04 g54665_u0 ( .a(n_13122), .o(n_13304) );
in01f06 g54666_u0 ( .a(n_12956), .o(n_13122) );
oa12f02 g54669_u0 ( .a(n_8727), .b(n_8730), .c(n_10825), .o(n_12170) );
na02f02 g54670_u0 ( .a(n_12947), .b(n_12948), .o(n_13041) );
na02f02 g54672_u0 ( .a(n_12942), .b(n_12941), .o(n_17028) );
na02f02 g54673_u0 ( .a(n_12937), .b(n_12938), .o(n_16600) );
na02f02 g54674_u0 ( .a(n_12935), .b(n_12934), .o(n_16602) );
no02f02 g54677_u0 ( .a(n_12814), .b(n_12904), .o(n_13034) );
na02f02 g54678_u0 ( .a(n_12894), .b(n_12895), .o(n_15440) );
na02f02 g54679_u0 ( .a(n_12893), .b(n_12892), .o(n_16588) );
na02f02 g54680_u0 ( .a(n_12878), .b(n_12879), .o(n_15438) );
na02f02 g54681_u0 ( .a(n_12876), .b(n_12875), .o(n_16591) );
no02f02 g54716_u0 ( .a(n_12166), .b(n_11014), .o(n_12591) );
no02f02 g54717_u0 ( .a(n_12165), .b(n_11741), .o(n_12590) );
no02f02 g54718_u0 ( .a(n_12164), .b(n_11740), .o(n_12589) );
no02f02 g54719_u0 ( .a(n_12163), .b(n_10987), .o(n_12588) );
no02f02 g54720_u0 ( .a(n_12162), .b(n_10764), .o(n_12587) );
no02f02 g54721_u0 ( .a(n_12161), .b(n_10978), .o(n_12586) );
no02f02 g54722_u0 ( .a(n_12160), .b(n_10976), .o(n_12585) );
no02f02 g54723_u0 ( .a(n_12159), .b(n_10975), .o(n_12584) );
no02f02 g54724_u0 ( .a(n_12158), .b(n_10971), .o(n_12583) );
no02f02 g54726_u0 ( .a(n_12156), .b(n_10963), .o(n_12581) );
no02f02 g54727_u0 ( .a(n_12155), .b(n_10962), .o(n_12580) );
no02f02 g54728_u0 ( .a(n_12154), .b(n_10952), .o(n_12579) );
no02f02 g54729_u0 ( .a(n_11847), .b(n_11738), .o(n_12442) );
no02f02 g54730_u0 ( .a(n_12153), .b(n_10943), .o(n_12578) );
no02f02 g54731_u0 ( .a(n_17041), .b(n_17042), .o(n_12577) );
no02f02 g54733_u0 ( .a(n_11846), .b(n_10932), .o(n_12441) );
no02f02 g54734_u0 ( .a(n_11736), .b(n_12439), .o(n_12772) );
no02f02 g54735_u0 ( .a(n_12148), .b(n_10923), .o(n_12575) );
no02f02 g54736_u0 ( .a(n_12147), .b(n_10638), .o(n_12574) );
no02f02 g54737_u0 ( .a(n_10631), .b(n_12146), .o(n_12573) );
no02f02 g54738_u0 ( .a(n_12145), .b(n_10919), .o(n_12572) );
no02f02 g54739_u0 ( .a(n_11845), .b(n_10917), .o(n_12440) );
no02f02 g54740_u0 ( .a(n_12144), .b(n_10913), .o(n_12571) );
no02f02 g54741_u0 ( .a(n_12143), .b(n_11734), .o(n_12570) );
no02f02 g54742_u0 ( .a(n_12141), .b(n_10906), .o(n_12569) );
no02f02 g54743_u0 ( .a(n_12140), .b(n_11731), .o(n_12568) );
no02f02 g54744_u0 ( .a(n_12139), .b(n_11727), .o(n_12567) );
no02f02 g54745_u0 ( .a(n_12137), .b(n_11880), .o(n_12566) );
no02f02 g54746_u0 ( .a(n_12135), .b(n_11724), .o(n_12565) );
no02f02 g54747_u0 ( .a(n_12134), .b(n_10882), .o(n_12564) );
no02f02 g54748_u0 ( .a(n_12133), .b(n_10876), .o(n_12563) );
no02f02 g54749_u0 ( .a(n_12132), .b(n_10867), .o(n_12562) );
no02f02 g54750_u0 ( .a(n_12130), .b(n_11718), .o(n_12561) );
no02f02 g54751_u0 ( .a(n_12129), .b(n_10860), .o(n_12560) );
no02f02 g54752_u0 ( .a(n_12128), .b(n_10856), .o(n_12559) );
no02f02 g54754_u0 ( .a(n_12768), .b(n_12767), .o(n_12950) );
no02f02 g54755_u0 ( .a(n_12765), .b(n_12766), .o(n_12949) );
no02f02 g54757_u0 ( .a(n_12763), .b(n_12762), .o(n_12948) );
no02f02 g54758_u0 ( .a(n_12761), .b(n_12760), .o(n_12947) );
no02f02 g54759_u0 ( .a(n_12757), .b(n_12758), .o(n_12946) );
no02f02 g54762_u0 ( .a(n_12750), .b(n_12751), .o(n_12943) );
no02f02 g54763_u0 ( .a(n_12749), .b(n_12748), .o(n_12942) );
no02f02 g54764_u0 ( .a(n_12746), .b(n_12747), .o(n_12941) );
no02f02 g54766_u0 ( .a(n_12744), .b(n_12745), .o(n_12940) );
no02f02 g54767_u0 ( .a(n_12743), .b(n_12742), .o(n_12939) );
no02f02 g54769_u0 ( .a(n_17036), .b(n_17035), .o(n_12938) );
no02f02 g54770_u0 ( .a(n_12738), .b(n_12527), .o(n_12937) );
no02f02 g54771_u0 ( .a(n_12526), .b(n_12737), .o(n_12936) );
no02f02 g54772_u0 ( .a(n_12734), .b(n_12735), .o(n_12935) );
no02f02 g54773_u0 ( .a(n_12733), .b(n_12525), .o(n_12934) );
no02f02 g54774_u0 ( .a(n_12732), .b(n_12524), .o(n_12933) );
no02f02 g54775_u0 ( .a(n_12523), .b(n_12729), .o(n_12932) );
no02f02 g54776_u0 ( .a(n_12728), .b(n_12727), .o(n_12931) );
no02f02 g54777_u0 ( .a(n_12726), .b(n_12522), .o(n_12930) );
no02f02 g54778_u0 ( .a(n_12723), .b(n_12724), .o(n_12929) );
no02f02 g54779_u0 ( .a(n_12521), .b(n_12722), .o(n_12928) );
no02f02 g54780_u0 ( .a(n_12520), .b(n_12720), .o(n_12927) );
no02f02 g54783_u0 ( .a(n_12518), .b(n_12715), .o(n_12924) );
no02f02 g54784_u0 ( .a(n_12517), .b(n_12713), .o(n_12923) );
no02f02 g54785_u0 ( .a(n_12712), .b(n_12711), .o(n_12922) );
no02f02 g54786_u0 ( .a(n_12710), .b(n_12516), .o(n_12921) );
no02f02 g54789_u0 ( .a(n_12515), .b(n_12706), .o(n_12919) );
no02f04 g54790_u0 ( .a(n_12703), .b(n_12704), .o(n_12918) );
no02f02 g54791_u0 ( .a(n_12701), .b(n_12702), .o(n_12917) );
no02f02 g54792_u0 ( .a(n_12700), .b(n_12514), .o(n_12916) );
no02f02 g54793_u0 ( .a(n_12513), .b(n_12697), .o(n_12915) );
no02f02 g54794_u0 ( .a(n_12512), .b(n_12696), .o(n_12914) );
no02f02 g54795_u0 ( .a(n_12510), .b(n_12511), .o(n_12815) );
no02f02 g54796_u0 ( .a(n_12509), .b(n_12692), .o(n_12913) );
no02f02 g54798_u0 ( .a(n_12689), .b(n_12508), .o(n_12911) );
no02f02 g54801_u0 ( .a(n_12683), .b(n_12684), .o(n_12908) );
no02f02 g54802_u0 ( .a(n_12506), .b(n_12680), .o(n_12907) );
no02f02 g54803_u0 ( .a(n_12679), .b(n_12505), .o(n_12906) );
no02f02 g54804_u0 ( .a(n_12504), .b(n_12678), .o(n_12905) );
na04f04 g54807_u0 ( .a(n_11957), .b(n_12378), .c(n_11956), .d(n_11818), .o(n_12813) );
no02f02 g54808_u0 ( .a(n_12500), .b(n_12675), .o(n_12903) );
no02f02 g54809_u0 ( .a(n_12674), .b(n_12673), .o(n_12902) );
na02f02 TIMEBOOST_cell_63912 ( .a(n_2693), .b(FE_OFN1700_n_5751), .o(TIMEBOOST_net_20942) );
no02f02 g54811_u0 ( .a(n_12670), .b(n_12671), .o(n_12900) );
no02f02 g54812_u0 ( .a(n_12668), .b(n_12669), .o(n_12899) );
no02f02 g54814_u0 ( .a(n_12665), .b(n_12666), .o(n_12897) );
no02f02 g54815_u0 ( .a(n_12664), .b(n_12663), .o(n_12896) );
no02f02 g54816_u0 ( .a(n_12498), .b(n_12499), .o(n_12812) );
no02f02 g54817_u0 ( .a(n_12661), .b(n_12660), .o(n_12895) );
no02f02 g54818_u0 ( .a(n_12658), .b(n_12659), .o(n_12894) );
na04f04 g54819_u0 ( .a(n_11938), .b(n_11814), .c(n_11937), .d(n_12075), .o(n_12811) );
no02f02 g54820_u0 ( .a(n_12655), .b(n_12656), .o(n_12893) );
no02f02 g54821_u0 ( .a(n_12654), .b(n_12653), .o(n_12892) );
no02f02 g54822_u0 ( .a(n_12496), .b(n_12652), .o(n_12891) );
no02f02 g54823_u0 ( .a(n_12494), .b(n_12651), .o(n_12890) );
no02f02 g54824_u0 ( .a(n_12649), .b(n_12650), .o(n_12889) );
no02f02 g54825_u0 ( .a(n_12648), .b(n_12493), .o(n_12888) );
no02f02 g54826_u0 ( .a(n_12492), .b(n_12646), .o(n_12887) );
no02f02 g54827_u0 ( .a(n_12645), .b(n_12644), .o(n_12886) );
no02f02 g54828_u0 ( .a(n_12643), .b(n_12491), .o(n_12885) );
no02f02 g54829_u0 ( .a(n_12641), .b(n_12640), .o(n_12884) );
no02f02 g54830_u0 ( .a(n_12639), .b(n_12638), .o(n_12883) );
no02f02 g54831_u0 ( .a(n_12637), .b(n_12490), .o(n_12882) );
no02f02 g54832_u0 ( .a(FE_OFN186_n_15768), .b(n_15759), .o(n_11450) );
na04f04 TIMEBOOST_cell_24654 ( .a(n_9712), .b(g57224_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q), .d(FE_OFN2188_n_8567), .o(n_11532) );
in01f10 g54834_u0 ( .a(n_13116), .o(n_13617) );
in01f08 g54838_u0 ( .a(n_16981), .o(n_13116) );
no02f02 g54840_u0 ( .a(n_12635), .b(n_12489), .o(n_12881) );
no02f02 g54841_u0 ( .a(n_12633), .b(n_12634), .o(n_12880) );
no02f02 g54843_u0 ( .a(n_12630), .b(n_12631), .o(n_12879) );
no02f02 g54844_u0 ( .a(n_12628), .b(n_12629), .o(n_12878) );
no02f02 g54846_u0 ( .a(n_12625), .b(n_12626), .o(n_12876) );
no02f02 g54847_u0 ( .a(n_12624), .b(n_12488), .o(n_12875) );
no02f02 g54849_u0 ( .a(n_12487), .b(n_12622), .o(n_12873) );
no02f02 g54850_u0 ( .a(n_12621), .b(n_12486), .o(n_12872) );
no02f02 g54851_u0 ( .a(n_12620), .b(n_12485), .o(n_12871) );
no02f02 g54852_u0 ( .a(n_12617), .b(n_12618), .o(n_12870) );
no02f02 g54853_u0 ( .a(n_12616), .b(n_12615), .o(n_12869) );
no02f02 g54855_u0 ( .a(n_12613), .b(n_12612), .o(n_12867) );
no02f02 g54856_u0 ( .a(n_12611), .b(n_12610), .o(n_12866) );
no02f02 g54857_u0 ( .a(n_16597), .b(n_16596), .o(n_12865) );
no02f02 g54858_u0 ( .a(n_12606), .b(n_12607), .o(n_12864) );
no02f02 g54859_u0 ( .a(n_12604), .b(n_12605), .o(n_12863) );
no02f02 g54860_u0 ( .a(n_12603), .b(n_12483), .o(n_12862) );
no02f02 g54863_u0 ( .a(n_12481), .b(n_12596), .o(n_12859) );
in01f01 g54864_u0 ( .a(n_12167), .o(n_12168) );
in01f02 g54865_u0 ( .a(n_15611), .o(n_12167) );
na04f02 g54867_u0 ( .a(n_17016), .b(n_11157), .c(n_11144), .d(n_17017), .o(n_12558) );
na04f02 g54868_u0 ( .a(n_11796), .b(n_11153), .c(n_11147), .d(n_11155), .o(n_12557) );
na04f02 g54869_u0 ( .a(n_11793), .b(n_11152), .c(n_11149), .d(n_11148), .o(n_12556) );
na04f02 g54870_u0 ( .a(n_11142), .b(n_11143), .c(n_11146), .d(n_11145), .o(n_12555) );
na04f02 g54872_u0 ( .a(n_11135), .b(n_11134), .c(n_11131), .d(n_11132), .o(n_12553) );
na04f02 g54874_u0 ( .a(n_11129), .b(n_11126), .c(n_16581), .d(n_16582), .o(n_12552) );
na04f02 g54875_u0 ( .a(n_10788), .b(n_11124), .c(n_11122), .d(n_11123), .o(n_12551) );
na04f02 g54876_u0 ( .a(n_11121), .b(n_11120), .c(n_11118), .d(n_11119), .o(n_12550) );
na04f02 g54877_u0 ( .a(n_16583), .b(n_11115), .c(n_11113), .d(n_16584), .o(n_12549) );
na04f02 g54878_u0 ( .a(n_11111), .b(n_11110), .c(n_11108), .d(n_11109), .o(n_12548) );
na04f02 g54879_u0 ( .a(n_11790), .b(n_11107), .c(n_11104), .d(n_11106), .o(n_12547) );
na04f02 g54883_u0 ( .a(n_11086), .b(n_11786), .c(n_11087), .d(n_10784), .o(n_12770) );
na04f02 g54884_u0 ( .a(n_11090), .b(n_11088), .c(n_11089), .d(n_10785), .o(n_12543) );
na04f02 g54885_u0 ( .a(n_11085), .b(n_11784), .c(n_11084), .d(n_11083), .o(n_12542) );
na04f02 g54886_u0 ( .a(n_16586), .b(n_16585), .c(n_11079), .d(n_11081), .o(n_12541) );
na04f02 g54887_u0 ( .a(n_11078), .b(n_11077), .c(n_11075), .d(n_11076), .o(n_12540) );
na04f02 g54888_u0 ( .a(n_11782), .b(n_11783), .c(n_11072), .d(n_11073), .o(n_12539) );
na04f02 g54890_u0 ( .a(n_11065), .b(n_10782), .c(n_11066), .d(n_11067), .o(n_12537) );
na04f02 g54891_u0 ( .a(n_11063), .b(n_11780), .c(n_11064), .d(n_11778), .o(n_12536) );
na04f02 g54893_u0 ( .a(n_11776), .b(n_11059), .c(n_11057), .d(n_11058), .o(n_12534) );
na04f02 g54895_u0 ( .a(n_11050), .b(n_11049), .c(n_11051), .d(n_11048), .o(n_12532) );
na04f02 g54896_u0 ( .a(n_11775), .b(n_11044), .c(n_11047), .d(n_11046), .o(n_12531) );
na04f02 g54897_u0 ( .a(n_10781), .b(n_11043), .c(n_11774), .d(n_11042), .o(n_12769) );
na04f02 g54899_u0 ( .a(n_11038), .b(n_11034), .c(n_11037), .d(n_11036), .o(n_12529) );
in01f03 g54903_u0 ( .a(n_16131), .o(n_12858) );
in01f02 g54907_u0 ( .a(n_15301), .o(n_10825) );
na02m02 TIMEBOOST_cell_69310 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q), .b(n_4447), .o(TIMEBOOST_net_21863) );
na02m02 TIMEBOOST_cell_68630 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q), .o(TIMEBOOST_net_21523) );
na04f04 TIMEBOOST_cell_24376 ( .a(n_9432), .b(g57551_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q), .d(FE_OFN1408_n_8567), .o(n_11193) );
ao12f02 g54936_u0 ( .a(n_12479), .b(FE_OFN1553_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q), .o(n_12809) );
na02s01 TIMEBOOST_cell_48902 ( .a(TIMEBOOST_net_14668), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_12788) );
na02m02 TIMEBOOST_cell_53817 ( .a(n_4519), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q), .o(TIMEBOOST_net_17126) );
no02f10 TIMEBOOST_cell_53982 ( .a(TIMEBOOST_net_17208), .b(FE_RN_503_0), .o(n_2253) );
na03f02 TIMEBOOST_cell_65926 ( .a(TIMEBOOST_net_20431), .b(FE_OFN1170_n_5592), .c(g62138_sb), .o(n_5555) );
na04f04 TIMEBOOST_cell_24382 ( .a(n_9802), .b(g57120_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q), .d(FE_OFN1424_n_8567), .o(n_11625) );
na02f02 TIMEBOOST_cell_70339 ( .a(TIMEBOOST_net_22377), .b(g63592_sb), .o(n_7203) );
ao12f02 g54945_u0 ( .a(n_12417), .b(FE_OFN1757_n_12681), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q), .o(n_12756) );
na03m02 TIMEBOOST_cell_73016 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .c(pci_target_unit_pcit_if_strd_addr_in_712), .o(TIMEBOOST_net_22181) );
na03m02 TIMEBOOST_cell_72635 ( .a(g65056_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q), .c(TIMEBOOST_net_10572), .o(TIMEBOOST_net_20545) );
na02s01 g58419_u2 ( .a(FE_OFN207_n_9865), .b(FE_OFN1651_n_9428), .o(g58419_db) );
na02m02 TIMEBOOST_cell_53653 ( .a(TIMEBOOST_net_13230), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_17044) );
ao12f02 g54953_u0 ( .a(n_12044), .b(FE_OFN1749_n_12004), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q), .o(n_12528) );
na02s02 g58409_u2 ( .a(FE_OFN1656_n_9502), .b(FE_OFN215_n_9856), .o(g58409_db) );
na02s02 g58408_u2 ( .a(FE_OFN254_n_9825), .b(FE_OFN579_n_9531), .o(g58408_db) );
na03s02 TIMEBOOST_cell_41714 ( .a(g58423_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q), .c(g58423_db), .o(n_8997) );
na02s01 TIMEBOOST_cell_43125 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q), .o(TIMEBOOST_net_12457) );
no02f10 TIMEBOOST_cell_62401 ( .a(TIMEBOOST_net_20147), .b(FE_RN_709_0), .o(n_15755) );
na02s01 TIMEBOOST_cell_49531 ( .a(FE_OFN1666_n_9477), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q), .o(TIMEBOOST_net_14983) );
na02s01 TIMEBOOST_cell_44113 ( .a(FE_OFN262_n_9851), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q), .o(TIMEBOOST_net_12951) );
na04f04 TIMEBOOST_cell_24392 ( .a(n_9007), .b(g57530_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q), .d(FE_OFN1385_n_8567), .o(n_10314) );
na04m02 TIMEBOOST_cell_67302 ( .a(n_4488), .b(g65088_sb), .c(FE_OFN659_n_4392), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q), .o(n_4302) );
ao12f02 g54964_u0 ( .a(n_12478), .b(FE_OFN1553_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q), .o(n_12805) );
na02m02 TIMEBOOST_cell_53030 ( .a(TIMEBOOST_net_16732), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_15314) );
na02s01 g58364_u2 ( .a(FE_OFN241_n_9830), .b(FE_OFN548_n_9477), .o(g58364_db) );
na02s02 TIMEBOOST_cell_48946 ( .a(TIMEBOOST_net_14690), .b(g63618_db), .o(TIMEBOOST_net_13017) );
na02s01 TIMEBOOST_cell_52629 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_16532) );
na03f02 TIMEBOOST_cell_68030 ( .a(TIMEBOOST_net_17449), .b(FE_OFN1268_n_4095), .c(g62554_sb), .o(n_6456) );
ao12f02 g54973_u0 ( .a(n_12300), .b(FE_OFN1734_n_16317), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q), .o(n_12736) );
na02m01 g58363_u2 ( .a(FE_OFN239_n_9832), .b(FE_OFN1668_n_9477), .o(g58363_db) );
na04f04 TIMEBOOST_cell_24400 ( .a(n_9761), .b(g57159_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q), .d(FE_OFN1384_n_8567), .o(n_11590) );
na02s01 g58361_u2 ( .a(FE_OFN1666_n_9477), .b(FE_OFN235_n_9834), .o(g58361_db) );
in01s01 TIMEBOOST_cell_45946 ( .a(TIMEBOOST_net_13906), .o(TIMEBOOST_net_13907) );
na04f04 TIMEBOOST_cell_24402 ( .a(n_9767), .b(g57155_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q), .d(FE_OFN1424_n_8567), .o(n_11595) );
na02f02 TIMEBOOST_cell_70056 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q), .b(FE_OFN704_n_8069), .o(TIMEBOOST_net_22236) );
ao12f02 g54981_u0 ( .a(n_12294), .b(FE_OFN1734_n_16317), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q), .o(n_12731) );
na04f04 TIMEBOOST_cell_24404 ( .a(n_9770), .b(g57151_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q), .d(FE_OFN1406_n_8567), .o(n_11599) );
na03f02 TIMEBOOST_cell_66953 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_16502), .c(FE_OFN2210_n_11027), .o(n_12702) );
ao12f02 g54986_u0 ( .a(n_12476), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q), .o(n_12801) );
na02f02 TIMEBOOST_cell_69173 ( .a(TIMEBOOST_net_21794), .b(TIMEBOOST_net_12634), .o(TIMEBOOST_net_17333) );
na04f04 TIMEBOOST_cell_24408 ( .a(n_9779), .b(g57145_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q), .d(FE_OFN1405_n_8567), .o(n_11605) );
na03f10 TIMEBOOST_cell_72383 ( .a(n_1442), .b(n_2914), .c(n_2397), .o(TIMEBOOST_net_12739) );
na02m04 TIMEBOOST_cell_69430 ( .a(g64796_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q), .o(TIMEBOOST_net_21923) );
na04f04 TIMEBOOST_cell_24412 ( .a(n_9897), .b(g57193_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q), .d(FE_OFN1385_n_8567), .o(n_11560) );
ao12f01 g54996_u0 ( .a(n_12003), .b(FE_OFN1562_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q), .o(n_12519) );
na03f02 TIMEBOOST_cell_66801 ( .a(n_7226), .b(g59370_sb), .c(TIMEBOOST_net_7726), .o(n_7694) );
na03f02 TIMEBOOST_cell_66323 ( .a(TIMEBOOST_net_13371), .b(n_6232), .c(g62655_sb), .o(n_6234) );
na02m01 TIMEBOOST_cell_69294 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q), .o(TIMEBOOST_net_21855) );
na03f02 TIMEBOOST_cell_73354 ( .a(n_2224), .b(FE_OFN1699_n_5751), .c(TIMEBOOST_net_9627), .o(TIMEBOOST_net_22957) );
ao12f02 g55005_u0 ( .a(n_12280), .b(FE_OFN1759_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q), .o(n_12714) );
na03m06 TIMEBOOST_cell_64801 ( .a(n_3761), .b(FE_OFN1663_n_4490), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q), .o(TIMEBOOST_net_16270) );
na02s04 TIMEBOOST_cell_68130 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_95), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_21273) );
na03m06 TIMEBOOST_cell_68406 ( .a(g64095_sb), .b(pci_target_unit_fifos_pciw_addr_data_in_140), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q), .o(TIMEBOOST_net_21411) );
na04f04 TIMEBOOST_cell_24420 ( .a(n_9494), .b(g57456_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q), .d(FE_OFN1376_n_8567), .o(n_11277) );
na02m04 TIMEBOOST_cell_25488 ( .a(TIMEBOOST_net_6848), .b(n_7835), .o(TIMEBOOST_net_686) );
ao12f02 g55018_u0 ( .a(n_12271), .b(FE_OFN1735_n_16317), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q), .o(n_12705) );
na02m01 g63616_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q), .b(FE_OFN1079_n_4778), .o(g63616_db) );
na04f04 TIMEBOOST_cell_24426 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .b(g58621_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .d(FE_OFN1369_n_8567), .o(n_9181) );
na02s01 g65858_u2 ( .a(pci_target_unit_del_sync_addr_in_221), .b(FE_OFN776_n_15366), .o(g65858_db) );
ao12f04 g55023_u0 ( .a(n_12459), .b(FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q), .o(n_12797) );
na03f02 TIMEBOOST_cell_34858 ( .a(TIMEBOOST_net_9430), .b(FE_OFN1374_n_8567), .c(g57038_sb), .o(n_11695) );
na02s01 g58352_u2 ( .a(FE_OFN1666_n_9477), .b(FE_OFN221_n_9846), .o(g58352_db) );
ao12f02 g55026_u0 ( .a(n_12430), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q), .o(n_12699) );
na04f04 TIMEBOOST_cell_24430 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .b(g58617_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_), .d(FE_OFN1369_n_8567), .o(n_9185) );
na04f04 TIMEBOOST_cell_24432 ( .a(n_9718), .b(g57216_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q), .d(FE_OFN1376_n_8567), .o(n_11542) );
ao12f02 g55031_u0 ( .a(n_12266), .b(FE_OFN1761_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q), .o(n_12695) );
na02f01 TIMEBOOST_cell_53334 ( .a(TIMEBOOST_net_16884), .b(g65212_db), .o(n_2676) );
na02s01 g58345_u2 ( .a(FE_OFN1666_n_9477), .b(FE_OFN211_n_9858), .o(g58345_db) );
ao12f02 g55034_u0 ( .a(n_12264), .b(FE_OFN1558_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q), .o(n_12693) );
na03f02 TIMEBOOST_cell_34783 ( .a(TIMEBOOST_net_9528), .b(FE_OFN1391_n_8567), .c(g57455_sb), .o(n_11279) );
na04f04 TIMEBOOST_cell_24434 ( .a(n_9685), .b(g57246_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q), .d(FE_OFN1408_n_8567), .o(n_11510) );
na02m02 TIMEBOOST_cell_37975 ( .a(TIMEBOOST_net_10599), .b(g64178_sb), .o(n_3988) );
na04f04 TIMEBOOST_cell_24268 ( .a(n_9583), .b(g57346_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q), .d(FE_OFN1384_n_8567), .o(n_11405) );
ao12f02 g55042_u0 ( .a(n_12258), .b(FE_OFN1760_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q), .o(n_12688) );
na02s01 g58328_u2 ( .a(FE_OFN239_n_9832), .b(FE_OFN572_n_9502), .o(g58328_db) );
na02f01 TIMEBOOST_cell_44370 ( .a(TIMEBOOST_net_13079), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_11410) );
na02s01 g58327_u2 ( .a(FE_OFN235_n_9834), .b(FE_OFN572_n_9502), .o(g58327_db) );
ao12f02 g55050_u0 ( .a(n_12382), .b(FE_OFN1757_n_12681), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q), .o(n_12682) );
na04f02 TIMEBOOST_cell_73208 ( .a(FE_OFN2022_n_4778), .b(TIMEBOOST_net_16657), .c(TIMEBOOST_net_639), .d(g63598_sb), .o(n_7177) );
na02f02 TIMEBOOST_cell_71069 ( .a(TIMEBOOST_net_22742), .b(g62669_sb), .o(n_6200) );
na04f04 TIMEBOOST_cell_24436 ( .a(n_9462), .b(g57501_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q), .d(FE_OFN1415_n_8567), .o(n_11236) );
na03f02 TIMEBOOST_cell_34859 ( .a(TIMEBOOST_net_9563), .b(FE_OFN1411_n_8567), .c(g57408_sb), .o(n_11336) );
ao12f02 g55055_u0 ( .a(n_12475), .b(FE_OFN1553_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q), .o(n_12792) );
na04f04 TIMEBOOST_cell_24270 ( .a(n_9584), .b(g57343_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q), .d(FE_OFN1385_n_8567), .o(n_11406) );
ao12m01 g55058_u0 ( .a(n_11964), .b(FE_OFN1562_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q), .o(n_12503) );
in01f02 g55059_u0 ( .a(n_12501), .o(n_12677) );
na02s01 TIMEBOOST_cell_53450 ( .a(TIMEBOOST_net_16942), .b(g58050_db), .o(TIMEBOOST_net_9577) );
na02s02 TIMEBOOST_cell_47921 ( .a(g58163_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q), .o(TIMEBOOST_net_14178) );
na02f02 TIMEBOOST_cell_72301 ( .a(TIMEBOOST_net_23358), .b(g62648_sb), .o(n_6252) );
na04f04 TIMEBOOST_cell_24444 ( .a(n_9826), .b(g57103_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q), .d(FE_OFN1425_n_8567), .o(n_11642) );
na04f04 TIMEBOOST_cell_67632 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q), .b(g62894_sb), .c(TIMEBOOST_net_15242), .d(FE_OFN1202_n_4090), .o(n_6089) );
na03f04 TIMEBOOST_cell_73209 ( .a(TIMEBOOST_net_7265), .b(FE_OFN1149_n_13249), .c(TIMEBOOST_net_22365), .o(n_13668) );
ao12f02 g55066_u0 ( .a(n_12455), .b(FE_OFN1563_n_12502), .c(n_7373), .o(n_12791) );
na03f06 TIMEBOOST_cell_73210 ( .a(TIMEBOOST_net_16955), .b(FE_OFN1147_n_13249), .c(g54144_sb), .o(n_13495) );
na04f04 TIMEBOOST_cell_24450 ( .a(n_9798), .b(g57124_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q), .d(FE_OFN1419_n_8567), .o(n_11622) );
na02m02 TIMEBOOST_cell_68638 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q), .b(g64878_sb), .o(TIMEBOOST_net_21527) );
na02f01 TIMEBOOST_cell_68245 ( .a(TIMEBOOST_net_21330), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_12914) );
na02f04 TIMEBOOST_cell_44040 ( .a(TIMEBOOST_net_12914), .b(FE_OFN1147_n_13249), .o(TIMEBOOST_net_11493) );
na04f04 TIMEBOOST_cell_35124 ( .a(n_9299), .b(n_10124), .c(n_9298), .d(n_10127), .o(n_12155) );
na04f04 TIMEBOOST_cell_73211 ( .a(TIMEBOOST_net_20878), .b(FE_OFN1149_n_13249), .c(n_2100), .d(g54238_sb), .o(n_13650) );
ao12f02 g55078_u0 ( .a(n_12452), .b(FE_OFN1564_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q), .o(n_12789) );
na04f04 TIMEBOOST_cell_24272 ( .a(n_9589), .b(g57339_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q), .d(FE_OFN1425_n_8567), .o(n_11413) );
na03f02 TIMEBOOST_cell_35125 ( .a(TIMEBOOST_net_5572), .b(n_10792), .c(n_10281), .o(n_12169) );
ao12f02 g55081_u0 ( .a(n_12429), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q), .o(n_12662) );
na02s01 TIMEBOOST_cell_44041 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q), .b(g58419_sb), .o(TIMEBOOST_net_12915) );
na04f04 TIMEBOOST_cell_24460 ( .a(n_9467), .b(g57495_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q), .d(FE_OFN1424_n_8567), .o(n_11242) );
na03m02 TIMEBOOST_cell_72834 ( .a(g65328_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q), .c(TIMEBOOST_net_10577), .o(TIMEBOOST_net_17081) );
na02f02 g58311_u2 ( .a(FE_OFN572_n_9502), .b(FE_OFN211_n_9858), .o(g58311_db) );
na02s01 TIMEBOOST_cell_53328 ( .a(TIMEBOOST_net_16881), .b(g54216_da), .o(TIMEBOOST_net_13449) );
na04f02 TIMEBOOST_cell_35126 ( .a(n_10029), .b(n_10916), .c(n_10617), .d(n_12440), .o(n_12773) );
na03s02 TIMEBOOST_cell_68346 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(FE_OFN1785_n_1699), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q), .o(TIMEBOOST_net_21381) );
na02s01 TIMEBOOST_cell_31091 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_9650) );
na02f02 TIMEBOOST_cell_53206 ( .a(TIMEBOOST_net_16820), .b(g61914_sb), .o(n_7993) );
ao12f02 g55095_u0 ( .a(n_12073), .b(FE_OCP_RBN2272_n_10268), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q), .o(n_12495) );
na04m06 TIMEBOOST_cell_72963 ( .a(TIMEBOOST_net_14540), .b(FE_OFN1810_n_4454), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q), .d(g65064_sb), .o(TIMEBOOST_net_17515) );
na04f02 TIMEBOOST_cell_35127 ( .a(n_10880), .b(n_10881), .c(n_11720), .d(n_12564), .o(n_12826) );
na03f02 TIMEBOOST_cell_66858 ( .a(TIMEBOOST_net_20664), .b(n_14971), .c(g58654_sb), .o(n_9235) );
ao12f02 g55100_u0 ( .a(n_12474), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q), .o(n_12787) );
na02s01 g58305_u2 ( .a(FE_OFN252_n_9868), .b(FE_OFN569_n_9528), .o(g58305_db) );
na04f04 TIMEBOOST_cell_24466 ( .a(n_9472), .b(g57488_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q), .d(FE_OFN1408_n_8567), .o(n_11249) );
na02s02 TIMEBOOST_cell_68500 ( .a(TIMEBOOST_net_20755), .b(g65784_sb), .o(TIMEBOOST_net_21458) );
na04f04 TIMEBOOST_cell_24468 ( .a(n_9475), .b(g57484_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q), .d(FE_OFN1415_n_8567), .o(n_11252) );
na02s01 TIMEBOOST_cell_44042 ( .a(TIMEBOOST_net_12915), .b(g58419_db), .o(n_9430) );
na02f02 TIMEBOOST_cell_70547 ( .a(TIMEBOOST_net_22481), .b(g62744_sb), .o(n_6135) );
ao12f02 g55108_u0 ( .a(n_12451), .b(FE_OFN1556_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q), .o(n_12786) );
ao12f02 g55110_u0 ( .a(n_12425), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q), .o(n_12642) );
na04m02 TIMEBOOST_cell_67324 ( .a(g65006_sb), .b(n_4479), .c(TIMEBOOST_net_12494), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q), .o(TIMEBOOST_net_20981) );
na02s02 TIMEBOOST_cell_48787 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q), .b(g58353_sb), .o(TIMEBOOST_net_14611) );
na02m02 TIMEBOOST_cell_68987 ( .a(TIMEBOOST_net_21701), .b(FE_OFN642_n_4677), .o(TIMEBOOST_net_12641) );
ao12f02 g55116_u0 ( .a(n_12450), .b(FE_OFN1564_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q), .o(n_12785) );
na04f04 TIMEBOOST_cell_24476 ( .a(n_9480), .b(g57479_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q), .d(FE_OFN1408_n_8567), .o(n_11258) );
na02s01 TIMEBOOST_cell_18155 ( .a(FE_OFN1780_parchk_pci_ad_reg_in_1221), .b(g65968_db), .o(TIMEBOOST_net_5441) );
na02s02 TIMEBOOST_cell_51952 ( .a(TIMEBOOST_net_16193), .b(g65731_sb), .o(n_1936) );
na02f02 TIMEBOOST_cell_54428 ( .a(TIMEBOOST_net_17431), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_15440) );
na03f01 TIMEBOOST_cell_65136 ( .a(n_3785), .b(FE_OFN1624_n_4438), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q), .o(TIMEBOOST_net_14398) );
na03f02 TIMEBOOST_cell_72626 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q), .c(TIMEBOOST_net_8679), .o(TIMEBOOST_net_17483) );
na04f04 g55132_u0 ( .a(n_10956), .b(n_9296), .c(n_10120), .d(n_9297), .o(n_12154) );
na02s01 TIMEBOOST_cell_18154 ( .a(TIMEBOOST_net_5440), .b(g65813_sb), .o(n_2576) );
na02s01 TIMEBOOST_cell_18143 ( .a(pci_target_unit_del_sync_be_out_reg_3__Q), .b(FE_OFN786_n_2678), .o(TIMEBOOST_net_5435) );
na04f04 g55136_u0 ( .a(n_9284), .b(n_9285), .c(n_10093), .d(n_10090), .o(n_12151) );
na02s02 TIMEBOOST_cell_51312 ( .a(TIMEBOOST_net_15873), .b(TIMEBOOST_net_11031), .o(TIMEBOOST_net_9464) );
na02s01 TIMEBOOST_cell_43161 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q), .o(TIMEBOOST_net_12475) );
na03m02 TIMEBOOST_cell_69796 ( .a(g65057_sb), .b(g65057_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q), .o(TIMEBOOST_net_22106) );
na02s01 TIMEBOOST_cell_52891 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q), .b(FE_OFN540_n_9690), .o(TIMEBOOST_net_16663) );
na03m02 TIMEBOOST_cell_72624 ( .a(g64829_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q), .c(TIMEBOOST_net_10393), .o(TIMEBOOST_net_17066) );
na02s01 TIMEBOOST_cell_18149 ( .a(pci_target_unit_del_sync_be_out_reg_0__Q), .b(FE_OFN786_n_2678), .o(TIMEBOOST_net_5438) );
na04f04 TIMEBOOST_cell_24843 ( .a(wbs_dat_o_25_), .b(g52520_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_124), .d(FE_OFN2242_g52675_p), .o(n_13738) );
na04f04 TIMEBOOST_cell_24842 ( .a(wbs_dat_o_1_), .b(g52514_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_100), .d(FE_OFN2243_g52675_p), .o(n_13809) );
na02m10 TIMEBOOST_cell_44449 ( .a(g58350_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q), .o(TIMEBOOST_net_13119) );
na03f02 TIMEBOOST_cell_24837 ( .a(n_14895), .b(n_13484), .c(n_14829), .o(n_14893) );
na02s01 TIMEBOOST_cell_63088 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q), .o(TIMEBOOST_net_20491) );
na02m02 TIMEBOOST_cell_69820 ( .a(g64834_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_22118) );
na02s01 TIMEBOOST_cell_52631 ( .a(n_366), .b(n_271), .o(TIMEBOOST_net_16533) );
ao12f02 g55161_u0 ( .a(n_12212), .b(FE_OFN1759_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q), .o(n_12632) );
na04f04 TIMEBOOST_cell_73693 ( .a(n_10575), .b(n_10572), .c(n_9988), .d(n_9992), .o(n_12135) );
na02s01 g58265_u2 ( .a(FE_OFN239_n_9832), .b(FE_OFN1649_n_9428), .o(g58265_db) );
na02f06 FE_RC_883_0 ( .a(wishbone_slave_unit_pcim_sm_data_in_658), .b(FE_OFN1611_n_2122), .o(FE_RN_579_0) );
na04f04 TIMEBOOST_cell_24478 ( .a(n_8996), .b(g57575_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q), .d(FE_OFN1389_n_8567), .o(n_10294) );
na02m10 TIMEBOOST_cell_45627 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q), .o(TIMEBOOST_net_13708) );
na03f02 TIMEBOOST_cell_33373 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_790), .b(g54314_sb), .c(g54314_db), .o(n_13102) );
na04m04 TIMEBOOST_cell_24486 ( .a(n_9106), .b(g57134_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q), .d(FE_OFN1396_n_8567), .o(n_10469) );
na02f02 TIMEBOOST_cell_70999 ( .a(TIMEBOOST_net_22707), .b(g62598_sb), .o(n_6355) );
na02s01 g65679_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q), .b(FE_OFN941_n_2047), .o(g65679_db) );
na04f04 TIMEBOOST_cell_24492 ( .a(n_9455), .b(g57515_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q), .d(FE_OFN1425_n_8567), .o(n_11226) );
ao12f02 g55179_u0 ( .a(n_12449), .b(FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q), .o(n_12781) );
na03m02 TIMEBOOST_cell_64409 ( .a(TIMEBOOST_net_17197), .b(FE_OFN936_n_2292), .c(g65687_sb), .o(n_2293) );
ao12f02 g55182_u0 ( .a(n_12423), .b(FE_OFN1552_n_12104), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q), .o(n_12619) );
na03m03 TIMEBOOST_cell_68654 ( .a(TIMEBOOST_net_21165), .b(g65671_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q), .o(TIMEBOOST_net_21535) );
na02m02 g65709_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q), .b(FE_OFN2109_n_2047), .o(g65709_db) );
ao12f02 g55187_u0 ( .a(n_12448), .b(FE_OFN1565_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q), .o(n_12780) );
na02s01 TIMEBOOST_cell_42771 ( .a(g54219_sb), .b(TIMEBOOST_net_6807), .o(TIMEBOOST_net_12280) );
na03m06 TIMEBOOST_cell_68898 ( .a(TIMEBOOST_net_13877), .b(g65888_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q), .o(TIMEBOOST_net_21657) );
na02s01 TIMEBOOST_cell_50018 ( .a(TIMEBOOST_net_15226), .b(TIMEBOOST_net_11461), .o(TIMEBOOST_net_9362) );
na03f02 TIMEBOOST_cell_65942 ( .a(TIMEBOOST_net_17306), .b(FE_OFN1171_n_5592), .c(g62131_sb), .o(n_5565) );
na02s02 TIMEBOOST_cell_68280 ( .a(g65789_sb), .b(TIMEBOOST_net_21169), .o(TIMEBOOST_net_21348) );
ao12f04 g55193_u0 ( .a(n_12447), .b(FE_OCP_RBN2013_FE_OCPN1895_FE_OFN1559_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q), .o(n_12779) );
ao12f02 g55196_u0 ( .a(n_11891), .b(FE_OFN1565_n_12502), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q), .o(n_12484) );
na02m04 TIMEBOOST_cell_49235 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_), .o(TIMEBOOST_net_14835) );
na02m01 TIMEBOOST_cell_68456 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q), .b(FE_OFN671_n_4505), .o(TIMEBOOST_net_21436) );
na02s01 TIMEBOOST_cell_62876 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q), .o(TIMEBOOST_net_20385) );
na03s02 TIMEBOOST_cell_32811 ( .a(n_2300), .b(g62003_sb), .c(g62003_db), .o(n_7889) );
na03m02 TIMEBOOST_cell_72510 ( .a(g65879_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q), .c(TIMEBOOST_net_14117), .o(TIMEBOOST_net_17009) );
na04f04 TIMEBOOST_cell_24278 ( .a(n_9593), .b(g57332_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q), .d(FE_OFN1417_n_8567), .o(n_11418) );
ao12f02 g55204_u0 ( .a(n_12186), .b(FE_OFN1760_n_10780), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q), .o(n_12602) );
na02f02 TIMEBOOST_cell_44623 ( .a(n_4160), .b(FE_OFN1700_n_5751), .o(TIMEBOOST_net_13206) );
na04f04 TIMEBOOST_cell_24506 ( .a(n_9796), .b(g57125_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q), .d(FE_OFN1415_n_8567), .o(n_11620) );
na04f04 TIMEBOOST_cell_24508 ( .a(n_9534), .b(g57584_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q), .d(FE_OFN1396_n_8567), .o(n_11165) );
na03s01 TIMEBOOST_cell_41741 ( .a(g58409_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q), .c(g58409_db), .o(n_9431) );
ao12f02 g55212_u0 ( .a(n_11885), .b(FE_OFN1749_n_12004), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q), .o(n_12480) );
no02f04 g55217_u0 ( .a(n_15001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56), .o(n_12479) );
na03f02 TIMEBOOST_cell_67951 ( .a(TIMEBOOST_net_13113), .b(FE_OFN1132_g64577_p), .c(g62736_sb), .o(n_5507) );
na02m01 TIMEBOOST_cell_68304 ( .a(TIMEBOOST_net_6803), .b(n_4725), .o(TIMEBOOST_net_21360) );
no02f04 g55221_u0 ( .a(n_15001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59), .o(n_12478) );
na02m02 TIMEBOOST_cell_69399 ( .a(TIMEBOOST_net_21907), .b(g64952_sb), .o(TIMEBOOST_net_17573) );
na02f02 TIMEBOOST_cell_51260 ( .a(TIMEBOOST_net_15847), .b(g61760_sb), .o(n_8293) );
no02f01 g55224_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62), .o(n_12476) );
na03f04 TIMEBOOST_cell_66657 ( .a(TIMEBOOST_net_17096), .b(FE_OFN1313_n_6624), .c(g62433_sb), .o(n_6731) );
na03s02 TIMEBOOST_cell_73495 ( .a(FE_OFN231_n_9839), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q), .c(FE_OFN1687_n_9528), .o(TIMEBOOST_net_20642) );
na02f02 g55228_u0 ( .a(FE_OCPN1827_n_14995), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q), .o(n_12122) );
no02f02 g55229_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67), .o(n_12430) );
na03s02 TIMEBOOST_cell_32815 ( .a(n_2161), .b(g61999_sb), .c(g61999_db), .o(n_7897) );
no02f04 g55233_u0 ( .a(n_15001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70), .o(n_12475) );
na02f02 g55234_u0 ( .a(FE_OCP_RBN1979_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q), .o(n_12117) );
na03m02 TIMEBOOST_cell_73212 ( .a(TIMEBOOST_net_22253), .b(FE_OFN1095_g64577_p), .c(g63077_sb), .o(n_7121) );
no02f01 g55237_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43), .o(n_12429) );
na02m01 TIMEBOOST_cell_52275 ( .a(TIMEBOOST_net_12703), .b(FE_OFN1049_n_16657), .o(TIMEBOOST_net_16355) );
no02f04 TIMEBOOST_cell_18039 ( .a(FE_RN_621_0), .b(FE_RN_609_0), .o(TIMEBOOST_net_5383) );
no02f02 g55240_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46), .o(n_12474) );
no02f01 g55241_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47), .o(n_12425) );
na03f01 TIMEBOOST_cell_68366 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q), .c(FE_OFN906_n_4736), .o(TIMEBOOST_net_21391) );
na02f02 TIMEBOOST_cell_43646 ( .a(TIMEBOOST_net_12717), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_11002) );
na03m02 TIMEBOOST_cell_68972 ( .a(TIMEBOOST_net_14229), .b(FE_OFN1013_n_4734), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q), .o(TIMEBOOST_net_21694) );
na03s02 TIMEBOOST_cell_72538 ( .a(g58160_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q), .c(g58166_db), .o(TIMEBOOST_net_16421) );
no02f02 g55246_u0 ( .a(FE_OCP_RBN1922_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51), .o(n_12423) );
na02f02 g55247_u0 ( .a(FE_OCP_RBN1924_n_10273), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q), .o(n_12112) );
na02m02 TIMEBOOST_cell_47885 ( .a(n_3747), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q), .o(TIMEBOOST_net_14160) );
na03f02 TIMEBOOST_cell_66955 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_16010), .c(FE_OFN2210_n_11027), .o(n_12621) );
na03f02 TIMEBOOST_cell_66719 ( .a(TIMEBOOST_net_17095), .b(FE_OFN1312_n_6624), .c(g62673_sb), .o(n_6193) );
na02s01 TIMEBOOST_cell_47920 ( .a(TIMEBOOST_net_14177), .b(FE_OFN950_n_2055), .o(TIMEBOOST_net_12490) );
na02m01 TIMEBOOST_cell_70131 ( .a(TIMEBOOST_net_22273), .b(FE_OFN577_n_9902), .o(TIMEBOOST_net_20404) );
na03f02 TIMEBOOST_cell_73769 ( .a(TIMEBOOST_net_13701), .b(FE_OFN1774_n_13800), .c(FE_OFN1770_n_14054), .o(g53203_p) );
na03s02 TIMEBOOST_cell_73047 ( .a(TIMEBOOST_net_23230), .b(FE_OFN707_n_8119), .c(g61926_sb), .o(n_7971) );
na02m02 TIMEBOOST_cell_51304 ( .a(TIMEBOOST_net_15869), .b(g63001_sb), .o(n_5880) );
na04f04 TIMEBOOST_cell_24375 ( .a(n_9407), .b(g57580_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q), .d(FE_OFN1389_n_8567), .o(n_11171) );
no02f02 g55257_u0 ( .a(n_12381), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330), .o(n_12417) );
na03f02 TIMEBOOST_cell_66518 ( .a(TIMEBOOST_net_16807), .b(FE_OFN1333_n_13547), .c(g53912_sb), .o(n_13529) );
na04m02 TIMEBOOST_cell_67268 ( .a(n_3741), .b(g65004_sb), .c(g65004_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q), .o(TIMEBOOST_net_21022) );
na02f02 TIMEBOOST_cell_50194 ( .a(TIMEBOOST_net_15314), .b(g60661_sb), .o(n_5658) );
na03m02 TIMEBOOST_cell_64408 ( .a(TIMEBOOST_net_17198), .b(FE_OFN936_n_2292), .c(g65712_sb), .o(n_2198) );
na02m04 TIMEBOOST_cell_54061 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q), .o(TIMEBOOST_net_17248) );
na03m04 TIMEBOOST_cell_72402 ( .a(n_817), .b(n_1283), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_), .o(TIMEBOOST_net_22257) );
in01s04 TIMEBOOST_cell_67100 ( .a(TIMEBOOST_net_21134), .o(FE_OFN518_n_9697) );
na02s01 TIMEBOOST_cell_48321 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_14378) );
na02f02 TIMEBOOST_cell_70039 ( .a(TIMEBOOST_net_22227), .b(g61823_sb), .o(n_8142) );
na02m02 TIMEBOOST_cell_52292 ( .a(TIMEBOOST_net_16363), .b(g65431_sb), .o(n_3506) );
na02f02 TIMEBOOST_cell_44381 ( .a(n_3852), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q), .o(TIMEBOOST_net_13085) );
na02m01 TIMEBOOST_cell_31511 ( .a(g64852_sb), .b(n_4482), .o(TIMEBOOST_net_9860) );
na03s02 TIMEBOOST_cell_72543 ( .a(FE_OFN563_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q), .c(TIMEBOOST_net_12793), .o(TIMEBOOST_net_16455) );
na03f02 TIMEBOOST_cell_72742 ( .a(TIMEBOOST_net_21573), .b(g64296_sb), .c(FE_OFN2106_g64577_p), .o(TIMEBOOST_net_22543) );
na03f02 TIMEBOOST_cell_65357 ( .a(TIMEBOOST_net_16313), .b(n_5633), .c(g62078_sb), .o(n_5632) );
na02s01 TIMEBOOST_cell_52633 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_16534) );
na03m02 TIMEBOOST_cell_72759 ( .a(TIMEBOOST_net_21538), .b(g64987_sb), .c(TIMEBOOST_net_21848), .o(TIMEBOOST_net_13237) );
in01f04 TIMEBOOST_cell_35476 ( .a(TIMEBOOST_net_10067), .o(n_7608) );
na04f01 TIMEBOOST_cell_67941 ( .a(n_3939), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q), .c(FE_OFN1134_g64577_p), .d(g63017_sb), .o(n_5214) );
na02m02 TIMEBOOST_cell_38695 ( .a(TIMEBOOST_net_10959), .b(g64091_sb), .o(n_4064) );
na02s01 TIMEBOOST_cell_50029 ( .a(configuration_pci_err_addr_489), .b(wbm_adr_o_19_), .o(TIMEBOOST_net_15232) );
na04f04 TIMEBOOST_cell_24415 ( .a(n_9732), .b(g57195_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q), .d(FE_OFN1385_n_8567), .o(n_11557) );
na02f02 g55292_u0 ( .a(FE_OFN1553_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q), .o(n_12393) );
na03f02 TIMEBOOST_cell_66646 ( .a(TIMEBOOST_net_17081), .b(FE_OFN2063_n_6391), .c(g62953_sb), .o(n_5975) );
na04f04 TIMEBOOST_cell_24419 ( .a(n_9024), .b(g57458_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q), .d(FE_OFN1385_n_8567), .o(n_10346) );
na02s01 TIMEBOOST_cell_62478 ( .a(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .b(g54171_sb), .o(TIMEBOOST_net_20186) );
na02s02 TIMEBOOST_cell_49083 ( .a(g58387_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q), .o(TIMEBOOST_net_14759) );
na02f02 TIMEBOOST_cell_68217 ( .a(TIMEBOOST_net_21316), .b(n_580), .o(TIMEBOOST_net_20667) );
na04f04 TIMEBOOST_cell_24423 ( .a(n_9498), .b(g57452_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q), .d(FE_OFN1408_n_8567), .o(n_11282) );
na02f02 g55299_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q), .o(n_12088) );
na04f04 TIMEBOOST_cell_24427 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .b(g58619_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_), .d(FE_OFN1369_n_8567), .o(n_9183) );
na02m02 TIMEBOOST_cell_50027 ( .a(wbm_adr_o_23_), .b(configuration_pci_err_addr_493), .o(TIMEBOOST_net_15231) );
na02m01 TIMEBOOST_cell_53997 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q), .o(TIMEBOOST_net_17216) );
na02f01 g55303_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q), .o(n_12084) );
na03s02 TIMEBOOST_cell_73281 ( .a(TIMEBOOST_net_22262), .b(n_8272), .c(g61893_sb), .o(n_8041) );
na02m04 TIMEBOOST_cell_68830 ( .a(n_4488), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q), .o(TIMEBOOST_net_21623) );
na03f02 TIMEBOOST_cell_66325 ( .a(TIMEBOOST_net_9947), .b(n_6287), .c(g62495_sb), .o(n_6594) );
no02f02 g55310_u0 ( .a(n_12381), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342), .o(n_12382) );
na02s01 TIMEBOOST_cell_53103 ( .a(g58115_sb), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_16769) );
na03m20 TIMEBOOST_cell_69580 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(FE_OFN918_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q), .o(TIMEBOOST_net_21998) );
na04f04 TIMEBOOST_cell_24431 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .b(g58616_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_), .d(FE_OFN1369_n_8567), .o(n_9187) );
na02f02 g55314_u0 ( .a(FE_OFN1551_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q), .o(n_12379) );
na02f04 g55315_u0 ( .a(FE_OCP_RBN1975_n_12381), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q), .o(n_12378) );
na03m02 TIMEBOOST_cell_73048 ( .a(TIMEBOOST_net_22044), .b(FE_OFN706_n_8119), .c(g61954_sb), .o(n_7917) );
na02m01 TIMEBOOST_cell_48682 ( .a(TIMEBOOST_net_14558), .b(FE_OFN912_n_4727), .o(TIMEBOOST_net_12839) );
na03m02 TIMEBOOST_cell_72995 ( .a(TIMEBOOST_net_21920), .b(g65017_sb), .c(TIMEBOOST_net_22086), .o(TIMEBOOST_net_17458) );
na03f02 TIMEBOOST_cell_66184 ( .a(TIMEBOOST_net_16731), .b(FE_OFN1182_n_3476), .c(g60621_sb), .o(n_4833) );
na03f02 TIMEBOOST_cell_65932 ( .a(TIMEBOOST_net_8786), .b(FE_OFN1169_n_5592), .c(g62109_sb), .o(n_5589) );
na02f01 TIMEBOOST_cell_70586 ( .a(TIMEBOOST_net_15073), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_22501) );
na03f02 TIMEBOOST_cell_66170 ( .a(TIMEBOOST_net_16440), .b(FE_OFN1184_n_3476), .c(g60617_sb), .o(n_4837) );
na04f04 TIMEBOOST_cell_24644 ( .a(n_9077), .b(g57249_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q), .d(FE_OFN2180_n_8567), .o(n_10423) );
na02s01 TIMEBOOST_cell_47726 ( .a(TIMEBOOST_net_14080), .b(FE_OFN602_n_9687), .o(TIMEBOOST_net_10229) );
na04f04 TIMEBOOST_cell_24437 ( .a(n_9683), .b(g57250_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q), .d(FE_OFN1384_n_8567), .o(n_11507) );
na03f02 TIMEBOOST_cell_66957 ( .a(FE_OFN1752_n_12086), .b(TIMEBOOST_net_16507), .c(FE_OFN2209_n_11027), .o(n_12758) );
na02s01 TIMEBOOST_cell_52635 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q), .o(TIMEBOOST_net_16535) );
na02m02 TIMEBOOST_cell_64091 ( .a(TIMEBOOST_net_21031), .b(g58079_sb), .o(TIMEBOOST_net_20602) );
na02f02 g55332_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q), .o(n_12075) );
na02m02 TIMEBOOST_cell_70023 ( .a(TIMEBOOST_net_22219), .b(g62027_sb), .o(n_7842) );
no02f02 g55335_u0 ( .a(FE_OCPN1907_n_11767), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6), .o(n_12073) );
na02f02 g55336_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q), .o(n_12072) );
in01f02 TIMEBOOST_cell_35477 ( .a(TIMEBOOST_net_10068), .o(TIMEBOOST_net_10067) );
na02m08 TIMEBOOST_cell_53035 ( .a(configuration_pci_err_addr_488), .b(wbm_adr_o_18_), .o(TIMEBOOST_net_16735) );
na03f02 TIMEBOOST_cell_67882 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(g64184_sb), .c(g64184_db), .o(n_3982) );
na03s02 TIMEBOOST_cell_46689 ( .a(TIMEBOOST_net_12774), .b(g58238_sb), .c(g58248_db), .o(TIMEBOOST_net_9344) );
na02m02 TIMEBOOST_cell_69865 ( .a(TIMEBOOST_net_22140), .b(g64256_sb), .o(n_3917) );
na02f02 g55346_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q), .o(n_12068) );
no03f10 TIMEBOOST_cell_64381 ( .a(FE_RN_103_0), .b(FE_RN_102_0), .c(n_16030), .o(n_1279) );
na02s01 TIMEBOOST_cell_48436 ( .a(TIMEBOOST_net_14435), .b(FE_OFN517_n_9697), .o(TIMEBOOST_net_10620) );
na02s01 TIMEBOOST_cell_52213 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q), .b(g58278_sb), .o(TIMEBOOST_net_16324) );
na02s02 TIMEBOOST_cell_52214 ( .a(TIMEBOOST_net_16324), .b(g58278_db), .o(n_9524) );
na02f04 g55351_u0 ( .a(n_12357), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q), .o(n_12349) );
no03f10 TIMEBOOST_cell_23949 ( .a(n_15512), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_), .c(FE_RN_540_0), .o(n_15514) );
na03f20 TIMEBOOST_cell_23951 ( .a(g75162_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .c(g75162_db), .o(n_16534) );
na02f04 g55357_u0 ( .a(n_12357), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q), .o(n_12345) );
na02f02 g55358_u0 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q), .o(n_12066) );
na02f01 TIMEBOOST_cell_72226 ( .a(TIMEBOOST_net_9913), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_23321) );
in01s01 TIMEBOOST_cell_72352 ( .a(TIMEBOOST_net_23385), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_93) );
na02m02 TIMEBOOST_cell_39975 ( .a(TIMEBOOST_net_11599), .b(g62589_sb), .o(n_6373) );
na03m02 TIMEBOOST_cell_68586 ( .a(FE_OFN624_n_4409), .b(g64906_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q), .o(TIMEBOOST_net_21501) );
na02f02 g55364_u0 ( .a(FE_OFN1553_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q), .o(n_12341) );
na02m02 TIMEBOOST_cell_50562 ( .a(TIMEBOOST_net_15498), .b(g62927_sb), .o(n_6027) );
na03f02 TIMEBOOST_cell_66529 ( .a(TIMEBOOST_net_16799), .b(FE_OFN1331_n_13547), .c(g53928_sb), .o(n_13517) );
na02s03 TIMEBOOST_cell_52637 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q), .o(TIMEBOOST_net_16536) );
na04m06 TIMEBOOST_cell_65898 ( .a(g57955_db), .b(g57964_sb), .c(FE_OFN262_n_9851), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q), .o(TIMEBOOST_net_17172) );
na02m10 TIMEBOOST_cell_69586 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_143), .o(TIMEBOOST_net_22001) );
na02s01 TIMEBOOST_cell_48442 ( .a(TIMEBOOST_net_14438), .b(FE_OFN2254_n_9687), .o(TIMEBOOST_net_10610) );
na04s04 TIMEBOOST_cell_66272 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q), .b(FE_OFN231_n_9839), .c(FE_OFN584_n_9692), .d(g58185_sb), .o(n_9602) );
na02f02 TIMEBOOST_cell_54410 ( .a(TIMEBOOST_net_17422), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_15500) );
na02f02 g55382_u0 ( .a(FE_OCPN1825_n_12030), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q), .o(n_12055) );
na02f04 g55383_u0 ( .a(FE_OFN1565_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q), .o(n_12054) );
na02f02 g55384_u0 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q), .o(n_12053) );
na02f04 g55385_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q), .o(n_12052) );
na03f02 TIMEBOOST_cell_66861 ( .a(FE_OFN1565_n_12502), .b(TIMEBOOST_net_16477), .c(n_12313), .o(n_12726) );
na04f04 TIMEBOOST_cell_24379 ( .a(n_9437), .b(g57539_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q), .d(FE_OFN1396_n_8567), .o(n_11203) );
na02m10 TIMEBOOST_cell_51681 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_16058) );
na02m10 TIMEBOOST_cell_45713 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q), .o(TIMEBOOST_net_13751) );
na02s01 TIMEBOOST_cell_43574 ( .a(TIMEBOOST_net_12681), .b(FE_OFN1057_n_4727), .o(TIMEBOOST_net_10950) );
na03f02 TIMEBOOST_cell_72958 ( .a(TIMEBOOST_net_21820), .b(g65280_sb), .c(TIMEBOOST_net_22026), .o(TIMEBOOST_net_20963) );
no02f02 TIMEBOOST_cell_51519 ( .a(TIMEBOOST_net_7530), .b(FE_RN_711_0), .o(TIMEBOOST_net_15977) );
na02s02 TIMEBOOST_cell_54024 ( .a(TIMEBOOST_net_17229), .b(g57893_sb), .o(TIMEBOOST_net_14340) );
na02m10 TIMEBOOST_cell_45645 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q), .o(TIMEBOOST_net_13717) );
na02s01 TIMEBOOST_cell_62477 ( .a(TIMEBOOST_net_20185), .b(g54205_sb), .o(TIMEBOOST_net_14105) );
na03s02 TIMEBOOST_cell_66332 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q), .b(FE_OFN241_n_9830), .c(FE_OFN543_n_9690), .o(TIMEBOOST_net_10858) );
na02s01 TIMEBOOST_cell_43600 ( .a(TIMEBOOST_net_12694), .b(g58052_sb), .o(n_9093) );
na02f02 TIMEBOOST_cell_53606 ( .a(TIMEBOOST_net_17020), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_15533) );
na02f04 g55404_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q), .o(n_11841) );
na02s01 TIMEBOOST_cell_52639 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q), .o(TIMEBOOST_net_16537) );
no02f01 g55407_u0 ( .a(FE_OCPN1834_n_11884), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487), .o(n_12044) );
na03f04 TIMEBOOST_cell_66863 ( .a(FE_OFN1583_n_12306), .b(TIMEBOOST_net_13519), .c(FE_OFN1762_n_10780), .o(n_12754) );
na02s03 TIMEBOOST_cell_53225 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_768), .o(TIMEBOOST_net_16830) );
na02s01 TIMEBOOST_cell_53209 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_792), .o(TIMEBOOST_net_16822) );
na04f02 TIMEBOOST_cell_67908 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q), .b(FE_OFN716_n_8176), .c(n_1610), .d(g61811_sb), .o(n_8171) );
na02f04 g55415_u0 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q), .o(n_12038) );
na02f04 g55416_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q), .o(n_12310) );
na02f02 g55417_u0 ( .a(n_12001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q), .o(n_12037) );
na02f04 g55418_u0 ( .a(FE_OFN1749_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q), .o(n_12036) );
na02f02 TIMEBOOST_cell_39373 ( .a(TIMEBOOST_net_11298), .b(g63046_sb), .o(n_5161) );
in01s01 TIMEBOOST_cell_73871 ( .a(TIMEBOOST_net_23435), .o(TIMEBOOST_net_23436) );
in01s01 TIMEBOOST_cell_73940 ( .a(wbm_dat_i_20_), .o(TIMEBOOST_net_23505) );
in01s01 TIMEBOOST_cell_73855 ( .a(TIMEBOOST_net_23419), .o(TIMEBOOST_net_23420) );
na02f04 g55424_u0 ( .a(FE_OFN1566_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q), .o(n_12032) );
na02f04 g55425_u0 ( .a(FE_OCPN1825_n_12030), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q), .o(n_12031) );
na02s02 TIMEBOOST_cell_43604 ( .a(TIMEBOOST_net_12696), .b(g65720_sb), .o(n_1942) );
na03f02 TIMEBOOST_cell_66496 ( .a(TIMEBOOST_net_17134), .b(FE_OFN1312_n_6624), .c(g62955_sb), .o(n_5971) );
na02m02 TIMEBOOST_cell_50025 ( .a(wbm_adr_o_22_), .b(configuration_pci_err_addr_492), .o(TIMEBOOST_net_15230) );
na03s02 TIMEBOOST_cell_70022 ( .a(n_1838), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q), .c(FE_OFN699_n_7845), .o(TIMEBOOST_net_22219) );
na02m01 TIMEBOOST_cell_62602 ( .a(n_3749), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q), .o(TIMEBOOST_net_20248) );
na02m02 TIMEBOOST_cell_43606 ( .a(TIMEBOOST_net_12697), .b(g64145_sb), .o(n_4522) );
na04f02 TIMEBOOST_cell_24821 ( .a(n_10032), .b(n_10035), .c(n_9262), .d(n_9261), .o(n_11845) );
na02f01 TIMEBOOST_cell_40256 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_0__Q), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_11740) );
no02f04 g55439_u0 ( .a(n_12293), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177), .o(n_12300) );
na04f04 TIMEBOOST_cell_24397 ( .a(n_9098), .b(g57168_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q), .d(FE_OFN1396_n_8567), .o(n_10457) );
na03m02 TIMEBOOST_cell_72761 ( .a(n_4442), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q), .c(TIMEBOOST_net_10803), .o(TIMEBOOST_net_17061) );
na02m02 TIMEBOOST_cell_68374 ( .a(g65310_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q), .o(TIMEBOOST_net_21395) );
na02m04 TIMEBOOST_cell_69722 ( .a(g65349_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q), .o(TIMEBOOST_net_22069) );
na04m02 TIMEBOOST_cell_67900 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(FE_OFN1041_n_2037), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q), .d(g65869_sb), .o(n_1872) );
no02f04 g55449_u0 ( .a(n_12293), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178), .o(n_12294) );
na04s02 TIMEBOOST_cell_65029 ( .a(n_4493), .b(g65033_sb), .c(g65033_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_17058) );
na02s04 TIMEBOOST_cell_52641 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q), .o(TIMEBOOST_net_16538) );
na02m02 TIMEBOOST_cell_53372 ( .a(TIMEBOOST_net_16903), .b(FE_OFN1017_n_2053), .o(TIMEBOOST_net_14495) );
na03s02 TIMEBOOST_cell_73213 ( .a(TIMEBOOST_net_12810), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q), .c(FE_OFN531_n_9823), .o(TIMEBOOST_net_20879) );
na03f02 TIMEBOOST_cell_70002 ( .a(n_2056), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q), .c(FE_OFN717_n_8176), .o(TIMEBOOST_net_22209) );
na03f02 TIMEBOOST_cell_66910 ( .a(FE_OFN1733_n_16317), .b(TIMEBOOST_net_16486), .c(FE_OFN1738_n_11019), .o(n_12663) );
na02f02 TIMEBOOST_cell_70619 ( .a(TIMEBOOST_net_22517), .b(g62834_sb), .o(n_5305) );
na02m06 TIMEBOOST_cell_52259 ( .a(g64250_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q), .o(TIMEBOOST_net_16347) );
na02m06 TIMEBOOST_cell_49227 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q), .b(g65884_sb), .o(TIMEBOOST_net_14831) );
na02f02 TIMEBOOST_cell_52482 ( .a(TIMEBOOST_net_16458), .b(g62354_sb), .o(n_6892) );
na03f02 TIMEBOOST_cell_73594 ( .a(TIMEBOOST_net_13066), .b(FE_OFN1135_g64577_p), .c(g63064_sb), .o(n_5122) );
na03m02 TIMEBOOST_cell_72691 ( .a(TIMEBOOST_net_21528), .b(g65052_sb), .c(TIMEBOOST_net_21782), .o(TIMEBOOST_net_17131) );
no02f04 TIMEBOOST_cell_48464 ( .a(TIMEBOOST_net_14449), .b(FE_RN_581_0), .o(TIMEBOOST_net_7488) );
no02f01 g55468_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258), .o(n_12003) );
na02f02 g55469_u0 ( .a(n_12001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q), .o(n_12002) );
na02s01 TIMEBOOST_cell_70739 ( .a(TIMEBOOST_net_22577), .b(TIMEBOOST_net_12433), .o(TIMEBOOST_net_16432) );
na02m02 TIMEBOOST_cell_49084 ( .a(TIMEBOOST_net_14759), .b(g58387_db), .o(n_9444) );
na02s02 TIMEBOOST_cell_72303 ( .a(TIMEBOOST_net_23359), .b(g58212_sb), .o(n_9573) );
no02f02 g55474_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376), .o(n_12461) );
na02m08 TIMEBOOST_cell_45287 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q), .o(TIMEBOOST_net_13538) );
no02f04 g55477_u0 ( .a(n_16587), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532), .o(n_12280) );
na03m04 TIMEBOOST_cell_64407 ( .a(TIMEBOOST_net_17199), .b(FE_OFN935_n_2292), .c(g65772_sb), .o(n_2194) );
na03m02 TIMEBOOST_cell_72696 ( .a(TIMEBOOST_net_21565), .b(FE_OFN646_n_4497), .c(TIMEBOOST_net_21901), .o(TIMEBOOST_net_20533) );
na02f02 TIMEBOOST_cell_68367 ( .a(TIMEBOOST_net_21391), .b(g64197_sb), .o(n_3972) );
na03f02 TIMEBOOST_cell_66531 ( .a(g53913_sb), .b(FE_OFN1332_n_13547), .c(TIMEBOOST_net_16801), .o(n_13528) );
na04f04 TIMEBOOST_cell_24409 ( .a(n_9807), .b(g57116_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q), .d(FE_OFN1406_n_8567), .o(n_11630) );
na02s01 TIMEBOOST_cell_70738 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q), .b(FE_OFN1649_n_9428), .o(TIMEBOOST_net_22577) );
in01s01 TIMEBOOST_cell_72359 ( .a(TIMEBOOST_net_23391), .o(TIMEBOOST_net_23392) );
na02f01 g55487_u0 ( .a(n_11881), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q), .o(n_12276) );
na02f02 g55488_u0 ( .a(FE_OFN1562_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q), .o(n_11992) );
na02f02 g55489_u0 ( .a(FE_OFN2202_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q), .o(n_12275) );
na02f04 g55490_u0 ( .a(FE_OFN1577_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q), .o(n_12274) );
na02f02 g55491_u0 ( .a(FE_OFN1762_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q), .o(n_11991) );
na02f02 g55492_u0 ( .a(FE_OFN1583_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q), .o(n_11990) );
na03f02 TIMEBOOST_cell_64817 ( .a(TIMEBOOST_net_16900), .b(FE_OFN1011_n_4734), .c(g64163_sb), .o(TIMEBOOST_net_13048) );
no02f04 g55495_u0 ( .a(n_12293), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183), .o(n_12271) );
na02m02 TIMEBOOST_cell_68918 ( .a(n_4447), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q), .o(TIMEBOOST_net_21667) );
na04m02 TIMEBOOST_cell_67210 ( .a(n_3739), .b(g64781_sb), .c(g64781_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q), .o(TIMEBOOST_net_21002) );
na04f04 TIMEBOOST_cell_24417 ( .a(n_9459), .b(g57508_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q), .d(FE_OFN1402_n_8567), .o(n_11232) );
in01s01 TIMEBOOST_cell_73856 ( .a(n_14622), .o(TIMEBOOST_net_23421) );
no02f04 g55502_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__379), .o(n_12459) );
na03f04 TIMEBOOST_cell_65936 ( .a(TIMEBOOST_net_20443), .b(FE_OFN1174_n_5592), .c(g62141_sb), .o(n_5552) );
na02m01 TIMEBOOST_cell_4011 ( .a(TIMEBOOST_net_565), .b(g65858_db), .o(n_2594) );
na04f02 TIMEBOOST_cell_73496 ( .a(FE_OFN233_n_9876), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q), .c(FE_OFN580_n_9531), .d(g58393_sb), .o(n_9440) );
no02f04 g55512_u0 ( .a(FE_OCP_RBN2293_FE_OFN1581_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536), .o(n_12266) );
na02s01 TIMEBOOST_cell_49499 ( .a(FE_OFN264_n_9849), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q), .o(TIMEBOOST_net_14967) );
no02f04 g55515_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380), .o(n_12264) );
na03s02 TIMEBOOST_cell_68684 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q), .c(FE_OFN951_n_2055), .o(TIMEBOOST_net_21550) );
na02f02 TIMEBOOST_cell_49944 ( .a(TIMEBOOST_net_15189), .b(g62752_sb), .o(n_5476) );
na03m02 TIMEBOOST_cell_69316 ( .a(n_4465), .b(g65303_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q), .o(TIMEBOOST_net_21866) );
na03f04 TIMEBOOST_cell_66960 ( .a(FE_OCP_RBN1973_n_12381), .b(n_11831), .c(TIMEBOOST_net_16510), .o(n_12703) );
na02s02 TIMEBOOST_cell_43610 ( .a(TIMEBOOST_net_12699), .b(g65702_sb), .o(n_1949) );
na02m04 TIMEBOOST_cell_68680 ( .a(g64749_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q), .o(TIMEBOOST_net_21548) );
no02f04 g55524_u0 ( .a(n_11762), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509), .o(n_12258) );
na02f02 g55525_u0 ( .a(FE_OFN1762_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q), .o(n_11975) );
na02f02 g55526_u0 ( .a(FE_OFN1583_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q), .o(n_12257) );
na02m02 TIMEBOOST_cell_49500 ( .a(TIMEBOOST_net_14967), .b(TIMEBOOST_net_11211), .o(TIMEBOOST_net_9412) );
na03f04 TIMEBOOST_cell_73282 ( .a(TIMEBOOST_net_23312), .b(g63045_sb), .c(FE_OFN1120_g64577_p), .o(n_5163) );
na02f02 TIMEBOOST_cell_51180 ( .a(TIMEBOOST_net_15807), .b(g62950_sb), .o(n_5981) );
na04f04 TIMEBOOST_cell_24435 ( .a(n_9682), .b(g57251_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q), .d(FE_OFN1376_n_8567), .o(n_11505) );
na03f08 TIMEBOOST_cell_62810 ( .a(n_2435), .b(n_2428), .c(n_1359), .o(TIMEBOOST_net_20352) );
na02m01 TIMEBOOST_cell_68564 ( .a(FE_OFN622_n_4409), .b(n_4396), .o(TIMEBOOST_net_21490) );
na02m02 TIMEBOOST_cell_49239 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q), .b(g65314_sb), .o(TIMEBOOST_net_14837) );
na04m06 TIMEBOOST_cell_73149 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(FE_OFN923_n_4740), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q), .d(g64212_sb), .o(n_3957) );
na03f02 TIMEBOOST_cell_72784 ( .a(n_4488), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q), .c(TIMEBOOST_net_12548), .o(TIMEBOOST_net_20969) );
na04f04 TIMEBOOST_cell_24429 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .b(g58618_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_), .d(FE_OFN1369_n_8567), .o(n_9184) );
na02m02 TIMEBOOST_cell_68087 ( .a(TIMEBOOST_net_21251), .b(TIMEBOOST_net_6761), .o(TIMEBOOST_net_8810) );
na03m02 TIMEBOOST_cell_69854 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q), .b(TIMEBOOST_net_12679), .c(FE_OFN1056_n_4727), .o(TIMEBOOST_net_22135) );
no02f01 g55544_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__265), .o(n_11964) );
na02f04 g55545_u0 ( .a(FE_OFN1760_n_10780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q), .o(n_11962) );
na02f02 g55546_u0 ( .a(FE_OFN1579_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q), .o(n_11961) );
na02f02 g55547_u0 ( .a(FE_OFN2204_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q), .o(n_12248) );
na02f02 g55548_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q), .o(n_12246) );
na02f02 g55549_u0 ( .a(FE_OCPN1825_n_12030), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q), .o(n_11960) );
na02f02 g55550_u0 ( .a(FE_OFN1563_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q), .o(n_11819) );
na03f02 TIMEBOOST_cell_65916 ( .a(TIMEBOOST_net_17307), .b(FE_OFN1171_n_5592), .c(g62130_sb), .o(n_5566) );
na02f02 TIMEBOOST_cell_44856 ( .a(TIMEBOOST_net_13322), .b(g62528_sb), .o(n_6518) );
na02f04 g55553_u0 ( .a(n_11823), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q), .o(n_11818) );
na02f04 g55554_u0 ( .a(FE_OFN1748_n_12004), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q), .o(n_11957) );
na02f01 g55555_u0 ( .a(n_12001), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q), .o(n_11956) );
na03f02 TIMEBOOST_cell_66206 ( .a(TIMEBOOST_net_17003), .b(FE_OFN1276_n_4096), .c(g62914_sb), .o(n_6051) );
na02m04 TIMEBOOST_cell_72104 ( .a(g64193_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q), .o(TIMEBOOST_net_23260) );
na04f04 TIMEBOOST_cell_24439 ( .a(n_9818), .b(g57108_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q), .d(FE_OFN1415_n_8567), .o(n_11638) );
no02f04 g55561_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271), .o(n_12455) );
na02f02 g55562_u0 ( .a(FE_OFN1574_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q), .o(n_12244) );
na02f04 g55563_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q), .o(n_12243) );
na04f04 TIMEBOOST_cell_24441 ( .a(n_9820), .b(g57106_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q), .d(FE_OFN1423_n_8567), .o(n_11639) );
na03f02 TIMEBOOST_cell_65901 ( .a(n_4064), .b(g62848_sb), .c(g62848_db), .o(n_5275) );
na02m02 TIMEBOOST_cell_68876 ( .a(n_4672), .b(n_14), .o(TIMEBOOST_net_21646) );
na03f02 TIMEBOOST_cell_66964 ( .a(FE_OCPN1866_n_12377), .b(FE_OFN1757_n_12681), .c(TIMEBOOST_net_13675), .o(n_12604) );
na03f04 TIMEBOOST_cell_66959 ( .a(TIMEBOOST_net_13668), .b(n_11831), .c(n_12357), .o(n_12728) );
na02m01 TIMEBOOST_cell_68246 ( .a(n_8884), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q), .o(TIMEBOOST_net_21331) );
na03f02 TIMEBOOST_cell_66656 ( .a(TIMEBOOST_net_16771), .b(FE_OFN1315_n_6624), .c(g62569_sb), .o(n_6417) );
na02f04 g55572_u0 ( .a(FE_OFN1574_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q), .o(n_12238) );
na03m06 TIMEBOOST_cell_72403 ( .a(pci_target_unit_fifos_pcir_flush_in), .b(g57780_sb), .c(n_7569), .o(TIMEBOOST_net_21355) );
na03f02 TIMEBOOST_cell_72693 ( .a(TIMEBOOST_net_21529), .b(g65023_sb), .c(TIMEBOOST_net_22119), .o(TIMEBOOST_net_20955) );
na03m04 TIMEBOOST_cell_73119 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q), .b(g63563_sb), .c(TIMEBOOST_net_16959), .o(TIMEBOOST_net_14892) );
na02m02 TIMEBOOST_cell_68368 ( .a(g65373_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q), .o(TIMEBOOST_net_21392) );
na03s02 TIMEBOOST_cell_46605 ( .a(TIMEBOOST_net_12829), .b(g63613_sb), .c(g63613_db), .o(n_7143) );
no02f04 g55581_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238), .o(n_12452) );
na03f02 TIMEBOOST_cell_70576 ( .a(n_7218), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q), .c(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_22496) );
na04f04 TIMEBOOST_cell_24271 ( .a(n_9585), .b(g57342_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q), .d(FE_OFN1408_n_8567), .o(n_11408) );
na04f04 TIMEBOOST_cell_24453 ( .a(n_9003), .b(g57546_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q), .d(FE_OFN1396_n_8567), .o(n_10308) );
na02s02 TIMEBOOST_cell_69746 ( .a(FE_OFN215_n_9856), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q), .o(TIMEBOOST_net_22081) );
na04f04 TIMEBOOST_cell_35225 ( .a(n_17045), .b(n_9329), .c(n_17046), .d(n_9330), .o(n_12164) );
na03f02 TIMEBOOST_cell_66761 ( .a(n_4044), .b(g62734_sb), .c(g62734_db), .o(n_5511) );
na04f04 TIMEBOOST_cell_24459 ( .a(n_9466), .b(g57496_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q), .d(FE_OFN1424_n_8567), .o(n_11241) );
na02m04 TIMEBOOST_cell_69867 ( .a(TIMEBOOST_net_22141), .b(g64339_sb), .o(TIMEBOOST_net_17318) );
na04f04 TIMEBOOST_cell_24455 ( .a(n_9463), .b(g57500_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q), .d(FE_OFN1419_n_8567), .o(n_11238) );
in01s01 TIMEBOOST_cell_67751 ( .a(pci_target_unit_fifos_pcir_data_in_174), .o(TIMEBOOST_net_21178) );
na02f02 g55594_u0 ( .a(FE_OFN1739_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q), .o(n_11938) );
na02f04 g55595_u0 ( .a(FE_OFN1734_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q), .o(n_11937) );
na02f02 g55596_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q), .o(n_11814) );
na04f04 TIMEBOOST_cell_24275 ( .a(n_9057), .b(g57335_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q), .d(FE_OFN1416_n_8567), .o(n_10394) );
na04f04 TIMEBOOST_cell_35221 ( .a(n_9269), .b(n_10054), .c(n_9270), .d(n_10057), .o(n_12146) );
na03f02 TIMEBOOST_cell_65255 ( .a(TIMEBOOST_net_16290), .b(g64350_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q), .o(TIMEBOOST_net_15069) );
na02f02 TIMEBOOST_cell_51292 ( .a(TIMEBOOST_net_15863), .b(g63147_sb), .o(n_5846) );
na03f02 TIMEBOOST_cell_68548 ( .a(FE_OFN1001_n_15978), .b(conf_wb_err_bc_in_848), .c(n_211), .o(TIMEBOOST_net_21482) );
na02m02 TIMEBOOST_cell_37941 ( .a(TIMEBOOST_net_10582), .b(g58319_db), .o(n_9493) );
na03m02 TIMEBOOST_cell_72819 ( .a(g65300_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q), .c(TIMEBOOST_net_16265), .o(TIMEBOOST_net_20535) );
na02s02 TIMEBOOST_cell_38545 ( .a(TIMEBOOST_net_10884), .b(g58209_db), .o(n_9576) );
na03m02 TIMEBOOST_cell_68914 ( .a(n_4470), .b(g64775_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q), .o(TIMEBOOST_net_21665) );
in01s01 TIMEBOOST_cell_63606 ( .a(TIMEBOOST_net_20786), .o(TIMEBOOST_net_20741) );
na03f02 TIMEBOOST_cell_66308 ( .a(TIMEBOOST_net_13374), .b(n_6554), .c(g62511_sb), .o(n_6556) );
na04f04 TIMEBOOST_cell_24463 ( .a(n_9469), .b(g57492_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q), .d(FE_OFN1406_n_8567), .o(n_11244) );
na03s02 TIMEBOOST_cell_72694 ( .a(TIMEBOOST_net_21209), .b(g65730_sb), .c(TIMEBOOST_net_7094), .o(n_1981) );
na02s02 TIMEBOOST_cell_49532 ( .a(TIMEBOOST_net_14983), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_12949) );
na02s01 TIMEBOOST_cell_53911 ( .a(g58206_sb), .b(FE_RN_484_0), .o(TIMEBOOST_net_17173) );
no02f04 g55623_u0 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359), .o(n_12451) );
na02m02 TIMEBOOST_cell_68853 ( .a(TIMEBOOST_net_21634), .b(n_4442), .o(TIMEBOOST_net_20344) );
na04m04 TIMEBOOST_cell_36027 ( .a(g62013_sb), .b(n_2155), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q), .d(FE_OFN712_n_8140), .o(n_7869) );
na03f02 TIMEBOOST_cell_73792 ( .a(FE_OFN1602_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q), .c(n_17021), .o(n_14504) );
na04f04 TIMEBOOST_cell_24467 ( .a(n_9474), .b(g57486_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q), .d(FE_OFN1405_n_8567), .o(n_11251) );
na02f02 TIMEBOOST_cell_49950 ( .a(TIMEBOOST_net_15192), .b(g63378_sb), .o(n_4138) );
na04f04 TIMEBOOST_cell_24469 ( .a(n_9486), .b(g57467_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q), .d(FE_OFN1396_n_8567), .o(n_11265) );
in01s01 TIMEBOOST_cell_73872 ( .a(n_8109), .o(TIMEBOOST_net_23437) );
no02f04 g55633_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243), .o(n_12450) );
na02m02 TIMEBOOST_cell_48564 ( .a(TIMEBOOST_net_14499), .b(FE_OFN569_n_9528), .o(TIMEBOOST_net_11146) );
na04f04 TIMEBOOST_cell_24471 ( .a(n_9487), .b(g57465_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q), .d(FE_OFN1376_n_8567), .o(n_11266) );
na02s02 TIMEBOOST_cell_48260 ( .a(TIMEBOOST_net_14347), .b(g57931_sb), .o(TIMEBOOST_net_10464) );
na02s02 TIMEBOOST_cell_53092 ( .a(TIMEBOOST_net_16763), .b(g58154_sb), .o(TIMEBOOST_net_9498) );
na03f06 TIMEBOOST_cell_64752 ( .a(n_2389), .b(n_4806), .c(n_3018), .o(n_3125) );
na02f02 TIMEBOOST_cell_70459 ( .a(TIMEBOOST_net_22437), .b(FE_OFN1632_n_9531), .o(n_9009) );
na02f02 TIMEBOOST_cell_50476 ( .a(TIMEBOOST_net_15455), .b(g62376_sb), .o(n_6851) );
na02f02 TIMEBOOST_cell_43943 ( .a(pciu_bar0_in_367), .b(n_15598), .o(TIMEBOOST_net_12866) );
no02f04 g55643_u0 ( .a(FE_OCP_RBN2293_FE_OFN1581_n_12306), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_), .o(n_12212) );
na02f02 g55644_u0 ( .a(FE_OCPN1825_n_12030), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q), .o(n_11915) );
na02f04 g55645_u0 ( .a(FE_OFN1564_n_12502), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q), .o(n_11914) );
na02f02 g55646_u0 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q), .o(n_11913) );
na02f04 g55647_u0 ( .a(FE_OFN1556_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q), .o(n_11912) );
na02s01 TIMEBOOST_cell_45435 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q), .o(TIMEBOOST_net_13612) );
na03m06 TIMEBOOST_cell_69898 ( .a(TIMEBOOST_net_17251), .b(FE_OFN1049_n_16657), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q), .o(TIMEBOOST_net_22157) );
na02s02 TIMEBOOST_cell_48566 ( .a(TIMEBOOST_net_14500), .b(FE_OFN1668_n_9477), .o(TIMEBOOST_net_11294) );
na04m02 TIMEBOOST_cell_72613 ( .a(n_3741), .b(FE_OFN653_n_4508), .c(TIMEBOOST_net_10648), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q), .o(TIMEBOOST_net_17387) );
na02m02 TIMEBOOST_cell_63250 ( .a(n_351), .b(n_4909), .o(TIMEBOOST_net_20572) );
na02f02 g55656_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q), .o(n_12206) );
na02f02 g55657_u0 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q), .o(n_11908) );
na02f02 g55658_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q), .o(n_11806) );
in01s01 TIMEBOOST_cell_67788 ( .a(TIMEBOOST_net_21215), .o(TIMEBOOST_net_21214) );
na02s01 TIMEBOOST_cell_43627 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_133), .o(TIMEBOOST_net_12708) );
na02s02 TIMEBOOST_cell_48568 ( .a(TIMEBOOST_net_14501), .b(FE_OFN1668_n_9477), .o(TIMEBOOST_net_11289) );
na02s01 TIMEBOOST_cell_62994 ( .a(configuration_wb_err_addr_551), .b(conf_wb_err_addr_in_960), .o(TIMEBOOST_net_20444) );
na02f02 g55665_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q), .o(n_12203) );
na02f02 g55666_u0 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q), .o(n_11903) );
na02f02 g55667_u0 ( .a(FE_OFN1757_n_12681), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q), .o(n_11805) );
na02m08 TIMEBOOST_cell_68990 ( .a(FE_OFN1644_n_4671), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q), .o(TIMEBOOST_net_21703) );
na02m02 TIMEBOOST_cell_54354 ( .a(TIMEBOOST_net_17394), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_15460) );
na02m02 TIMEBOOST_cell_68833 ( .a(TIMEBOOST_net_21624), .b(n_4482), .o(TIMEBOOST_net_16232) );
na02s01 TIMEBOOST_cell_49275 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q), .b(FE_OFN601_n_9687), .o(TIMEBOOST_net_14855) );
na02s01 TIMEBOOST_cell_37626 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q), .b(pci_target_unit_fifos_pcir_data_in_168), .o(TIMEBOOST_net_10425) );
no02f04 g55675_u0 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__363), .o(n_12449) );
na02s06 TIMEBOOST_cell_68249 ( .a(TIMEBOOST_net_21332), .b(wbu_addr_in_277), .o(TIMEBOOST_net_12393) );
na02s02 TIMEBOOST_cell_48570 ( .a(TIMEBOOST_net_14502), .b(FE_OFN1690_n_9528), .o(TIMEBOOST_net_11114) );
na02f02 TIMEBOOST_cell_70047 ( .a(TIMEBOOST_net_22231), .b(g61790_sb), .o(n_8220) );
na04m04 TIMEBOOST_cell_24487 ( .a(n_9105), .b(g57133_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q), .d(FE_OFN1416_n_8567), .o(n_10470) );
na03f02 TIMEBOOST_cell_73450 ( .a(TIMEBOOST_net_13249), .b(FE_OFN1273_n_4096), .c(g62358_sb), .o(n_6883) );
na02m02 TIMEBOOST_cell_45006 ( .a(TIMEBOOST_net_13397), .b(g58394_db), .o(n_9439) );
no02f04 g55685_u0 ( .a(n_12453), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247), .o(n_12448) );
na02f02 g55686_u0 ( .a(FE_OFN1559_n_12042), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q), .o(n_12196) );
na02f02 g55687_u0 ( .a(FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q), .o(n_12195) );
na04f04 TIMEBOOST_cell_24495 ( .a(n_9408), .b(g57595_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q), .d(FE_OFN1423_n_8567), .o(n_11158) );
na02f02 TIMEBOOST_cell_64097 ( .a(TIMEBOOST_net_21034), .b(FE_OFN1214_n_4151), .o(TIMEBOOST_net_15417) );
na03m02 TIMEBOOST_cell_46703 ( .a(TIMEBOOST_net_12790), .b(g58266_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q), .o(TIMEBOOST_net_9435) );
na02s01 TIMEBOOST_cell_68349 ( .a(TIMEBOOST_net_21382), .b(g65713_db), .o(n_1612) );
no02f04 g55695_u0 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__365), .o(n_12447) );
na04f04 TIMEBOOST_cell_24561 ( .a(n_9207), .b(g57552_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q), .d(FE_OFN1402_n_8567), .o(n_10810) );
na02s02 TIMEBOOST_cell_48572 ( .a(TIMEBOOST_net_14503), .b(FE_OFN1668_n_9477), .o(TIMEBOOST_net_11080) );
no02f01 g55698_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__248), .o(n_11891) );
na02s01 TIMEBOOST_cell_45289 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q), .o(TIMEBOOST_net_13539) );
na03f02 TIMEBOOST_cell_47283 ( .a(FE_OFN1735_n_16317), .b(TIMEBOOST_net_13581), .c(FE_OFN1741_n_11019), .o(n_12768) );
no03f02 TIMEBOOST_cell_66865 ( .a(FE_RN_241_0), .b(TIMEBOOST_net_16479), .c(n_12453), .o(n_12778) );
na02f02 TIMEBOOST_cell_70183 ( .a(TIMEBOOST_net_22299), .b(g54323_sb), .o(TIMEBOOST_net_15953) );
na02f02 TIMEBOOST_cell_49960 ( .a(TIMEBOOST_net_15197), .b(TIMEBOOST_net_329), .o(TIMEBOOST_net_11571) );
na02f02 TIMEBOOST_cell_63147 ( .a(TIMEBOOST_net_20520), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_15699) );
na02m02 TIMEBOOST_cell_54521 ( .a(TIMEBOOST_net_13234), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_17478) );
no02m02 g55707_u0 ( .a(n_11762), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522), .o(n_12186) );
na03f02 TIMEBOOST_cell_70038 ( .a(n_4520), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q), .c(FE_OFN712_n_8140), .o(TIMEBOOST_net_22227) );
na04f04 TIMEBOOST_cell_24497 ( .a(n_9423), .b(g57569_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q), .d(FE_OFN1408_n_8567), .o(n_11182) );
na02s02 TIMEBOOST_cell_48506 ( .a(TIMEBOOST_net_14470), .b(TIMEBOOST_net_12459), .o(TIMEBOOST_net_9402) );
na02m02 TIMEBOOST_cell_68810 ( .a(FE_OFN678_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_21613) );
na02s02 TIMEBOOST_cell_48574 ( .a(TIMEBOOST_net_14504), .b(FE_OFN1687_n_9528), .o(TIMEBOOST_net_11079) );
na02f02 g55714_u0 ( .a(FE_OFN1741_n_11019), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q), .o(n_11887) );
na04f04 TIMEBOOST_cell_23817 ( .a(g62030_da), .b(g62030_db), .c(g52446_sb), .d(g52446_db), .o(n_14846) );
na02f02 TIMEBOOST_cell_70341 ( .a(TIMEBOOST_net_22378), .b(g63589_sb), .o(n_7209) );
no02f02 g55717_u0 ( .a(FE_OCPN1834_n_11884), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484), .o(n_11885) );
ao22f02 g55720_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q), .o(n_11157) );
ao22f02 g55721_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q), .o(n_17016) );
ao22f02 g55722_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q), .o(n_11155) );
ao22f02 g55723_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q), .o(n_11153) );
ao22f02 g55725_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q), .o(n_11793) );
ao22f02 g55726_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q), .o(n_11152) );
ao22f02 g55727_u0 ( .a(FE_OFN1431_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q), .o(n_11149) );
ao22f02 g55728_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q), .o(n_11148) );
ao22f02 g55729_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q), .o(n_11147) );
ao22f02 g55730_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q), .o(n_11146) );
ao22f02 g55731_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q), .o(n_11145) );
ao22f02 g55732_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q), .o(n_11144) );
ao22f02 g55733_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q), .o(n_11143) );
ao22f02 g55734_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q), .o(n_11142) );
ao22f02 g55735_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q), .o(n_11140) );
ao22f02 g55738_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q), .o(n_11136) );
ao22f02 g55739_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q), .o(n_11135) );
ao22f02 g55740_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q), .o(n_11134) );
ao22f02 g55741_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q), .o(n_11132) );
ao22f02 g55742_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q), .o(n_11131) );
ao22f02 g55744_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q), .o(n_11792) );
ao22f02 g55745_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q), .o(n_11130) );
ao22f02 g55746_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q), .o(n_11791) );
ao22f02 g55747_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q), .o(n_16582) );
ao22f02 g55748_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q), .o(n_11129) );
ao22f02 g55749_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q), .o(n_16581) );
ao22f02 g55750_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q), .o(n_11126) );
ao22f02 g55751_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q), .o(n_10788) );
ao22f02 g55752_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q), .o(n_11124) );
ao22f02 g55753_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q), .o(n_11123) );
ao22f02 g55754_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q), .o(n_11122) );
ao22f02 g55755_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q), .o(n_11121) );
ao22f02 g55756_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q), .o(n_11120) );
ao22f02 g55757_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q), .o(n_11119) );
ao22f02 g55759_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q), .o(n_16584) );
ao22f02 g55760_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q), .o(n_11115) );
ao22f02 g55761_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q), .c(FE_OFN1450_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q), .o(n_16583) );
ao22f02 g55763_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q), .c(FE_OFN1450_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q), .o(n_11111) );
ao22f02 g55764_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q), .o(n_11110) );
ao22f02 g55765_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q), .c(n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q), .o(n_11109) );
ao22f02 g55766_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q), .o(n_11108) );
ao22f02 g55767_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q), .o(n_11790) );
ao22f02 g55771_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q), .o(n_11102) );
ao22f02 g55772_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q), .o(n_11101) );
ao22f02 g55773_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q), .o(n_11100) );
ao22f02 g55774_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q), .o(n_11099) );
ao22f02 g55775_u0 ( .a(FE_OFN1431_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q), .o(n_11788) );
ao22f02 g55776_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q), .o(n_11097) );
ao22f02 g55777_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q), .o(n_11096) );
ao22f02 g55778_u0 ( .a(FE_OFN1716_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q), .o(n_11095) );
ao22f02 g55779_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q), .o(n_11094) );
ao22f02 g55781_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q), .o(n_11092) );
ao22f02 g55783_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q), .o(n_10785) );
ao22f02 g55784_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q), .o(n_11090) );
ao22f02 g55785_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q), .o(n_11089) );
ao22f02 g55786_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q), .o(n_11088) );
ao22f02 g55787_u0 ( .a(FE_OCP_RBN2009_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q), .c(FE_OFN1466_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q), .o(n_10784) );
ao22f02 g55788_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q), .o(n_11786) );
ao22f02 g55789_u0 ( .a(FE_OFN1478_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q), .c(FE_OFN2193_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q), .o(n_11087) );
ao22f02 g55790_u0 ( .a(FE_OFN2192_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q), .o(n_11086) );
ao22f02 g55791_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q), .o(n_11784) );
ao22f02 g55792_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q), .o(n_11085) );
ao22f02 g55793_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q), .c(FE_OFN1450_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q), .o(n_11084) );
ao22f02 g55794_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q), .o(n_11083) );
ao22f02 g55795_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q), .o(n_16586) );
ao22f02 g55796_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q), .o(n_11081) );
ao22f02 g55797_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q), .o(n_16585) );
ao22f04 g55798_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q), .o(n_11079) );
ao22f02 g55799_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q), .o(n_11078) );
ao22f02 g55801_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q), .o(n_11076) );
ao22f02 g55802_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q), .o(n_11075) );
ao22f02 g55803_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q), .o(n_11783) );
ao22f02 g55804_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q), .o(n_11782) );
ao22f02 g55806_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q), .o(n_11072) );
ao22f02 g55807_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q), .o(n_11781) );
ao22f02 g55808_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q), .o(n_11071) );
ao22f02 g55809_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q), .o(n_11070) );
ao22f02 g55810_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q), .o(n_11069) );
ao22f02 g55811_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q), .o(n_10782) );
ao22f02 g55812_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q), .o(n_11067) );
ao22f02 g55813_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q), .o(n_11066) );
ao22f02 g55814_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q), .o(n_11065) );
ao22f02 g55815_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q), .o(n_11780) );
ao22f02 g55816_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q), .o(n_11778) );
ao22f02 g55817_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q), .o(n_11064) );
ao22f02 g55818_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q), .o(n_11063) );
ao22f02 g55820_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q), .o(n_11062) );
ao22f02 g55821_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q), .o(n_11061) );
ao22f02 g55822_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q), .o(n_11060) );
ao22f02 g55823_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q), .o(n_11776) );
ao22f02 g55826_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q), .o(n_11057) );
ao22f02 g55827_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q), .o(n_11056) );
ao22f02 g55828_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q), .o(n_11055) );
ao22f02 g55829_u0 ( .a(FE_OFN2208_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q), .c(FE_OFN1455_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q), .o(n_11054) );
ao22f02 g55830_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q), .o(n_11053) );
ao22f02 g55832_u0 ( .a(FE_OCP_RBN2012_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q), .c(FE_OFN1465_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q), .o(n_11050) );
ao22f02 g55833_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q), .o(n_11049) );
ao22f02 g55835_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q), .o(n_11775) );
ao22f02 g55836_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q), .o(n_11047) );
ao22f02 g55837_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q), .o(n_11046) );
ao22f02 g55838_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q), .c(FE_OFN2195_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q), .o(n_11044) );
ao22f02 g55839_u0 ( .a(FE_OCP_RBN2010_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q), .o(n_10781) );
ao22f02 g55840_u0 ( .a(n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q), .c(FE_OFN2194_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q), .o(n_11043) );
ao22f02 g55841_u0 ( .a(FE_OFN1432_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q), .c(FE_OFN1445_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q), .o(n_11042) );
ao22f02 g55842_u0 ( .a(FE_OFN1460_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q), .c(FE_OFN1456_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q), .o(n_11774) );
ao22f02 g55843_u0 ( .a(FE_OFN1431_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q), .c(FE_OFN1444_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q), .o(n_11773) );
ao22f02 g55844_u0 ( .a(FE_OFN1716_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q), .c(FE_OFN1467_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q), .o(n_11041) );
ao22f02 g55845_u0 ( .a(FE_OFN1461_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q), .c(FE_OFN1458_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q), .o(n_11040) );
ao22f02 g55846_u0 ( .a(FE_OFN1477_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q), .c(FE_OFN1449_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q), .o(n_11039) );
ao22f02 g55847_u0 ( .a(FE_OFN1479_n_16637), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q), .c(FE_OFN2196_n_9163), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q), .o(n_11038) );
ao22f02 g55848_u0 ( .a(FE_OFN1433_n_16779), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q), .c(FE_OFN1446_n_11125), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q), .o(n_11037) );
ao22f02 g55849_u0 ( .a(FE_OCP_RBN2011_n_16698), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q), .c(FE_OFN1468_n_10789), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q), .o(n_11036) );
ao22f02 g55850_u0 ( .a(FE_OFN1462_n_11795), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q), .c(FE_OFN1457_n_11138), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q), .o(n_11034) );
in01f02 g55851_u0 ( .a(n_9177), .o(g55851_sb) );
na02m02 TIMEBOOST_cell_54630 ( .a(TIMEBOOST_net_17532), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_15525) );
na03m02 TIMEBOOST_cell_72496 ( .a(n_3761), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q), .c(FE_OFN654_n_4508), .o(TIMEBOOST_net_12569) );
na02f01 TIMEBOOST_cell_26639 ( .a(conf_wb_err_addr_in_954), .b(FE_OFN2069_n_15978), .o(TIMEBOOST_net_7424) );
in01f02 g55852_u0 ( .a(n_9177), .o(g55852_sb) );
na04f04 TIMEBOOST_cell_24663 ( .a(n_9750), .b(g57174_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q), .d(FE_OFN1428_n_8567), .o(n_11582) );
na02m02 TIMEBOOST_cell_53654 ( .a(TIMEBOOST_net_17044), .b(g62546_sb), .o(n_6475) );
na02m04 TIMEBOOST_cell_69020 ( .a(g65059_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q), .o(TIMEBOOST_net_21718) );
in01f02 g55853_u0 ( .a(n_9177), .o(g55853_sb) );
na04f04 TIMEBOOST_cell_24665 ( .a(n_9210), .b(g57505_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q), .d(FE_OFN2184_n_8567), .o(n_10817) );
na02f02 TIMEBOOST_cell_26640 ( .a(TIMEBOOST_net_7424), .b(FE_OFN1145_n_15261), .o(TIMEBOOST_net_597) );
na02f01 TIMEBOOST_cell_27105 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_7657) );
no02f01 g56438_u0 ( .a(FE_OFN778_n_4152), .b(n_4697), .o(n_5744) );
no02f02 g56439_u0 ( .a(n_4800), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8579) );
in01f02 g56450_u0 ( .a(n_9338), .o(n_10780) );
na02f02 g56451_u0 ( .a(n_16313), .b(FE_OCP_RBN2226_g75174_p), .o(n_9338) );
na02f04 g56461_u0 ( .a(n_16334), .b(n_16445), .o(n_10273) );
in01f08 g56466_u0 ( .a(n_12381), .o(n_12357) );
in01f10 g56468_u0 ( .a(n_12099), .o(n_12381) );
in01f08 g56469_u0 ( .a(n_10270), .o(n_12099) );
na02f06 g56470_u0 ( .a(n_16334), .b(n_10258), .o(n_10270) );
in01f06 g56471_u0 ( .a(FE_OCPN1890_n_16553), .o(n_11831) );
in01f06 g56472_u0 ( .a(FE_OCPN1890_n_16553), .o(n_11823) );
in01f04 g56473_u0 ( .a(n_16553), .o(n_12681) );
na02f04 g56485_u0 ( .a(n_16552), .b(n_16445), .o(n_10268) );
in01f04 g56491_u0 ( .a(FE_OCPN1907_n_11767), .o(n_12362) );
in01f06 g56509_u0 ( .a(n_10261), .o(n_12004) );
na02f06 g56510_u0 ( .a(FE_OCP_RBN2282_g74996_p), .b(FE_OCP_RBN2226_g75174_p), .o(n_10261) );
in01f02 g56516_u0 ( .a(FE_OFN1584_n_12306), .o(n_16587) );
in01f04 g56517_u0 ( .a(FE_OFN1579_n_12306), .o(n_11762) );
na02f02 g56522_u0 ( .a(n_16313), .b(n_10258), .o(n_10259) );
in01f02 g56529_u0 ( .a(n_9336), .o(n_12502) );
na02f02 g56530_u0 ( .a(n_16313), .b(n_16364), .o(n_9336) );
in01f02 g56554_u0 ( .a(n_10254), .o(n_12104) );
na02f02 g56555_u0 ( .a(n_16445), .b(FE_OCP_RBN2281_g74996_p), .o(n_10254) );
in01f06 g56556_u0 ( .a(FE_OFN1739_n_11019), .o(n_12293) );
in01f04 g56564_u0 ( .a(n_10252), .o(n_11019) );
na02f04 g56565_u0 ( .a(n_16552), .b(n_16364), .o(n_10252) );
in01f04 g56566_u0 ( .a(n_11884), .o(n_12010) );
in01f03 g56567_u0 ( .a(n_11884), .o(n_11977) );
in01f06 g56568_u0 ( .a(FE_OCPN1834_n_11884), .o(n_12228) );
in01m06 g56572_u0 ( .a(n_11884), .o(n_12001) );
na02f06 g56575_u0 ( .a(FE_OCP_RBN2283_g74996_p), .b(n_10258), .o(n_11884) );
in01f08 g56577_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .o(n_12313) );
in01f10 g56580_u0 ( .a(n_11881), .o(n_12453) );
in01f08 g56582_u0 ( .a(FE_OCP_RBN2286_FE_RN_494_0), .o(n_11881) );
in01f02 g56598_u0 ( .a(n_10244), .o(n_12028) );
na02f02 g56599_u0 ( .a(n_16552), .b(n_10258), .o(n_10244) );
ao22f02 g56600_u0 ( .a(FE_OCPN1879_FE_OFN470_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q), .o(n_16987) );
ao22f02 g56601_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q), .o(n_9335) );
ao22f02 g56602_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q), .o(n_9334) );
ao22f02 g56603_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q), .c(FE_OCPN1872_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q), .o(n_16986) );
in01f02 g56604_u0 ( .a(n_10777), .o(n_11014) );
ao22f02 g56605_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q), .o(n_10777) );
ao22f04 g56606_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q), .c(FE_OFN2206_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q), .o(n_10774) );
ao22f02 g56607_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q), .o(n_10771) );
ao22f02 g56608_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q), .o(n_11013) );
ao22f02 g56609_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q), .o(n_11008) );
ao22f02 g56611_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q), .o(n_9331) );
ao22f02 g56612_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q), .c(n_10232), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q), .o(n_10235) );
in01f02 g56613_u0 ( .a(n_11005), .o(n_11741) );
ao22f02 g56614_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q), .o(n_11005) );
ao22f02 g56615_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q), .o(n_10768) );
ao22f02 g56616_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q), .o(n_10230) );
ao22f02 g56617_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q), .o(n_11002) );
ao22f02 g56619_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q), .o(n_9330) );
ao22f02 g56621_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q), .o(n_9329) );
in01f02 g56622_u0 ( .a(n_10994), .o(n_11740) );
ao22f02 g56623_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q), .o(n_10994) );
ao22f04 g56624_u0 ( .a(FE_OCPN1886_FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q), .o(n_10221) );
ao22f02 g56625_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q), .o(n_10216) );
ao22f02 g56626_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q), .o(n_10991) );
ao22f01 g56627_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q), .c(n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q), .o(n_16843) );
ao22f01 g56629_u0 ( .a(n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q), .o(n_16842) );
ao22f02 g56630_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q), .c(n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q), .o(n_9325) );
in01f02 g56631_u0 ( .a(n_10765), .o(n_10987) );
ao22f02 g56632_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q), .o(n_10765) );
ao22f04 g56633_u0 ( .a(FE_OFN1491_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q), .o(n_10205) );
ao22f02 g56634_u0 ( .a(FE_OFN1728_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q), .c(FE_OCP_RBN1933_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q), .o(n_10202) );
ao22f02 g56635_u0 ( .a(n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q), .o(n_10986) );
ao22f02 g56636_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q), .c(FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q), .o(n_10985) );
ao22f02 g56637_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q), .o(n_9322) );
ao22f02 g56638_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q), .o(n_9321) );
ao22f02 g56639_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q), .c(FE_OCPN2015_n_10195), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q), .o(n_10198) );
in01f02 g56640_u0 ( .a(n_10193), .o(n_10764) );
ao22f02 g56641_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q), .o(n_10193) );
ao22f02 g56642_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q), .o(n_10763) );
ao22f02 g56644_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q), .o(n_10981) );
ao22f02 g56647_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q), .o(n_10183) );
in01f02 g56648_u0 ( .a(n_10755), .o(n_10978) );
ao22f02 g56650_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q), .o(n_9315) );
ao22f02 g56652_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q), .o(n_10754) );
ao22f02 g56653_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q), .o(n_10977) );
ao22f02 g56654_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q), .o(n_9312) );
ao22f02 g56655_u0 ( .a(FE_OCP_RBN1968_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q), .c(n_10185), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q), .o(n_10176) );
in01f02 g56658_u0 ( .a(n_10753), .o(n_10976) );
ao22f02 g56659_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q), .c(n_10693), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q), .o(n_10753) );
ao22f02 g56660_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q), .o(n_10750) );
ao22f04 g56661_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q), .o(n_10747) );
ao22f02 g56662_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q), .o(n_10744) );
ao22f02 g56663_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q), .o(n_9309) );
ao22f02 g56664_u0 ( .a(n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q), .o(n_16849) );
ao22f02 g56665_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q), .c(FE_OFN2143_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q), .o(n_16848) );
ao22f04 g56666_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q), .o(n_10163) );
in01f02 g56667_u0 ( .a(n_10741), .o(n_10975) );
ao22f02 g56669_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q), .c(FE_OFN2206_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q), .o(n_10738) );
ao22f02 g56670_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q), .o(n_10974) );
ao22f04 g56671_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q), .o(n_10160) );
ao22f02 g56672_u0 ( .a(FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q), .o(n_9307) );
ao22f02 g56673_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q), .c(FE_OFN2139_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q), .o(n_10154) );
ao22f02 g56674_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q), .c(FE_OFN1500_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q), .o(n_9306) );
ao22f02 g56675_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q), .o(n_10151) );
in01f02 g56676_u0 ( .a(n_10734), .o(n_10971) );
ao22f02 g56677_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q), .o(n_10734) );
ao22f02 g56678_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q), .o(n_10970) );
ao22f02 g56679_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q), .o(n_10731) );
ao22f04 g56680_u0 ( .a(FE_OCPN1892_FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q), .o(n_10147) );
ao22f02 g56681_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q), .o(n_9305) );
ao22f02 g56683_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q), .c(n_10141), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q), .o(n_10144) );
in01f02 g56685_u0 ( .a(n_10967), .o(n_11739) );
ao22f04 g56686_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q), .o(n_10967) );
ao22f02 g56690_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q), .c(FE_OCP_RBN1934_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q), .o(n_17051) );
ao22f02 g56691_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q), .c(FE_OFN1545_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q), .o(n_9301) );
ao22f02 g56692_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q), .o(n_17050) );
ao22f02 g56693_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q), .o(n_10134) );
in01f02 g56694_u0 ( .a(n_10715), .o(n_10963) );
ao22f01 g56695_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q), .o(n_10715) );
ao22f02 g56696_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q), .o(n_10131) );
ao22f02 g56697_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q), .o(n_10711) );
ao22f02 g56698_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q), .o(n_10708) );
ao22f04 g56699_u0 ( .a(FE_OCPN1879_FE_OFN470_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q), .o(n_10127) );
ao22f02 g56700_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q), .o(n_9299) );
ao22f02 g56701_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q), .o(n_9298) );
ao22f02 g56702_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q), .c(FE_OCPN1872_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q), .o(n_10124) );
in01f02 g56703_u0 ( .a(n_10705), .o(n_10962) );
ao22f02 g56704_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q), .o(n_10705) );
ao22f02 g56706_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q), .c(FE_OFN2206_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q), .o(n_10699) );
ao22f02 g56707_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q), .o(n_10961) );
ao22f02 g56708_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q), .o(n_10956) );
ao22f02 g56710_u0 ( .a(FE_OCP_RBN1968_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q), .c(n_10232), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q), .o(n_10120) );
ao22f02 g56711_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q), .o(n_9296) );
in01f02 g56712_u0 ( .a(n_10696), .o(n_10952) );
ao22f02 g56713_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q), .c(n_10693), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q), .o(n_10696) );
ao22f04 g56715_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q), .o(n_10691) );
ao22f02 g56716_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q), .o(n_10688) );
ao22f02 g56717_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q), .o(n_10116) );
ao22f02 g56718_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q), .o(n_10112) );
ao22f02 g56719_u0 ( .a(n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q), .c(FE_OFN1501_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q), .o(n_9295) );
ao22f02 g56720_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q), .c(FE_OFN1723_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q), .o(n_9294) );
in01f02 g56721_u0 ( .a(n_10947), .o(n_11738) );
ao22f02 g56723_u0 ( .a(FE_OFN1728_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q), .c(FE_OCP_RBN1933_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q), .o(n_10109) );
ao22f02 g56724_u0 ( .a(FE_OFN1539_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q), .c(FE_OFN1521_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q), .o(n_10685) );
ao22f02 g56725_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q), .o(n_10105) );
ao22f02 g56726_u0 ( .a(FE_OFN2148_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q), .o(n_10944) );
ao22f02 g56727_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q), .c(n_10185), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q), .o(n_10102) );
ao22f02 g56728_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q), .o(n_9293) );
ao22f02 g56729_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q), .o(n_9290) );
in01f02 g56730_u0 ( .a(n_10682), .o(n_10943) );
ao22f02 g56731_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q), .o(n_10682) );
ao22f02 g56732_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q), .o(n_10681) );
ao22f02 g56733_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q), .c(n_15568), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q), .o(n_10679) );
ao22f02 g56734_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q), .o(n_10676) );
ao22f02 g56735_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q), .c(FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q), .o(n_10942) );
ao22f02 g56737_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q), .c(n_10141), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q), .o(n_10099) );
ao22f02 g56738_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q), .o(n_9286) );
in01f02 g56739_u0 ( .a(n_10939), .o(n_17042) );
ao22f02 g56740_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q), .o(n_10939) );
ao22f02 g56741_u0 ( .a(FE_OCPN1886_FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q), .o(n_10096) );
ao22f02 g56742_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q), .c(n_15568), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q), .o(n_10675) );
ao22f02 g56743_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q), .o(n_10672) );
ao22f02 g56744_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q), .o(n_9285) );
ao22f02 g56745_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q), .o(n_9284) );
ao22m02 g56746_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q), .c(FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q), .o(n_10093) );
ao22f02 g56747_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q), .c(FE_OCPN2015_n_10195), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q), .o(n_10090) );
in01f02 g56748_u0 ( .a(n_10087), .o(n_10669) );
ao22f02 g56749_u0 ( .a(FE_OCPN1886_FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q), .o(n_10087) );
ao22f02 g56753_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q), .o(n_10084) );
ao22f02 g56754_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q), .o(n_10081) );
ao22f02 g56755_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q), .o(n_9283) );
ao22f02 g56756_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q), .c(FE_OFN1500_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q), .o(n_9280) );
in01f02 g56757_u0 ( .a(n_10662), .o(n_10932) );
ao22f02 g56758_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q), .o(n_10662) );
ao22f02 g56759_u0 ( .a(FE_OFN1728_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q), .c(FE_OCP_RBN1933_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q), .o(n_10661) );
ao22f02 g56761_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q), .o(n_10660) );
ao22f02 g56762_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q), .o(n_9277) );
ao22f02 g56764_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q), .o(n_9276) );
in01f02 g56766_u0 ( .a(n_10927), .o(n_11736) );
ao22f02 g56767_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q), .o(n_10927) );
ao22f02 g56768_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q), .o(n_10075) );
ao22f02 g56769_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q), .o(n_10659) );
ao22f02 g56770_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q), .o(n_10656) );
ao22f02 g56772_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q), .o(n_9274) );
ao22f02 g56773_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q), .c(n_10141), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q), .o(n_17043) );
ao22f02 g56774_u0 ( .a(FE_OFN2149_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q), .c(FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q), .o(n_10069) );
in01f02 g56775_u0 ( .a(n_10653), .o(n_10923) );
ao22f02 g56776_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q), .o(n_10653) );
ao22f02 g56777_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q), .o(n_10650) );
ao22f04 g56778_u0 ( .a(n_10680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q), .o(n_10647) );
ao22f02 g56779_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q), .c(n_15568), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q), .o(n_10644) );
ao22f02 g56780_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q), .o(n_9272) );
ao22f02 g56781_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q), .o(n_10641) );
ao22f02 g56782_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q), .o(n_9271) );
ao22f02 g56783_u0 ( .a(FE_OCP_RBN1968_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q), .c(n_10232), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q), .o(n_10066) );
in01f02 g56784_u0 ( .a(n_10063), .o(n_10638) );
ao22f01 g56785_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q), .o(n_10063) );
ao22f04 g56786_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q), .o(n_10637) );
ao22f04 g56787_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q), .o(n_10060) );
ao22f02 g56788_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q), .c(FE_OCPN1863_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q), .o(n_10634) );
ao22f02 g56789_u0 ( .a(FE_OCP_RBN1969_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q), .c(n_10185), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q), .o(n_10057) );
ao22f02 g56790_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q), .o(n_9270) );
in01f02 g56792_u0 ( .a(n_10051), .o(n_10631) );
ao22f02 g56793_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q), .o(n_10051) );
ao22f02 g56794_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q), .c(FE_OCP_RBN2005_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q), .o(n_9269) );
ao22f04 g56795_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q), .c(FE_OCPN1863_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q), .o(n_10922) );
ao22f02 g56796_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q), .o(n_10630) );
ao22f02 g56797_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q), .c(n_15568), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q), .o(n_10627) );
ao22f02 g56798_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q), .c(FE_OFN1723_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q), .o(n_16835) );
ao22f02 g56799_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q), .o(n_10048) );
in01f02 g56801_u0 ( .a(n_10624), .o(n_10919) );
ao22f02 g56802_u0 ( .a(FE_OFN1539_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q), .c(FE_OFN1521_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q), .o(n_10624) );
ao22f02 g56804_u0 ( .a(FE_OFN1728_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q), .c(FE_OCP_RBN1933_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q), .o(n_10041) );
ao22f02 g56805_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q), .o(n_10038) );
ao22f02 g56806_u0 ( .a(FE_OFN1535_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q), .o(n_10918) );
ao22f02 g56807_u0 ( .a(FE_OFN1453_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q), .c(FE_OFN1529_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q), .o(n_10035) );
ao22f02 g56808_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q), .c(FE_OFN2140_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q), .o(n_10032) );
ao22f02 g56809_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q), .o(n_9262) );
in01f02 g56810_u0 ( .a(n_10622), .o(n_10917) );
ao22f02 g56811_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q), .o(n_10622) );
ao22m02 g56812_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q), .o(n_9261) );
ao22f02 g56813_u0 ( .a(FE_OFN1539_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q), .c(FE_OFN1521_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q), .o(n_10617) );
ao22f02 g56814_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q), .o(n_10029) );
ao22f02 g56815_u0 ( .a(FE_OFN1535_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q), .o(n_10916) );
ao22f02 g56816_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q), .o(n_9260) );
ao22f02 g56818_u0 ( .a(FE_OFN2147_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q), .c(FE_OFN1523_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q), .o(n_10614) );
in01f02 g56820_u0 ( .a(n_10611), .o(n_10913) );
ao22f02 g56821_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q), .o(n_10611) );
ao22f04 g56822_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q), .o(n_11735) );
ao22f02 g56823_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q), .c(FE_OCPN1863_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q), .o(n_10912) );
ao22f04 g56824_u0 ( .a(FE_OCPN1884_n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q), .o(n_10608) );
ao22f02 g56825_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q), .o(n_10020) );
ao22f02 g56826_u0 ( .a(FE_OCPN1879_FE_OFN470_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q), .o(n_10605) );
ao22f02 g56827_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q), .o(n_10017) );
ao22f02 g56828_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q), .c(FE_OCPN1872_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q), .o(n_10602) );
in01f02 g56829_u0 ( .a(n_10909), .o(n_11734) );
ao22f02 g56830_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q), .o(n_10909) );
ao22f02 g56831_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q), .o(n_10908) );
ao22f02 g56833_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q), .o(n_10907) );
ao22f02 g56835_u0 ( .a(FE_OFN2146_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q), .c(FE_OFN1547_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q), .o(n_10014) );
ao22f02 g56837_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q), .o(n_10010) );
in01f02 g56838_u0 ( .a(n_10592), .o(n_10906) );
ao22f02 g56839_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q), .o(n_10592) );
ao22f04 g56840_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q), .o(n_11732) );
ao22f02 g56841_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q), .o(n_10905) );
ao22f02 g56842_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q), .o(n_10904) );
ao22f02 g56843_u0 ( .a(FE_OFN2131_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q), .o(n_16841) );
ao22f02 g56844_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q), .c(FE_OFN2142_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q), .o(n_16840) );
ao22f02 g56845_u0 ( .a(FE_OFN1511_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q), .o(n_10007) );
in01f02 g56846_u0 ( .a(n_10903), .o(n_11731) );
ao22f02 g56849_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q), .o(n_10902) );
ao22f02 g56850_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q), .o(n_10901) );
ao22f02 g56851_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q), .o(n_11730) );
ao22m02 g56853_u0 ( .a(FE_OFN2131_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q), .o(n_10584) );
ao22f02 g56854_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q), .o(n_9997) );
in01f02 g56856_u0 ( .a(n_10898), .o(n_11727) );
ao22f02 g56857_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q), .o(n_10898) );
ao22f02 g56858_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q), .o(n_10579) );
ao22f02 g56860_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q), .o(n_10895) );
ao22f02 g56862_u0 ( .a(n_9991), .b(n_337), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q), .o(n_9993) );
ao22f02 g56863_u0 ( .a(FE_OFN2137_n_15534), .b(n_354), .c(FE_OFN2145_n_16992), .d(n_393), .o(n_16844) );
ao22f02 g56864_u0 ( .a(FE_OFN2131_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q), .c(FE_OFN1528_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q), .o(n_10577) );
in01f02 g56865_u0 ( .a(n_11725), .o(n_11880) );
ao22f02 g56866_u0 ( .a(FE_OFN2216_n_10143), .b(n_251), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q), .o(n_11725) );
ao22f02 g56867_u0 ( .a(FE_OFN2150_n_10595), .b(n_317), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q), .o(n_10891) );
ao22f02 g56868_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q), .o(n_10576) );
ao22f02 g56869_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q), .o(n_10890) );
ao22f02 g56870_u0 ( .a(FE_OCPN1882_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q), .o(n_9992) );
ao22f02 g56871_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q), .o(n_10575) );
ao22f02 g56873_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q), .o(n_10572) );
in01f02 g56874_u0 ( .a(n_10889), .o(n_11724) );
ao22f02 g56875_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q), .o(n_10889) );
ao22f02 g56876_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q), .o(n_11723) );
ao22f02 g56877_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q), .c(FE_OFN1545_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q), .o(n_10569) );
ao22f02 g56878_u0 ( .a(FE_OCPN1892_FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q), .c(FE_OCP_RBN1934_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q), .o(n_10885) );
ao22f02 g56879_u0 ( .a(n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q), .o(n_16851) );
ao22f01 g56880_u0 ( .a(FE_OFN2131_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q), .c(n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q), .o(n_10564) );
ao22f02 g56881_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q), .c(FE_OFN2141_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q), .o(n_16850) );
in01f02 g56883_u0 ( .a(n_10561), .o(n_10882) );
ao22f02 g56884_u0 ( .a(FE_OFN1730_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q), .c(FE_OFN2205_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q), .o(n_10561) );
ao22f02 g56885_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q), .o(n_11720) );
ao22f02 g56886_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q), .c(FE_OFN2207_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q), .o(n_10881) );
ao22f02 g56887_u0 ( .a(FE_OFN1490_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q), .o(n_10880) );
ao22f02 g56890_u0 ( .a(FE_OFN1731_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q), .c(FE_OCP_RBN2006_FE_RN_459_0), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q), .o(n_9976) );
ao22f02 g56891_u0 ( .a(FE_OCP_RBN1968_FE_OFN1532_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q), .c(n_10232), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q), .o(n_10560) );
in01f02 g56892_u0 ( .a(n_10559), .o(n_10876) );
ao22f02 g56893_u0 ( .a(FE_OCPN1881_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q), .c(FE_OFN1498_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q), .o(n_10559) );
ao22f02 g56894_u0 ( .a(FE_OFN2130_n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q), .c(FE_OFN1530_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q), .o(n_10875) );
ao22f04 g56895_u0 ( .a(FE_OCPN1861_FE_OFN468_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q), .c(FE_OCPN1873_FE_OFN474_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q), .o(n_10873) );
ao22f02 g56896_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q), .c(FE_OFN1724_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q), .o(n_10870) );
ao22f02 g56897_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q), .o(n_10556) );
ao22f02 g56898_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q), .c(FE_OFN1723_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q), .o(n_9971) );
ao22f01 g56899_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q), .c(n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q), .o(n_10554) );
ao22f02 g56900_u0 ( .a(n_15566), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q), .c(FE_OFN1501_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q), .o(n_9968) );
in01f02 g56901_u0 ( .a(n_10553), .o(n_10867) );
ao22f02 g56902_u0 ( .a(FE_OCPN1892_FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q), .c(FE_OCP_RBN1934_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q), .o(n_10553) );
ao22f02 g56903_u0 ( .a(FE_OFN1539_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q), .c(FE_OFN1521_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q), .o(n_10866) );
ao22f02 g56904_u0 ( .a(FE_OFN1535_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q), .o(n_11719) );
ao22f02 g56905_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q), .o(n_10865) );
ao22f04 g56906_u0 ( .a(FE_OCPN1882_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q), .c(FE_OFN1500_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q), .o(n_16837) );
ao22f02 g56907_u0 ( .a(FE_OFN1509_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q), .o(n_9962) );
ao22f02 g56908_u0 ( .a(FE_OFN1484_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q), .c(n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q), .o(n_16836) );
ao22f02 g56909_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q), .o(n_10547) );
in01f02 g56910_u0 ( .a(n_10864), .o(n_11718) );
ao22f02 g56911_u0 ( .a(FE_OFN1538_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q), .c(FE_OCPN1915_FE_OFN1522_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q), .o(n_10864) );
ao22f02 g56912_u0 ( .a(FE_OFN1491_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q), .c(n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q), .o(n_10544) );
ao22f04 g56913_u0 ( .a(FE_OCPN1892_FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q), .c(FE_OCP_RBN1934_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q), .o(n_10541) );
ao22f02 g56914_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q), .o(n_11717) );
ao22f02 g56915_u0 ( .a(n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q), .c(FE_OFN1499_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q), .o(n_16839) );
ao22f02 g56916_u0 ( .a(FE_OFN1510_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q), .c(FE_OFN1725_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q), .o(n_9956) );
ao22f02 g56917_u0 ( .a(FE_OFN2137_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q), .c(FE_OFN2142_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q), .o(n_16838) );
in01f02 g56919_u0 ( .a(n_10530), .o(n_10860) );
ao22f02 g56921_u0 ( .a(FE_OFN1493_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q), .c(FE_OFN1546_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q), .o(n_10527) );
ao22f02 g56922_u0 ( .a(FE_OFN2150_n_10595), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q), .c(FE_OFN2206_n_10892), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q), .o(n_10859) );
ao22f02 g56923_u0 ( .a(FE_OFN2216_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q), .c(n_11728), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q), .o(n_11716) );
ao22f02 g56924_u0 ( .a(FE_OFN1727_n_9975), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q), .c(FE_OCP_RBN1932_FE_OFN1515_n_10538), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q), .o(n_9953) );
ao22f02 g56925_u0 ( .a(FE_OFN1489_n_9320), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q), .c(FE_OFN1548_n_10566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q), .o(n_9950) );
ao22f02 g56927_u0 ( .a(FE_OFN1536_n_10143), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q), .c(FE_OCPN2015_n_10195), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q), .o(n_10521) );
in01f02 g56928_u0 ( .a(n_10518), .o(n_10856) );
ao22f02 g56929_u0 ( .a(FE_OCPN1882_n_9991), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q), .c(FE_OFN1502_n_15558), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q), .o(n_10518) );
ao22f04 g56930_u0 ( .a(FE_OFN1485_n_15534), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q), .c(FE_OCPN1888_FE_OFN473_n_16992), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q), .o(n_11715) );
ao22f02 g56931_u0 ( .a(n_10588), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q), .c(FE_OFN1527_n_10853), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q), .o(n_10855) );
ao22f02 g56932_u0 ( .a(FE_OCPN1886_FE_OFN1508_n_15587), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q), .c(FE_OFN1720_n_16891), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q), .o(n_10851) );
in01m20 g56933_u0 ( .a(pci_target_unit_fifos_pcir_flush_in), .o(g56933_sb) );
na02s02 TIMEBOOST_cell_38989 ( .a(TIMEBOOST_net_11106), .b(g58328_db), .o(n_9486) );
in01f10 g56934_u0 ( .a(FE_OFN276_n_9941), .o(g56934_sb) );
na02f04 TIMEBOOST_cell_51581 ( .a(n_13784), .b(FE_OFN1714_n_13650), .o(TIMEBOOST_net_16008) );
na02f01 TIMEBOOST_cell_54198 ( .a(TIMEBOOST_net_17316), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_15169) );
in01f02 g56959_u0 ( .a(n_8934), .o(n_8875) );
no02f06 g56960_u0 ( .a(n_8800), .b(n_2878), .o(n_8934) );
na02m02 TIMEBOOST_cell_18210 ( .a(TIMEBOOST_net_5468), .b(g61829_sb), .o(n_8128) );
in01f08 g56975_u0 ( .a(n_8941), .o(n_10789) );
na02f08 g56976_u0 ( .a(n_9152), .b(n_8939), .o(n_8941) );
na02f10 g56978_u0 ( .a(n_16605), .b(n_9173), .o(n_9256) );
na02f08 g56980_u0 ( .a(n_9173), .b(n_8939), .o(n_8940) );
no02f04 g56985_u0 ( .a(n_9173), .b(n_8924), .o(n_9163) );
in01f06 g56991_u0 ( .a(n_9174), .o(n_11795) );
na02f06 g56992_u0 ( .a(n_9173), .b(n_9171), .o(n_9174) );
in01f06 g56999_u0 ( .a(n_9172), .o(n_11138) );
na02f06 g57000_u0 ( .a(n_9152), .b(n_9171), .o(n_9172) );
in01f06 g57003_u0 ( .a(n_9153), .o(n_11125) );
na02f04 g57009_u0 ( .a(n_9152), .b(n_15516), .o(n_9153) );
na02f04 g57011_u0 ( .a(n_9173), .b(n_15516), .o(n_9170) );
oa12f02 g57019_u0 ( .a(n_8871), .b(pci_target_unit_fifos_pcir_flush_in), .c(n_8876), .o(n_9168) );
oa12f02 g57020_u0 ( .a(n_9160), .b(FE_OFN276_n_9941), .c(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(n_9942) );
oa12f02 g57021_u0 ( .a(n_8950), .b(FE_OFN1394_n_8567), .c(n_9928), .o(n_11710) );
oa12f02 g57022_u0 ( .a(n_8949), .b(FE_OFN2184_n_8567), .c(n_9926), .o(n_11708) );
oa12m02 g57023_u0 ( .a(n_8890), .b(FE_OFN2184_n_8567), .c(n_9924), .o(n_11707) );
oa12f02 g57024_u0 ( .a(n_8889), .b(FE_OFN1403_n_8567), .c(n_9922), .o(n_11706) );
oa12m02 g57025_u0 ( .a(n_8888), .b(FE_OFN1403_n_8567), .c(n_9920), .o(n_11705) );
oa12m02 g57026_u0 ( .a(n_8947), .b(FE_OFN1402_n_8567), .c(n_9918), .o(n_11712) );
oa12m02 g57027_u0 ( .a(n_8946), .b(FE_OFN2184_n_8567), .c(n_9916), .o(n_11703) );
oa12m02 g57028_u0 ( .a(n_8945), .b(FE_OFN1402_n_8567), .c(n_9914), .o(n_11702) );
oa12m02 g57029_u0 ( .a(n_8944), .b(FE_OFN2184_n_8567), .c(n_9912), .o(n_11701) );
no02f04 g57030_u0 ( .a(n_3463), .b(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .o(g57030_p) );
ao12f02 g57030_u1 ( .a(g57030_p), .b(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .c(n_3463), .o(n_4697) );
oa12m02 g57031_u0 ( .a(n_8943), .b(FE_OFN1402_n_8567), .c(n_9910), .o(n_11700) );
oa12m02 g57032_u0 ( .a(n_8887), .b(FE_OFN2184_n_8567), .c(n_9908), .o(n_11699) );
no02f04 g57033_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .b(n_3462), .o(g57033_p) );
ao12f02 g57033_u1 ( .a(g57033_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .c(n_3462), .o(n_4800) );
in01f02 g57034_u0 ( .a(FE_OFN1420_n_8567), .o(g57034_sb) );
na02f02 TIMEBOOST_cell_70193 ( .a(TIMEBOOST_net_22304), .b(g54325_sb), .o(n_12992) );
na02f02 TIMEBOOST_cell_51474 ( .a(TIMEBOOST_net_15954), .b(g52455_da), .o(n_14834) );
na02m01 TIMEBOOST_cell_69822 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q), .o(TIMEBOOST_net_22119) );
in01f02 g57035_u0 ( .a(FE_OFN2179_n_8567), .o(g57035_sb) );
na02f02 TIMEBOOST_cell_70685 ( .a(TIMEBOOST_net_22550), .b(g62827_sb), .o(n_5323) );
na03f02 TIMEBOOST_cell_73355 ( .a(FE_RN_401_0), .b(FE_RN_403_0), .c(FE_RN_402_0), .o(FE_RN_404_0) );
in01f02 g57036_u0 ( .a(FE_OFN1422_n_8567), .o(g57036_sb) );
na02f02 TIMEBOOST_cell_27790 ( .a(TIMEBOOST_net_7999), .b(n_14392), .o(n_14397) );
na03m01 TIMEBOOST_cell_71840 ( .a(TIMEBOOST_net_6772), .b(g54209_sb), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q), .o(TIMEBOOST_net_23128) );
in01f02 g57037_u0 ( .a(FE_OFN1397_n_8567), .o(g57037_sb) );
na02s01 TIMEBOOST_cell_53211 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_796), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q), .o(TIMEBOOST_net_16823) );
na04f02 TIMEBOOST_cell_67580 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q), .b(FE_OFN2104_g64577_p), .c(TIMEBOOST_net_14984), .d(g62808_sb), .o(n_5136) );
na03s02 TIMEBOOST_cell_65528 ( .a(g58275_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q), .c(TIMEBOOST_net_11525), .o(TIMEBOOST_net_9326) );
in01f02 g57038_u0 ( .a(FE_OFN1374_n_8567), .o(g57038_sb) );
na02m10 TIMEBOOST_cell_45647 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q), .o(TIMEBOOST_net_13718) );
na02f01 TIMEBOOST_cell_39561 ( .a(TIMEBOOST_net_11392), .b(g62771_sb), .o(n_5452) );
in01f02 g57039_u0 ( .a(FE_OFN2170_n_8567), .o(g57039_sb) );
na03f02 TIMEBOOST_cell_24997 ( .a(FE_RN_182_0), .b(n_10870), .c(n_12563), .o(n_12825) );
na02s01 TIMEBOOST_cell_42804 ( .a(TIMEBOOST_net_12296), .b(FE_OFN936_n_2292), .o(TIMEBOOST_net_10235) );
na02m02 TIMEBOOST_cell_71892 ( .a(n_3761), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q), .o(TIMEBOOST_net_23154) );
in01f02 g57040_u0 ( .a(FE_OFN2170_n_8567), .o(g57040_sb) );
na03f02 TIMEBOOST_cell_24987 ( .a(n_10763), .b(FE_RN_480_0), .c(n_12587), .o(n_12849) );
na04s02 TIMEBOOST_cell_67373 ( .a(g65215_sb), .b(pci_target_unit_del_sync_bc_in), .c(FE_OFN787_n_2678), .d(pci_target_unit_pcit_if_strd_bc_in), .o(n_2644) );
in01f02 g57041_u0 ( .a(FE_OFN1385_n_8567), .o(g57041_sb) );
na02s01 TIMEBOOST_cell_53213 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_795), .o(TIMEBOOST_net_16824) );
na03f02 TIMEBOOST_cell_66640 ( .a(TIMEBOOST_net_8541), .b(FE_OCPN1847_n_14981), .c(g59118_sb), .o(n_8692) );
in01f02 g57042_u0 ( .a(FE_OFN1423_n_8567), .o(g57042_sb) );
na02s01 TIMEBOOST_cell_68141 ( .a(TIMEBOOST_net_21278), .b(g61989_db), .o(TIMEBOOST_net_14690) );
na02m02 TIMEBOOST_cell_50290 ( .a(TIMEBOOST_net_15362), .b(g62373_sb), .o(n_6857) );
in01f02 g57043_u0 ( .a(FE_OFN1389_n_8567), .o(g57043_sb) );
na04f02 TIMEBOOST_cell_67190 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(g64167_sb), .c(g64167_db), .d(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q), .o(TIMEBOOST_net_15061) );
in01m04 TIMEBOOST_cell_35478 ( .a(TIMEBOOST_net_10108), .o(TIMEBOOST_net_10069) );
na02f04 TIMEBOOST_cell_72215 ( .a(TIMEBOOST_net_23315), .b(TIMEBOOST_net_360), .o(TIMEBOOST_net_11922) );
in01f02 g57044_u0 ( .a(FE_OFN1349_n_8567), .o(g57044_sb) );
na04f04 TIMEBOOST_cell_34997 ( .a(n_9448), .b(g57524_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q), .d(FE_OFN1408_n_8567), .o(n_11217) );
na02s01 TIMEBOOST_cell_47665 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q), .b(g65951_sb), .o(TIMEBOOST_net_14050) );
na02m01 TIMEBOOST_cell_69816 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q), .o(TIMEBOOST_net_22116) );
in01f02 g57045_u0 ( .a(FE_OFN1420_n_8567), .o(g57045_sb) );
na02m10 TIMEBOOST_cell_45649 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q), .o(TIMEBOOST_net_13719) );
in01f02 g57046_u0 ( .a(FE_OFN2177_n_8567), .o(g57046_sb) );
na02s02 TIMEBOOST_cell_37119 ( .a(TIMEBOOST_net_10171), .b(g65268_da), .o(TIMEBOOST_net_8563) );
na02m01 TIMEBOOST_cell_62972 ( .a(configuration_wb_err_addr_560), .b(conf_wb_err_addr_in_969), .o(TIMEBOOST_net_20433) );
in01f02 g57047_u0 ( .a(FE_OFN1390_n_8567), .o(g57047_sb) );
na03f02 TIMEBOOST_cell_65846 ( .a(TIMEBOOST_net_12842), .b(g64244_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q), .o(TIMEBOOST_net_15876) );
in01f02 g57048_u0 ( .a(FE_OFN1407_n_8567), .o(g57048_sb) );
na02s03 TIMEBOOST_cell_53215 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_770), .o(TIMEBOOST_net_16825) );
in01m04 TIMEBOOST_cell_35480 ( .a(TIMEBOOST_net_10110), .o(TIMEBOOST_net_10071) );
in01f02 g57049_u0 ( .a(FE_OFN2190_n_8567), .o(g57049_sb) );
na02m01 TIMEBOOST_cell_25294 ( .a(TIMEBOOST_net_6751), .b(n_574), .o(TIMEBOOST_net_5360) );
na02s01 TIMEBOOST_cell_48831 ( .a(FE_OFN211_n_9858), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q), .o(TIMEBOOST_net_14633) );
in01f02 g57050_u0 ( .a(FE_OFN2190_n_8567), .o(g57050_sb) );
na02s01 TIMEBOOST_cell_48013 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q), .b(FE_OFN1649_n_9428), .o(TIMEBOOST_net_14224) );
na02s02 TIMEBOOST_cell_51311 ( .a(g58231_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q), .o(TIMEBOOST_net_15873) );
in01f02 g57051_u0 ( .a(FE_OFN1397_n_8567), .o(g57051_sb) );
na03m02 TIMEBOOST_cell_66580 ( .a(n_4594), .b(g61959_sb), .c(g61959_db), .o(n_6953) );
na03m02 TIMEBOOST_cell_72832 ( .a(g64872_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q), .c(TIMEBOOST_net_17233), .o(TIMEBOOST_net_17439) );
in01f02 g57052_u0 ( .a(FE_OFN1383_n_8567), .o(g57052_sb) );
in01s01 TIMEBOOST_cell_73925 ( .a(TIMEBOOST_net_23489), .o(TIMEBOOST_net_23490) );
na02f01 TIMEBOOST_cell_53040 ( .a(TIMEBOOST_net_16737), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_15293) );
in01f02 g57053_u0 ( .a(FE_OFN1385_n_8567), .o(g57053_sb) );
in01s01 TIMEBOOST_cell_73960 ( .a(wbm_dat_i_2_), .o(TIMEBOOST_net_23525) );
na02f08 TIMEBOOST_cell_37123 ( .a(TIMEBOOST_net_10173), .b(n_2753), .o(TIMEBOOST_net_217) );
no03f04 TIMEBOOST_cell_67094 ( .a(FE_RN_818_0), .b(FE_RN_817_0), .c(FE_RN_816_0), .o(n_14438) );
in01f02 g57055_u0 ( .a(FE_OFN2179_n_8567), .o(g57055_sb) );
na02s01 TIMEBOOST_cell_47513 ( .a(parchk_pci_ad_reg_in_1205), .b(g67083_db), .o(TIMEBOOST_net_13974) );
na03f02 TIMEBOOST_cell_51575 ( .a(n_17050), .b(n_17051), .c(n_9301), .o(TIMEBOOST_net_16005) );
in01f02 g57056_u0 ( .a(FE_OFN1368_n_8567), .o(g57056_sb) );
na02m02 TIMEBOOST_cell_48832 ( .a(TIMEBOOST_net_14633), .b(FE_OFN580_n_9531), .o(TIMEBOOST_net_12805) );
in01s01 TIMEBOOST_cell_45948 ( .a(TIMEBOOST_net_13908), .o(TIMEBOOST_net_13909) );
in01f02 g57057_u0 ( .a(FE_OFN1392_n_8567), .o(g57057_sb) );
na03f02 TIMEBOOST_cell_66444 ( .a(TIMEBOOST_net_16772), .b(FE_OFN1311_n_6624), .c(g62983_sb), .o(n_5916) );
na02s01 TIMEBOOST_cell_28983 ( .a(pci_target_unit_fifos_outGreyCount_reg_1__Q), .b(n_996), .o(TIMEBOOST_net_8596) );
in01f02 g57058_u0 ( .a(FE_OFN2174_n_8567), .o(g57058_sb) );
na02f02 TIMEBOOST_cell_51002 ( .a(TIMEBOOST_net_15718), .b(g63185_sb), .o(n_5782) );
na02m02 TIMEBOOST_cell_53821 ( .a(n_4222), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q), .o(TIMEBOOST_net_17128) );
na03m06 TIMEBOOST_cell_68728 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(FE_OFN917_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q), .o(TIMEBOOST_net_21572) );
in01f02 g57059_u0 ( .a(FE_OFN2178_n_8567), .o(g57059_sb) );
na02s02 TIMEBOOST_cell_63067 ( .a(TIMEBOOST_net_20480), .b(FE_OFN1632_n_9531), .o(TIMEBOOST_net_10772) );
na02f01 TIMEBOOST_cell_53167 ( .a(n_13175), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q), .o(TIMEBOOST_net_16801) );
in01f02 g57060_u0 ( .a(FE_OFN2174_n_8567), .o(g57060_sb) );
na02f01 TIMEBOOST_cell_31738 ( .a(TIMEBOOST_net_9973), .b(FE_OFN881_g64577_p), .o(TIMEBOOST_net_7342) );
na02m01 TIMEBOOST_cell_68974 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q), .b(FE_OFN618_n_4490), .o(TIMEBOOST_net_21695) );
na02s01 TIMEBOOST_cell_52643 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q), .o(TIMEBOOST_net_16539) );
in01f02 g57061_u0 ( .a(FE_OFN1377_n_8567), .o(g57061_sb) );
na02m10 TIMEBOOST_cell_45655 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q), .o(TIMEBOOST_net_13722) );
na02m02 TIMEBOOST_cell_53647 ( .a(TIMEBOOST_net_13229), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_17041) );
in01f02 g57062_u0 ( .a(FE_OFN1399_n_8567), .o(g57062_sb) );
na03f02 TIMEBOOST_cell_70588 ( .a(n_4729), .b(n_255), .c(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_22502) );
na02s01 TIMEBOOST_cell_47774 ( .a(TIMEBOOST_net_14104), .b(FE_OFN941_n_2047), .o(TIMEBOOST_net_12392) );
in01f01 g57063_u0 ( .a(FE_OFN1394_n_8567), .o(g57063_sb) );
na03m06 TIMEBOOST_cell_69080 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN908_n_4734), .c(TIMEBOOST_net_16604), .o(TIMEBOOST_net_21748) );
in01f02 g57064_u0 ( .a(FE_OFN2167_n_8567), .o(g57064_sb) );
na03m02 TIMEBOOST_cell_72804 ( .a(n_4476), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q), .c(TIMEBOOST_net_12551), .o(TIMEBOOST_net_20617) );
na02s01 g54207_u1 ( .a(g54207_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_395), .o(g54207_da) );
in01f02 g57065_u0 ( .a(FE_OFN1412_n_8567), .o(g57065_sb) );
na02s03 TIMEBOOST_cell_53217 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_793), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q), .o(TIMEBOOST_net_16826) );
na04f04 TIMEBOOST_cell_67920 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q), .b(FE_OFN707_n_8119), .c(g61952_sb), .d(n_1707), .o(n_7921) );
in01f02 g57066_u0 ( .a(FE_OFN1397_n_8567), .o(g57066_sb) );
na02s01 TIMEBOOST_cell_49512 ( .a(TIMEBOOST_net_14973), .b(g58019_sb), .o(TIMEBOOST_net_9502) );
na02f02 TIMEBOOST_cell_4209 ( .a(TIMEBOOST_net_664), .b(n_14387), .o(n_14388) );
in01f02 g57067_u0 ( .a(FE_OFN2173_n_8567), .o(g57067_sb) );
na02s01 TIMEBOOST_cell_44451 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q), .b(g58291_sb), .o(TIMEBOOST_net_13120) );
na02f02 TIMEBOOST_cell_70533 ( .a(TIMEBOOST_net_22474), .b(g63392_sb), .o(n_4134) );
na02m20 TIMEBOOST_cell_62924 ( .a(pci_target_unit_pcit_if_strd_addr_in_703), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67), .o(TIMEBOOST_net_20409) );
in01f02 g57068_u0 ( .a(FE_OFN1423_n_8567), .o(g57068_sb) );
na02s01 TIMEBOOST_cell_45657 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q), .o(TIMEBOOST_net_13723) );
na02f02 TIMEBOOST_cell_4211 ( .a(TIMEBOOST_net_665), .b(n_14392), .o(n_14393) );
in01f02 g57069_u0 ( .a(FE_OFN1421_n_8567), .o(g57069_sb) );
na02s01 TIMEBOOST_cell_48151 ( .a(g58181_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_14293) );
na02f02 TIMEBOOST_cell_4213 ( .a(TIMEBOOST_net_666), .b(n_14390), .o(n_14391) );
na02f01 TIMEBOOST_cell_40080 ( .a(FE_OFN1179_n_3476), .b(configuration_pci_err_addr_478), .o(TIMEBOOST_net_11652) );
in01f02 g57070_u0 ( .a(FE_OFN1404_n_8567), .o(g57070_sb) );
na03s02 TIMEBOOST_cell_67859 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q), .b(FE_OFN217_n_9889), .c(FE_OFN588_n_9692), .o(TIMEBOOST_net_12466) );
in01f02 g57071_u0 ( .a(FE_OFN1425_n_8567), .o(g57071_sb) );
na03f02 TIMEBOOST_cell_73595 ( .a(TIMEBOOST_net_17435), .b(FE_OFN1285_n_4097), .c(g62391_sb), .o(n_6816) );
na03f04 TIMEBOOST_cell_66437 ( .a(TIMEBOOST_net_17120), .b(FE_OFN1311_n_6624), .c(g62660_sb), .o(n_6223) );
in01f02 g57072_u0 ( .a(FE_OFN1370_n_8567), .o(g57072_sb) );
na03f02 TIMEBOOST_cell_65165 ( .a(TIMEBOOST_net_16252), .b(g64181_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q), .o(TIMEBOOST_net_15060) );
in01f02 g57073_u0 ( .a(FE_OFN1415_n_8567), .o(g57073_sb) );
na02s01 TIMEBOOST_cell_53219 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_794), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q), .o(TIMEBOOST_net_16827) );
na02f02 TIMEBOOST_cell_4221 ( .a(TIMEBOOST_net_670), .b(n_8529), .o(n_8530) );
na02f01 g64648_u0 ( .a(n_2799), .b(n_12179), .o(n_3269) );
in01f02 g57074_u0 ( .a(FE_OFN2169_n_8567), .o(g57074_sb) );
na04m02 TIMEBOOST_cell_72817 ( .a(g64881_sb), .b(n_3777), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q), .d(TIMEBOOST_net_12737), .o(TIMEBOOST_net_17449) );
in01f02 g57075_u0 ( .a(FE_OFN1405_n_8567), .o(g57075_sb) );
na02s01 TIMEBOOST_cell_53223 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_767), .o(TIMEBOOST_net_16829) );
na03m02 TIMEBOOST_cell_72853 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q), .b(g65367_sb), .c(TIMEBOOST_net_22082), .o(TIMEBOOST_net_17443) );
in01f02 g57076_u0 ( .a(FE_OFN2182_n_8567), .o(g57076_sb) );
na02m01 TIMEBOOST_cell_70342 ( .a(TIMEBOOST_net_16954), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_22379) );
na03f02 TIMEBOOST_cell_73566 ( .a(TIMEBOOST_net_17495), .b(FE_OFN1232_n_6391), .c(g62455_sb), .o(n_6686) );
in01f02 g57077_u0 ( .a(FE_OFN1408_n_8567), .o(g57077_sb) );
na02f01 TIMEBOOST_cell_26085 ( .a(pci_target_unit_pcit_if_strd_addr_in_703), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7147) );
na03m04 TIMEBOOST_cell_73087 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q), .b(g65355_sb), .c(TIMEBOOST_net_22276), .o(TIMEBOOST_net_17500) );
in01f02 g57078_u0 ( .a(FE_OFN1389_n_8567), .o(g57078_sb) );
na03f02 TIMEBOOST_cell_73596 ( .a(TIMEBOOST_net_17466), .b(FE_OFN1285_n_4097), .c(g62385_sb), .o(n_6830) );
na02m02 TIMEBOOST_cell_69403 ( .a(TIMEBOOST_net_21909), .b(g64988_sb), .o(TIMEBOOST_net_12690) );
in01f02 g57079_u0 ( .a(FE_OFN1349_n_8567), .o(g57079_sb) );
na04f04 TIMEBOOST_cell_34999 ( .a(n_9890), .b(g57041_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q), .d(FE_OFN1376_n_8567), .o(n_11693) );
na03m02 TIMEBOOST_cell_67166 ( .a(n_3755), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q), .c(FE_OFN1663_n_4490), .o(TIMEBOOST_net_10576) );
na02m01 TIMEBOOST_cell_53998 ( .a(TIMEBOOST_net_17216), .b(FE_OFN687_n_4417), .o(TIMEBOOST_net_14314) );
in01f02 g57080_u0 ( .a(FE_OFN1421_n_8567), .o(g57080_sb) );
na03f02 TIMEBOOST_cell_67953 ( .a(TIMEBOOST_net_13104), .b(FE_OFN1132_g64577_p), .c(g62765_sb), .o(n_5465) );
na03m02 TIMEBOOST_cell_73150 ( .a(TIMEBOOST_net_14702), .b(g64265_sb), .c(g63052_sb), .o(TIMEBOOST_net_22372) );
in01f02 g57081_u0 ( .a(FE_OFN1392_n_8567), .o(g57081_sb) );
na02m08 TIMEBOOST_cell_53037 ( .a(wbm_adr_o_15_), .b(configuration_pci_err_addr_485), .o(TIMEBOOST_net_16736) );
na02f08 g75178_u1 ( .a(FE_OCP_RBN2232_n_16273), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .o(g75178_da) );
in01f02 g57082_u0 ( .a(FE_OFN1406_n_8567), .o(g57082_sb) );
na02f01 TIMEBOOST_cell_70578 ( .a(TIMEBOOST_net_13044), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_22497) );
na02f01 TIMEBOOST_cell_37450 ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_10337) );
in01f02 g57083_u0 ( .a(FE_OFN1406_n_8567), .o(g57083_sb) );
na02f01 TIMEBOOST_cell_37451 ( .a(TIMEBOOST_net_10337), .b(g53940_sb), .o(TIMEBOOST_net_587) );
in01f02 g57084_u0 ( .a(FE_OFN1424_n_8567), .o(g57084_sb) );
na04f06 TIMEBOOST_cell_64282 ( .a(n_16284), .b(n_16285), .c(conf_w_addr_in_938), .d(n_16696), .o(n_16286) );
na03f02 TIMEBOOST_cell_33379 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_791), .b(g54315_sb), .c(g54315_db), .o(n_13012) );
in01f02 g57085_u0 ( .a(FE_OFN1422_n_8567), .o(g57085_sb) );
na03f02 TIMEBOOST_cell_66958 ( .a(TIMEBOOST_net_16509), .b(n_11831), .c(n_12357), .o(n_12645) );
na03m02 TIMEBOOST_cell_64604 ( .a(n_3636), .b(FE_OFN622_n_4409), .c(n_3783), .o(TIMEBOOST_net_12426) );
in01f02 g57086_u0 ( .a(FE_OFN1370_n_8567), .o(g57086_sb) );
na02f01 TIMEBOOST_cell_26095 ( .a(pci_target_unit_pcit_if_strd_addr_in_711), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7152) );
na02f01 TIMEBOOST_cell_51852 ( .a(TIMEBOOST_net_16143), .b(n_261), .o(n_9834) );
in01f02 g57087_u0 ( .a(FE_OFN1414_n_8567), .o(g57087_sb) );
na02m06 TIMEBOOST_cell_68988 ( .a(FE_OFN615_n_4501), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q), .o(TIMEBOOST_net_21702) );
na03s01 TIMEBOOST_cell_41723 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q), .b(g58430_sb), .c(g58430_db), .o(n_8996) );
na02m02 TIMEBOOST_cell_4242 ( .a(pci_target_unit_fifos_pcir_flush_in), .b(g57787_da), .o(TIMEBOOST_net_681) );
in01f02 g57088_u0 ( .a(FE_OFN1414_n_8567), .o(g57088_sb) );
na02f01 TIMEBOOST_cell_26111 ( .a(pci_target_unit_pcit_if_strd_addr_in_713), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_7160) );
in01f02 g57089_u0 ( .a(FE_OFN1419_n_8567), .o(g57089_sb) );
na02f01 TIMEBOOST_cell_26109 ( .a(pci_target_unit_pcit_if_strd_addr_in_700), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7159) );
na03m02 TIMEBOOST_cell_64603 ( .a(FE_OFN624_n_4409), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q), .c(n_3770), .o(TIMEBOOST_net_10637) );
na02m02 TIMEBOOST_cell_4246 ( .a(pci_target_unit_fifos_pcir_flush_in), .b(g57788_da), .o(TIMEBOOST_net_683) );
in01f02 g57090_u0 ( .a(FE_OFN1415_n_8567), .o(g57090_sb) );
na02f01 TIMEBOOST_cell_26097 ( .a(pci_target_unit_pcit_if_strd_addr_in_714), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_7153) );
in01f02 g57091_u0 ( .a(FE_OFN1368_n_8567), .o(g57091_sb) );
na02f02 TIMEBOOST_cell_40845 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_12034), .o(TIMEBOOST_net_476) );
in01f02 g57092_u0 ( .a(FE_OFN1401_n_8567), .o(g57092_sb) );
na02f02 TIMEBOOST_cell_4251 ( .a(TIMEBOOST_net_685), .b(n_15517), .o(n_8853) );
na02m02 TIMEBOOST_cell_68298 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q), .b(n_4669), .o(TIMEBOOST_net_21357) );
in01f02 g57093_u0 ( .a(FE_OFN2169_n_8567), .o(g57093_sb) );
na02s01 TIMEBOOST_cell_53104 ( .a(TIMEBOOST_net_16769), .b(g58121_db), .o(n_9671) );
na02f01 TIMEBOOST_cell_44382 ( .a(TIMEBOOST_net_13085), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_11415) );
in01f02 g57094_u0 ( .a(FE_OFN2184_n_8567), .o(g57094_sb) );
na02s01 TIMEBOOST_cell_71370 ( .a(FE_OFN221_n_9846), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q), .o(TIMEBOOST_net_22893) );
na02s01 TIMEBOOST_cell_31093 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_9651) );
in01f02 g57095_u0 ( .a(FE_OFN1417_n_8567), .o(g57095_sb) );
na03f02 TIMEBOOST_cell_34890 ( .a(TIMEBOOST_net_9378), .b(FE_OFN1404_n_8567), .c(g57309_sb), .o(n_11441) );
in01f02 g57096_u0 ( .a(FE_OFN1377_n_8567), .o(g57096_sb) );
na02f02 TIMEBOOST_cell_40841 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_12032), .o(n_12752) );
na03f02 TIMEBOOST_cell_66505 ( .a(TIMEBOOST_net_16783), .b(FE_OFN1317_n_6624), .c(g63161_sb), .o(n_5814) );
no02f06 TIMEBOOST_cell_4256 ( .a(n_1513), .b(FE_RN_281_0), .o(TIMEBOOST_net_688) );
in01f02 g57097_u0 ( .a(FE_OFN1403_n_8567), .o(g57097_sb) );
na03f02 TIMEBOOST_cell_65895 ( .a(n_3872), .b(g63086_sb), .c(g63086_db), .o(n_5082) );
na03f02 TIMEBOOST_cell_34851 ( .a(TIMEBOOST_net_9490), .b(FE_OFN1420_n_8567), .c(g57034_sb), .o(n_11698) );
na03m02 TIMEBOOST_cell_72650 ( .a(TIMEBOOST_net_21492), .b(g64841_sb), .c(TIMEBOOST_net_21672), .o(TIMEBOOST_net_20538) );
in01f02 g57098_u0 ( .a(FE_OFN1405_n_8567), .o(g57098_sb) );
na02s02 TIMEBOOST_cell_4259 ( .a(TIMEBOOST_net_689), .b(n_16332), .o(g58582_p) );
in01f02 g57099_u0 ( .a(FE_OFN1380_n_8567), .o(g57099_sb) );
na02s01 TIMEBOOST_cell_70461 ( .a(TIMEBOOST_net_22438), .b(FE_OFN209_n_9126), .o(TIMEBOOST_net_10566) );
na02f10 TIMEBOOST_cell_38730 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_792), .o(TIMEBOOST_net_10977) );
na03f03 TIMEBOOST_cell_54733 ( .a(FE_RN_641_0), .b(FE_RN_666_0), .c(FE_RN_631_0), .o(TIMEBOOST_net_17584) );
in01f02 g57100_u0 ( .a(FE_OFN1400_n_8567), .o(g57100_sb) );
na02f02 TIMEBOOST_cell_70687 ( .a(TIMEBOOST_net_22551), .b(g63028_sb), .o(n_5190) );
na02f02 TIMEBOOST_cell_4263 ( .a(TIMEBOOST_net_691), .b(n_8897), .o(n_9932) );
na02s01 TIMEBOOST_cell_4264 ( .a(g59126_db), .b(g59126_sb), .o(TIMEBOOST_net_692) );
in01f02 g57101_u0 ( .a(FE_OFN1382_n_8567), .o(g57101_sb) );
na02f02 TIMEBOOST_cell_4265 ( .a(TIMEBOOST_net_692), .b(n_8582), .o(n_8583) );
in01f02 g57102_u0 ( .a(FE_OFN1420_n_8567), .o(g57102_sb) );
na02f02 TIMEBOOST_cell_4267 ( .a(n_10106), .b(TIMEBOOST_net_693), .o(n_11858) );
na03f02 TIMEBOOST_cell_34837 ( .a(TIMEBOOST_net_9421), .b(FE_OFN1407_n_8567), .c(g57361_sb), .o(n_11385) );
in01f02 g57103_u0 ( .a(FE_OFN1425_n_8567), .o(g57103_sb) );
na03f02 TIMEBOOST_cell_34892 ( .a(TIMEBOOST_net_9433), .b(FE_OFN1391_n_8567), .c(g57560_sb), .o(n_10298) );
na02f08 TIMEBOOST_cell_4269 ( .a(TIMEBOOST_net_694), .b(n_16331), .o(n_8820) );
na02f01 TIMEBOOST_cell_4270 ( .a(FE_OFN1023_n_11877), .b(g52479_da), .o(TIMEBOOST_net_695) );
in01f02 g57104_u0 ( .a(FE_OFN1411_n_8567), .o(g57104_sb) );
na03f02 TIMEBOOST_cell_72945 ( .a(pci_target_unit_del_sync_addr_in_224), .b(g65226_sb), .c(TIMEBOOST_net_7154), .o(n_2661) );
na02s01 TIMEBOOST_cell_48577 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q), .o(TIMEBOOST_net_14506) );
in01f02 g57105_u0 ( .a(FE_OFN1404_n_8567), .o(g57105_sb) );
na02s01 TIMEBOOST_cell_62422 ( .a(n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_20158) );
na03f40 TIMEBOOST_cell_72376 ( .a(conf_wb_err_bc_in_846), .b(g67048_sb), .c(TIMEBOOST_net_13990), .o(n_1211) );
na03m02 TIMEBOOST_cell_72773 ( .a(n_4493), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q), .c(TIMEBOOST_net_12756), .o(TIMEBOOST_net_17063) );
in01f02 g57106_u0 ( .a(FE_OFN1423_n_8567), .o(g57106_sb) );
na02f01 TIMEBOOST_cell_26091 ( .a(pci_target_unit_pcit_if_strd_addr_in_701), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7150) );
na03f20 TIMEBOOST_cell_72382 ( .a(pci_cbe_i_0_), .b(g67044_sb), .c(parchk_pci_cbe_en_in), .o(TIMEBOOST_net_23126) );
na03f02 TIMEBOOST_cell_65396 ( .a(wbs_we_i), .b(g63588_sb), .c(g63588_db), .o(n_4100) );
in01f02 g57107_u0 ( .a(FE_OFN1381_n_8567), .o(g57107_sb) );
na03f02 TIMEBOOST_cell_34894 ( .a(TIMEBOOST_net_9374), .b(FE_OFN1370_n_8567), .c(g57447_sb), .o(n_10349) );
na04f01 TIMEBOOST_cell_72392 ( .a(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .b(wishbone_slave_unit_delayed_write_data_comp_wdata_out_80), .c(g54205_sb), .d(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q), .o(TIMEBOOST_net_21275) );
na02f02 TIMEBOOST_cell_54476 ( .a(TIMEBOOST_net_17455), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_15428) );
in01f02 g57108_u0 ( .a(FE_OFN1415_n_8567), .o(g57108_sb) );
na02s01 TIMEBOOST_cell_53491 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q), .o(TIMEBOOST_net_16963) );
na03m04 TIMEBOOST_cell_72388 ( .a(n_947), .b(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .c(wishbone_slave_unit_del_sync_comp_cycle_count_5_), .o(TIMEBOOST_net_31) );
na02f02 TIMEBOOST_cell_70371 ( .a(TIMEBOOST_net_22393), .b(g63594_sb), .o(n_7205) );
in01f02 g57109_u0 ( .a(FE_OFN2167_n_8567), .o(g57109_sb) );
na03f02 TIMEBOOST_cell_73597 ( .a(TIMEBOOST_net_13242), .b(FE_OFN1243_n_4092), .c(g62508_sb), .o(n_6563) );
na02s01 TIMEBOOST_cell_31095 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_9652) );
na03m01 TIMEBOOST_cell_72424 ( .a(TIMEBOOST_net_14007), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q), .c(wbu_addr_in_256), .o(n_9789) );
in01f02 g57110_u0 ( .a(FE_OFN1405_n_8567), .o(g57110_sb) );
na04f20 TIMEBOOST_cell_72386 ( .a(conf_wb_err_addr_in_971), .b(conf_wb_err_addr_in_970), .c(n_1442), .d(n_1441), .o(n_1443) );
in01f02 g57111_u0 ( .a(FE_OFN2182_n_8567), .o(g57111_sb) );
na03f02 TIMEBOOST_cell_73811 ( .a(TIMEBOOST_net_16546), .b(FE_OFN1773_n_13800), .c(FE_OFN1769_n_14054), .o(g53254_p) );
na02m02 TIMEBOOST_cell_50394 ( .a(TIMEBOOST_net_15414), .b(g62989_sb), .o(n_5904) );
in01f02 g57112_u0 ( .a(FE_OFN1409_n_8567), .o(g57112_sb) );
na03f02 TIMEBOOST_cell_72780 ( .a(n_4470), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q), .c(TIMEBOOST_net_10591), .o(TIMEBOOST_net_17396) );
na03s02 TIMEBOOST_cell_64919 ( .a(FE_OFN540_n_9690), .b(g58232_sb), .c(TIMEBOOST_net_12781), .o(n_9546) );
in01f02 g57113_u0 ( .a(FE_OFN1388_n_8567), .o(g57113_sb) );
na03f20 TIMEBOOST_cell_72380 ( .a(pci_cbe_i_3_), .b(g67046_sb), .c(parchk_pci_cbe_en_in), .o(TIMEBOOST_net_23124) );
na02f02 TIMEBOOST_cell_54692 ( .a(TIMEBOOST_net_17563), .b(FE_OFN1257_n_4143), .o(TIMEBOOST_net_15398) );
in01f02 g57114_u0 ( .a(FE_OFN1421_n_8567), .o(g57114_sb) );
na03f01 TIMEBOOST_cell_68080 ( .a(pci_ad_i_15_), .b(n_574), .c(parchk_pci_ad_reg_in_1219), .o(TIMEBOOST_net_21248) );
no04f40 TIMEBOOST_cell_72372 ( .a(n_544), .b(n_715), .c(conf_wb_err_bc_in_848), .d(TIMEBOOST_net_12242), .o(TIMEBOOST_net_10180) );
na03f02 TIMEBOOST_cell_65397 ( .a(TIMEBOOST_net_16621), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .c(g52628_sb), .o(n_14678) );
in01f02 g57115_u0 ( .a(FE_OFN1345_n_8567), .o(g57115_sb) );
na02s01 TIMEBOOST_cell_43659 ( .a(pci_target_unit_del_sync_addr_in_233), .b(n_2509), .o(TIMEBOOST_net_12724) );
in01f02 g57116_u0 ( .a(FE_OFN1406_n_8567), .o(g57116_sb) );
na03f02 TIMEBOOST_cell_66400 ( .a(TIMEBOOST_net_21024), .b(n_8590), .c(g59089_sb), .o(n_8589) );
na03s01 TIMEBOOST_cell_72378 ( .a(pci_target_unit_fifos_pcir_whole_waddr_94), .b(pci_target_unit_fifos_pcir_flush_in), .c(g57780_sb), .o(TIMEBOOST_net_685) );
in01f02 g57117_u0 ( .a(FE_OFN1389_n_8567), .o(g57117_sb) );
in01s01 TIMEBOOST_cell_73929 ( .a(TIMEBOOST_net_23493), .o(TIMEBOOST_net_23494) );
na04f04 TIMEBOOST_cell_67596 ( .a(TIMEBOOST_net_13849), .b(g62104_sb), .c(FE_OFN1163_n_5615), .d(configuration_wb_err_data_573), .o(n_5597) );
in01f02 g57118_u0 ( .a(FE_OFN1368_n_8567), .o(g57118_sb) );
na03m10 TIMEBOOST_cell_72374 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q), .b(TIMEBOOST_net_12733), .c(FE_OFN1034_n_4732), .o(TIMEBOOST_net_23279) );
in01f02 g57119_u0 ( .a(FE_OFN2191_n_8567), .o(g57119_sb) );
na02f02 TIMEBOOST_cell_50880 ( .a(TIMEBOOST_net_15657), .b(g62474_sb), .o(n_6641) );
na03f02 TIMEBOOST_cell_66950 ( .a(FE_OFN1572_n_11027), .b(TIMEBOOST_net_16504), .c(FE_OFN1752_n_12086), .o(n_12706) );
in01f02 g57120_u0 ( .a(FE_OFN1424_n_8567), .o(g57120_sb) );
na02m04 TIMEBOOST_cell_69407 ( .a(TIMEBOOST_net_21911), .b(FE_OFN1058_n_4727), .o(TIMEBOOST_net_16958) );
na03s02 TIMEBOOST_cell_72370 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q), .c(FE_OFN953_n_2055), .o(TIMEBOOST_net_16193) );
in01f02 g57121_u0 ( .a(FE_OFN1380_n_8567), .o(g57121_sb) );
na02f02 TIMEBOOST_cell_71111 ( .a(TIMEBOOST_net_22763), .b(g62684_sb), .o(n_6171) );
na03f10 TIMEBOOST_cell_72384 ( .a(n_1409), .b(n_3007), .c(n_1549), .o(TIMEBOOST_net_17203) );
na02f02 TIMEBOOST_cell_70375 ( .a(TIMEBOOST_net_22395), .b(g63600_sb), .o(n_7189) );
in01f02 g57122_u0 ( .a(FE_OFN1383_n_8567), .o(g57122_sb) );
na02m04 TIMEBOOST_cell_69409 ( .a(TIMEBOOST_net_21912), .b(FE_OFN1058_n_4727), .o(TIMEBOOST_net_16959) );
na03f02 TIMEBOOST_cell_72390 ( .a(FE_RN_262_0), .b(n_5755), .c(TIMEBOOST_net_84), .o(TIMEBOOST_net_21322) );
na02m02 TIMEBOOST_cell_70343 ( .a(TIMEBOOST_net_22379), .b(g63606_sb), .o(n_7163) );
in01f02 g57123_u0 ( .a(FE_OFN1345_n_8567), .o(g57123_sb) );
na02m04 TIMEBOOST_cell_52258 ( .a(TIMEBOOST_net_16346), .b(g64337_db), .o(n_3840) );
in01f02 g57124_u0 ( .a(FE_OFN1419_n_8567), .o(g57124_sb) );
na04f04 TIMEBOOST_cell_35195 ( .a(n_10602), .b(n_10020), .c(n_10017), .d(n_10605), .o(n_12143) );
na03m06 TIMEBOOST_cell_72396 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .b(n_882), .c(n_1689), .o(n_883) );
na02s01 TIMEBOOST_cell_4298 ( .a(FE_OFN1022_n_11877), .b(g52472_da), .o(TIMEBOOST_net_709) );
in01f02 g57125_u0 ( .a(FE_OFN1415_n_8567), .o(g57125_sb) );
na02f01 TIMEBOOST_cell_53592 ( .a(TIMEBOOST_net_17013), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_15523) );
in01f02 g57126_u0 ( .a(FE_OFN1368_n_8567), .o(g57126_sb) );
na03s02 TIMEBOOST_cell_72550 ( .a(TIMEBOOST_net_13887), .b(g65734_sb), .c(g65734_db), .o(n_1934) );
na03s02 TIMEBOOST_cell_72394 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_98), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .c(g54205_sb), .o(TIMEBOOST_net_20793) );
na02s01 TIMEBOOST_cell_4302 ( .a(FE_OFN1021_n_11877), .b(g52464_da), .o(TIMEBOOST_net_711) );
in01f02 g57127_u0 ( .a(FE_OFN1401_n_8567), .o(g57127_sb) );
na03f02 TIMEBOOST_cell_66648 ( .a(TIMEBOOST_net_17074), .b(FE_OFN1231_n_6391), .c(g62346_sb), .o(n_6908) );
na02m02 TIMEBOOST_cell_71991 ( .a(TIMEBOOST_net_23203), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_10577) );
in01f02 g57128_u0 ( .a(FE_OFN1417_n_8567), .o(g57128_sb) );
na02f02 TIMEBOOST_cell_50933 ( .a(TIMEBOOST_net_7423), .b(FE_OFN1142_n_15261), .o(TIMEBOOST_net_15684) );
na02s02 TIMEBOOST_cell_48848 ( .a(TIMEBOOST_net_14641), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_9497) );
in01f02 g57129_u0 ( .a(FE_OFN1402_n_8567), .o(g57129_sb) );
na02f01 TIMEBOOST_cell_48001 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q), .b(n_3783), .o(TIMEBOOST_net_14218) );
na02f02 TIMEBOOST_cell_4307 ( .a(TIMEBOOST_net_713), .b(n_8896), .o(n_9931) );
na02s02 TIMEBOOST_cell_48012 ( .a(TIMEBOOST_net_14223), .b(g58036_sb), .o(TIMEBOOST_net_10380) );
in01f02 g57130_u0 ( .a(FE_OFN1417_n_8567), .o(g57130_sb) );
na03m04 TIMEBOOST_cell_72398 ( .a(n_1992), .b(n_245), .c(n_1993), .o(TIMEBOOST_net_126) );
na03m02 TIMEBOOST_cell_73497 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q), .b(FE_OFN231_n_9839), .c(FE_OFN575_n_9902), .o(TIMEBOOST_net_20559) );
in01f02 g57131_u0 ( .a(FE_OFN1377_n_8567), .o(g57131_sb) );
na02s02 TIMEBOOST_cell_48086 ( .a(TIMEBOOST_net_14260), .b(g58021_sb), .o(TIMEBOOST_net_10407) );
na03s02 TIMEBOOST_cell_72397 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_83), .b(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source), .c(g54167_sb), .o(TIMEBOOST_net_12275) );
na02s02 TIMEBOOST_cell_43786 ( .a(TIMEBOOST_net_12787), .b(FE_OFN1801_n_9690), .o(TIMEBOOST_net_11031) );
in01f02 g57132_u0 ( .a(FE_OFN1409_n_8567), .o(g57132_sb) );
na02m02 TIMEBOOST_cell_69317 ( .a(TIMEBOOST_net_21866), .b(TIMEBOOST_net_12504), .o(TIMEBOOST_net_17378) );
na02s01 TIMEBOOST_cell_31557 ( .a(FE_OFN1666_n_9477), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_9883) );
in01f02 g57133_u0 ( .a(FE_OFN1416_n_8567), .o(g57133_sb) );
na02s01 TIMEBOOST_cell_71308 ( .a(FE_OFN264_n_9849), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q), .o(TIMEBOOST_net_22862) );
na02s02 TIMEBOOST_cell_49459 ( .a(g57939_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q), .o(TIMEBOOST_net_14947) );
in01f02 g57134_u0 ( .a(FE_OFN1396_n_8567), .o(g57134_sb) );
na03f02 TIMEBOOST_cell_66882 ( .a(FE_OFN1566_n_12502), .b(TIMEBOOST_net_16482), .c(FE_OCPN1825_n_12030), .o(n_12525) );
na02m01 TIMEBOOST_cell_31559 ( .a(FE_OFN1690_n_9528), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_9884) );
in01f02 g57135_u0 ( .a(FE_OFN1413_n_8567), .o(g57135_sb) );
na03f02 TIMEBOOST_cell_35067 ( .a(TIMEBOOST_net_9613), .b(FE_OFN1437_n_9372), .c(g58466_sb), .o(n_9383) );
na04m02 TIMEBOOST_cell_67874 ( .a(n_4493), .b(g64909_sb), .c(g64909_db), .d(n_4403), .o(TIMEBOOST_net_17427) );
in01f02 g57136_u0 ( .a(FE_OFN1400_n_8567), .o(g57136_sb) );
na02m01 TIMEBOOST_cell_68264 ( .a(n_12179), .b(n_8486), .o(TIMEBOOST_net_21340) );
in01f02 g57137_u0 ( .a(FE_OFN2174_n_8567), .o(g57137_sb) );
na02m02 TIMEBOOST_cell_68336 ( .a(n_75), .b(n_3780), .o(TIMEBOOST_net_21376) );
in01s01 TIMEBOOST_cell_45989 ( .a(TIMEBOOST_net_13950), .o(TIMEBOOST_net_13853) );
in01f02 g57138_u0 ( .a(FE_OFN1425_n_8567), .o(g57138_sb) );
na03f02 TIMEBOOST_cell_35002 ( .a(TIMEBOOST_net_9572), .b(g57227_sb), .c(FE_OFN1383_n_8567), .o(n_11530) );
na03f02 TIMEBOOST_cell_66562 ( .a(TIMEBOOST_net_17483), .b(n_6319), .c(g62404_sb), .o(n_6791) );
in01f02 g57139_u0 ( .a(FE_OFN1411_n_8567), .o(g57139_sb) );
na03f02 TIMEBOOST_cell_67978 ( .a(TIMEBOOST_net_8841), .b(FE_OFN1183_n_3476), .c(g60636_sb), .o(n_5699) );
in01f02 g57140_u0 ( .a(FE_OFN1406_n_8567), .o(g57140_sb) );
na02s02 TIMEBOOST_cell_53492 ( .a(TIMEBOOST_net_16963), .b(FE_OFN1657_n_9502), .o(TIMEBOOST_net_11171) );
na03f02 TIMEBOOST_cell_73214 ( .a(FE_OCPN1875_n_14526), .b(n_16452), .c(n_7399), .o(TIMEBOOST_net_15048) );
in01f02 g57141_u0 ( .a(FE_OFN1423_n_8567), .o(g57141_sb) );
na03m02 TIMEBOOST_cell_68576 ( .a(g64814_db), .b(g64814_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q), .o(TIMEBOOST_net_21496) );
na02s02 TIMEBOOST_cell_43658 ( .a(TIMEBOOST_net_12723), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_11008) );
in01f02 g57142_u0 ( .a(FE_OFN1381_n_8567), .o(g57142_sb) );
in01s01 TIMEBOOST_cell_35482 ( .a(TIMEBOOST_net_10073), .o(wbs_dat_i_29_) );
na04f04 TIMEBOOST_cell_24528 ( .a(n_9783), .b(g57141_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q), .d(FE_OFN1423_n_8567), .o(n_11607) );
na02m06 TIMEBOOST_cell_68690 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q), .b(FE_OFN648_n_4497), .o(TIMEBOOST_net_21553) );
in01f02 g57143_u0 ( .a(FE_OFN1345_n_8567), .o(g57143_sb) );
na02m02 TIMEBOOST_cell_53048 ( .a(TIMEBOOST_net_16741), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_15290) );
na03f02 TIMEBOOST_cell_34896 ( .a(TIMEBOOST_net_9434), .b(FE_OFN1422_n_8567), .c(g57036_sb), .o(n_11696) );
in01f02 g57144_u0 ( .a(FE_OFN2167_n_8567), .o(g57144_sb) );
na03s02 TIMEBOOST_cell_41733 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q), .b(g58327_sb), .c(g58327_db), .o(n_9487) );
na03f02 TIMEBOOST_cell_73770 ( .a(TIMEBOOST_net_16054), .b(FE_OFN1774_n_13800), .c(FE_OFN1771_n_14054), .o(g53214_p) );
in01f02 g57145_u0 ( .a(FE_OFN1405_n_8567), .o(g57145_sb) );
na03f02 TIMEBOOST_cell_73356 ( .a(parchk_pci_cbe_out_in_1202), .b(FE_OFN1705_n_4868), .c(g59093_sb), .o(TIMEBOOST_net_15661) );
na04f08 TIMEBOOST_cell_73151 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q), .b(FE_OFN1074_n_4740), .c(pci_target_unit_fifos_pciw_cbe_in), .d(g64111_sb), .o(n_4741) );
na03f20 TIMEBOOST_cell_72366 ( .a(conf_wb_err_addr_in_947), .b(conf_wb_err_addr_in_950), .c(n_1165), .o(n_1972) );
in01f02 g57146_u0 ( .a(FE_OFN2182_n_8567), .o(g57146_sb) );
na02f02 TIMEBOOST_cell_70055 ( .a(TIMEBOOST_net_22235), .b(g61712_sb), .o(n_8402) );
in01s01 TIMEBOOST_cell_45986 ( .a(TIMEBOOST_net_13947), .o(TIMEBOOST_net_13946) );
na03f02 TIMEBOOST_cell_73283 ( .a(TIMEBOOST_net_8783), .b(g62746_sb), .c(FE_OFN1118_g64577_p), .o(n_5489) );
in01f02 g57147_u0 ( .a(FE_OFN1409_n_8567), .o(g57147_sb) );
na04f04 TIMEBOOST_cell_35004 ( .a(n_9706), .b(g57233_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q), .d(FE_OFN1392_n_8567), .o(n_11521) );
na03f04 TIMEBOOST_cell_73336 ( .a(TIMEBOOST_net_17344), .b(FE_OCPN1911_FE_OFN1152_n_13249), .c(g54148_sb), .o(n_13661) );
in01f02 g57148_u0 ( .a(FE_OFN1345_n_8567), .o(g57148_sb) );
in01s01 TIMEBOOST_cell_67756 ( .a(TIMEBOOST_net_21182), .o(TIMEBOOST_net_21183) );
na03m08 TIMEBOOST_cell_72996 ( .a(TIMEBOOST_net_17254), .b(FE_OFN1046_n_16657), .c(g64110_sb), .o(n_4047) );
na03f02 TIMEBOOST_cell_35001 ( .a(TIMEBOOST_net_9571), .b(FE_OFN2171_n_8567), .c(FE_OFN2177_n_8567), .o(n_11682) );
in01f02 g57149_u0 ( .a(FE_OFN1388_n_8567), .o(g57149_sb) );
in01s01 TIMEBOOST_cell_35483 ( .a(TIMEBOOST_net_10074), .o(TIMEBOOST_net_10073) );
na02f02 TIMEBOOST_cell_49932 ( .a(TIMEBOOST_net_15183), .b(g63115_sb), .o(n_5025) );
in01f02 g57150_u0 ( .a(FE_OFN1421_n_8567), .o(g57150_sb) );
na02m08 TIMEBOOST_cell_52961 ( .a(wishbone_slave_unit_pcim_sm_data_in_649), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q), .o(TIMEBOOST_net_16698) );
na03f02 TIMEBOOST_cell_67904 ( .a(TIMEBOOST_net_16935), .b(FE_OFN1056_n_4727), .c(g64238_sb), .o(TIMEBOOST_net_13079) );
in01f02 g57151_u0 ( .a(FE_OFN1406_n_8567), .o(g57151_sb) );
na03f02 TIMEBOOST_cell_66805 ( .a(TIMEBOOST_net_16847), .b(FE_OFN1345_n_8567), .c(g57178_sb), .o(n_11577) );
in01s01 TIMEBOOST_cell_35484 ( .a(TIMEBOOST_net_10075), .o(wbs_dat_i_5_) );
na04s02 TIMEBOOST_cell_33416 ( .a(g58149_sb), .b(FE_OFN266_n_9884), .c(g58149_db), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q), .o(TIMEBOOST_net_9507) );
in01f02 g57152_u0 ( .a(FE_OFN1392_n_8567), .o(g57152_sb) );
in01s01 TIMEBOOST_cell_35486 ( .a(TIMEBOOST_net_10077), .o(wbs_dat_i_18_) );
na03f02 TIMEBOOST_cell_34785 ( .a(TIMEBOOST_net_9530), .b(FE_OFN1383_n_8567), .c(g57381_sb), .o(n_11365) );
in01f02 g57153_u0 ( .a(FE_OFN1389_n_8567), .o(g57153_sb) );
na04f02 TIMEBOOST_cell_67595 ( .a(conf_wb_err_addr_in_963), .b(g62123_sb), .c(configuration_wb_err_addr_554), .d(FE_OFN1170_n_5592), .o(n_5573) );
na03f02 TIMEBOOST_cell_73799 ( .a(n_13997), .b(TIMEBOOST_net_8118), .c(FE_OFN1602_n_13995), .o(g53268_p) );
in01f02 g57154_u0 ( .a(FE_OFN2191_n_8567), .o(g57154_sb) );
na03m02 TIMEBOOST_cell_67958 ( .a(TIMEBOOST_net_15028), .b(g62729_sb), .c(FE_OFN1139_g64577_p), .o(n_5521) );
na03f04 TIMEBOOST_cell_72458 ( .a(TIMEBOOST_net_534), .b(n_4078), .c(n_3337), .o(n_4080) );
na02m02 TIMEBOOST_cell_48863 ( .a(g58096_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q), .o(TIMEBOOST_net_14649) );
in01f02 g57155_u0 ( .a(FE_OFN1424_n_8567), .o(g57155_sb) );
na03f02 TIMEBOOST_cell_70182 ( .a(TIMEBOOST_net_12850), .b(FE_OFN2127_n_16497), .c(g54039_sb), .o(TIMEBOOST_net_22299) );
na02s01 TIMEBOOST_cell_62449 ( .a(TIMEBOOST_net_20171), .b(FE_OFN1786_n_1699), .o(TIMEBOOST_net_16155) );
in01f02 g57156_u0 ( .a(FE_OFN1380_n_8567), .o(g57156_sb) );
na03m02 TIMEBOOST_cell_72760 ( .a(TIMEBOOST_net_21598), .b(g65078_sb), .c(TIMEBOOST_net_21994), .o(TIMEBOOST_net_21028) );
na03m02 TIMEBOOST_cell_72869 ( .a(TIMEBOOST_net_21731), .b(g64767_sb), .c(TIMEBOOST_net_21972), .o(TIMEBOOST_net_17153) );
na03f02 TIMEBOOST_cell_66965 ( .a(FE_OCP_RBN1973_n_12381), .b(TIMEBOOST_net_16512), .c(FE_OFN1755_n_12681), .o(n_12713) );
in01f02 g57157_u0 ( .a(FE_OFN2191_n_8567), .o(g57157_sb) );
na02f04 TIMEBOOST_cell_50711 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_389), .b(FE_OFN2070_n_15978), .o(TIMEBOOST_net_15573) );
na02m06 TIMEBOOST_cell_68989 ( .a(TIMEBOOST_net_21702), .b(g64865_sb), .o(TIMEBOOST_net_9763) );
in01f02 g57158_u0 ( .a(FE_OFN1345_n_8567), .o(g57158_sb) );
na02s02 TIMEBOOST_cell_39183 ( .a(TIMEBOOST_net_11203), .b(g58048_db), .o(n_9741) );
na02f01 TIMEBOOST_cell_26119 ( .a(pci_target_unit_pcit_if_strd_addr_in_708), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7164) );
na02m02 g61987_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61987_db) );
in01f02 g57159_u0 ( .a(FE_OFN1384_n_8567), .o(g57159_sb) );
na03m02 TIMEBOOST_cell_72860 ( .a(TIMEBOOST_net_21695), .b(g65036_sb), .c(TIMEBOOST_net_21958), .o(TIMEBOOST_net_20980) );
na03m02 TIMEBOOST_cell_70080 ( .a(n_4450), .b(g64864_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q), .o(TIMEBOOST_net_22248) );
in01f02 g57160_u0 ( .a(FE_OFN1345_n_8567), .o(g57160_sb) );
na02m02 TIMEBOOST_cell_70881 ( .a(TIMEBOOST_net_22648), .b(g57932_sb), .o(n_9878) );
na02s02 TIMEBOOST_cell_48504 ( .a(TIMEBOOST_net_14469), .b(g57998_db), .o(TIMEBOOST_net_9477) );
na02m02 g62021_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g62021_db) );
in01f02 g57161_u0 ( .a(FE_OFN1368_n_8567), .o(g57161_sb) );
na03f02 TIMEBOOST_cell_66867 ( .a(n_12228), .b(FE_OFN1749_n_12004), .c(TIMEBOOST_net_13522), .o(n_12707) );
na02s01 TIMEBOOST_cell_37609 ( .a(TIMEBOOST_net_10416), .b(g58154_db), .o(n_9637) );
na02s01 TIMEBOOST_cell_48161 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_14298) );
in01f02 g57162_u0 ( .a(FE_OFN1401_n_8567), .o(g57162_sb) );
na02m04 TIMEBOOST_cell_54063 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q), .b(pci_target_unit_fifos_pciw_cbe_in), .o(TIMEBOOST_net_17249) );
in01f02 g57163_u0 ( .a(FE_OFN2169_n_8567), .o(g57163_sb) );
na03f02 TIMEBOOST_cell_66568 ( .a(TIMEBOOST_net_17129), .b(FE_OFN1310_n_6624), .c(g62408_sb), .o(n_6783) );
na02m04 TIMEBOOST_cell_68622 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q), .o(TIMEBOOST_net_21519) );
in01f02 g57164_u0 ( .a(FE_OFN1377_n_8567), .o(g57164_sb) );
na03f01 TIMEBOOST_cell_65096 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q), .c(FE_OFN686_n_4417), .o(TIMEBOOST_net_16253) );
na04f04 TIMEBOOST_cell_24530 ( .a(n_9788), .b(g57138_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q), .d(FE_OFN1425_n_8567), .o(n_11611) );
na04f04 TIMEBOOST_cell_36842 ( .a(n_9095), .b(g57177_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q), .d(FE_OFN1398_n_8567), .o(n_10451) );
in01f02 g57165_u0 ( .a(FE_OFN1416_n_8567), .o(g57165_sb) );
na02f02 TIMEBOOST_cell_71068 ( .a(TIMEBOOST_net_17577), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_22742) );
na04f04 TIMEBOOST_cell_36843 ( .a(n_9563), .b(g57369_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q), .d(FE_OFN1397_n_8567), .o(n_11381) );
na02f02 TIMEBOOST_cell_49832 ( .a(TIMEBOOST_net_15133), .b(g63019_sb), .o(n_5210) );
in01f02 g57166_u0 ( .a(FE_OFN1377_n_8567), .o(g57166_sb) );
na02s01 TIMEBOOST_cell_68778 ( .a(n_3780), .b(g64752_sb), .o(TIMEBOOST_net_21597) );
na03m02 TIMEBOOST_cell_64601 ( .a(FE_OFN624_n_4409), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q), .c(n_3774), .o(TIMEBOOST_net_10572) );
in01f02 g57167_u0 ( .a(FE_OFN1409_n_8567), .o(g57167_sb) );
na02f01 TIMEBOOST_cell_70538 ( .a(TIMEBOOST_net_13110), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_22477) );
na03f02 TIMEBOOST_cell_73498 ( .a(g60634_sb), .b(wbm_adr_o_8_), .c(TIMEBOOST_net_11652), .o(n_5702) );
in01f02 g57168_u0 ( .a(FE_OFN1396_n_8567), .o(g57168_sb) );
na04m02 TIMEBOOST_cell_72775 ( .a(TIMEBOOST_net_20332), .b(n_4444), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q), .d(g65391_sb), .o(TIMEBOOST_net_17570) );
na02s01 TIMEBOOST_cell_43750 ( .a(TIMEBOOST_net_12769), .b(g58111_db), .o(n_9077) );
in01f02 g57169_u0 ( .a(FE_OFN1416_n_8567), .o(g57169_sb) );
na03f02 TIMEBOOST_cell_73357 ( .a(parchk_pci_cbe_out_in_1203), .b(FE_OFN1705_n_4868), .c(g52877_sb), .o(TIMEBOOST_net_7998) );
na02m01 TIMEBOOST_cell_63306 ( .a(n_8272), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_20600) );
na02f02 TIMEBOOST_cell_39109 ( .a(TIMEBOOST_net_11166), .b(g64253_da), .o(TIMEBOOST_net_9913) );
in01f02 g57170_u0 ( .a(FE_OFN1413_n_8567), .o(g57170_sb) );
na04f04 TIMEBOOST_cell_24284 ( .a(n_9604), .b(g57324_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q), .d(FE_OFN1424_n_8567), .o(n_11425) );
in01f02 g57171_u0 ( .a(FE_OFN1370_n_8567), .o(g57171_sb) );
in01s01 TIMEBOOST_cell_73873 ( .a(TIMEBOOST_net_23437), .o(TIMEBOOST_net_23438) );
na04m08 TIMEBOOST_cell_67293 ( .a(n_4645), .b(FE_OFN647_n_4497), .c(g64974_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q), .o(n_4369) );
in01f02 g57172_u0 ( .a(FE_OFN2173_n_8567), .o(g57172_sb) );
na02m02 TIMEBOOST_cell_68814 ( .a(n_4488), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q), .o(TIMEBOOST_net_21615) );
in01f02 g57173_u0 ( .a(FE_OFN1425_n_8567), .o(g57173_sb) );
na02f02 TIMEBOOST_cell_53630 ( .a(TIMEBOOST_net_17032), .b(FE_OFN1252_n_4143), .o(TIMEBOOST_net_15431) );
na03m04 TIMEBOOST_cell_47242 ( .a(FE_OFN1566_n_12502), .b(TIMEBOOST_net_13527), .c(n_12313), .o(n_12660) );
na02s01 TIMEBOOST_cell_43752 ( .a(TIMEBOOST_net_12770), .b(FE_OFN233_n_9876), .o(n_9763) );
in01f02 g57174_u0 ( .a(FE_OFN1427_n_8567), .o(g57174_sb) );
na02m04 TIMEBOOST_cell_68656 ( .a(g64798_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q), .o(TIMEBOOST_net_21536) );
no02f20 TIMEBOOST_cell_37137 ( .a(TIMEBOOST_net_10180), .b(n_832), .o(g65808_p) );
in01f02 g57175_u0 ( .a(FE_OFN2177_n_8567), .o(g57175_sb) );
na03m02 TIMEBOOST_cell_69864 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q), .b(pci_target_unit_fifos_pciw_cbe_in_153), .c(FE_OFN912_n_4727), .o(TIMEBOOST_net_22140) );
na03f02 TIMEBOOST_cell_66638 ( .a(TIMEBOOST_net_8538), .b(FE_OCPN1847_n_14981), .c(g59098_sb), .o(n_8713) );
in01f02 g57176_u0 ( .a(FE_OFN1408_n_8567), .o(g57176_sb) );
na02m02 TIMEBOOST_cell_68782 ( .a(FE_OFN1625_n_4438), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q), .o(TIMEBOOST_net_21599) );
na04f04 TIMEBOOST_cell_24286 ( .a(n_9612), .b(g57320_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q), .d(FE_OFN1389_n_8567), .o(n_11431) );
na02s01 TIMEBOOST_cell_4376 ( .a(FE_OFN1021_n_11877), .b(g52468_da), .o(TIMEBOOST_net_748) );
in01f02 g57177_u0 ( .a(FE_OFN1370_n_8567), .o(g57177_sb) );
na03f02 TIMEBOOST_cell_72678 ( .a(TIMEBOOST_net_16185), .b(FE_OFN787_n_2678), .c(g65230_sb), .o(n_2657) );
na03f02 TIMEBOOST_cell_66592 ( .a(TIMEBOOST_net_17433), .b(FE_OFN1218_n_6886), .c(g62624_sb), .o(n_6308) );
in01f02 g57178_u0 ( .a(FE_OFN1345_n_8567), .o(g57178_sb) );
na03m02 TIMEBOOST_cell_73039 ( .a(TIMEBOOST_net_23211), .b(FE_OFN1677_n_4655), .c(TIMEBOOST_net_22060), .o(TIMEBOOST_net_20536) );
na02m02 g61974_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61974_db) );
in01f02 g57179_u0 ( .a(FE_OFN2180_n_8567), .o(g57179_sb) );
na02f02 TIMEBOOST_cell_47926 ( .a(TIMEBOOST_net_14180), .b(FE_OFN918_n_4725), .o(TIMEBOOST_net_12478) );
na02s02 TIMEBOOST_cell_37141 ( .a(TIMEBOOST_net_10182), .b(FE_OFN935_n_2292), .o(TIMEBOOST_net_8199) );
na03s02 TIMEBOOST_cell_46433 ( .a(TIMEBOOST_net_12458), .b(g58236_sb), .c(TIMEBOOST_net_12711), .o(TIMEBOOST_net_9333) );
in01f02 g57180_u0 ( .a(FE_OFN1406_n_8567), .o(g57180_sb) );
na02m02 TIMEBOOST_cell_68786 ( .a(TIMEBOOST_net_12381), .b(FE_OFN917_n_4725), .o(TIMEBOOST_net_21601) );
in01s01 TIMEBOOST_cell_35488 ( .a(TIMEBOOST_net_10079), .o(wbs_dat_i_19_) );
na03f02 TIMEBOOST_cell_66807 ( .a(TIMEBOOST_net_16838), .b(FE_OFN1344_n_8567), .c(g57300_sb), .o(n_11451) );
in01f01 g57181_u0 ( .a(FE_OFN1394_n_8567), .o(g57181_sb) );
na03s01 TIMEBOOST_cell_64711 ( .a(pci_target_unit_del_sync_addr_in_234), .b(g66415_sb), .c(g66429_db), .o(n_2497) );
na02s02 TIMEBOOST_cell_70463 ( .a(TIMEBOOST_net_22439), .b(TIMEBOOST_net_20513), .o(TIMEBOOST_net_16428) );
in01f02 g57182_u0 ( .a(FE_OFN1408_n_8567), .o(g57182_sb) );
na02f02 TIMEBOOST_cell_69079 ( .a(TIMEBOOST_net_21747), .b(TIMEBOOST_net_14389), .o(TIMEBOOST_net_13377) );
na03f02 TIMEBOOST_cell_66685 ( .a(TIMEBOOST_net_13368), .b(n_6232), .c(g62973_sb), .o(n_5936) );
in01f02 g57183_u0 ( .a(FE_OFN1387_n_8567), .o(g57183_sb) );
na02m02 TIMEBOOST_cell_50250 ( .a(TIMEBOOST_net_15342), .b(g62568_sb), .o(n_6420) );
in01f02 g57184_u0 ( .a(FE_OFN1349_n_8567), .o(g57184_sb) );
na02s02 TIMEBOOST_cell_43364 ( .a(FE_OFN588_n_9692), .b(TIMEBOOST_net_12576), .o(TIMEBOOST_net_10627) );
na02m08 TIMEBOOST_cell_54111 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_142), .o(TIMEBOOST_net_17273) );
na02m02 g61976_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61976_db) );
in01f02 g57185_u0 ( .a(FE_OFN1391_n_8567), .o(g57185_sb) );
na04f04 TIMEBOOST_cell_73535 ( .a(n_3677), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q), .c(FE_OFN1233_n_6391), .d(g62644_sb), .o(n_6261) );
na03f02 TIMEBOOST_cell_73598 ( .a(TIMEBOOST_net_17429), .b(FE_OFN1270_n_4095), .c(g62555_sb), .o(n_6453) );
in01f02 g57186_u0 ( .a(FE_OFN1406_n_8567), .o(g57186_sb) );
na03f02 TIMEBOOST_cell_66637 ( .a(g62755_sb), .b(FE_OFN1233_n_6391), .c(TIMEBOOST_net_16764), .o(n_6127) );
na04m04 TIMEBOOST_cell_72606 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q), .c(FE_OFN1640_n_4671), .d(g65916_sb), .o(n_1852) );
in01s01 TIMEBOOST_cell_72360 ( .a(pci_target_unit_fifos_pcir_data_in_168), .o(TIMEBOOST_net_23393) );
in01f02 g57187_u0 ( .a(FE_OFN1392_n_8567), .o(g57187_sb) );
na02f02 TIMEBOOST_cell_37213 ( .a(TIMEBOOST_net_10218), .b(n_2125), .o(n_4720) );
na02m02 TIMEBOOST_cell_69444 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q), .b(g65032_sb), .o(TIMEBOOST_net_21930) );
na04f02 TIMEBOOST_cell_67956 ( .a(n_14741), .b(n_14839), .c(TIMEBOOST_net_20992), .d(g52449_sb), .o(n_14842) );
in01f02 g57188_u0 ( .a(FE_OFN1389_n_8567), .o(g57188_sb) );
na02s02 TIMEBOOST_cell_49229 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q), .b(g65882_sb), .o(TIMEBOOST_net_14832) );
na02f06 TIMEBOOST_cell_43690 ( .a(TIMEBOOST_net_12739), .b(n_2691), .o(n_2915) );
in01f02 g57189_u0 ( .a(FE_OFN1387_n_8567), .o(g57189_sb) );
na03f02 TIMEBOOST_cell_65221 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q), .b(FE_OFN1689_n_9528), .c(g58300_sb), .o(TIMEBOOST_net_14929) );
in01f02 g57190_u0 ( .a(FE_OFN1387_n_8567), .o(g57190_sb) );
na02m08 TIMEBOOST_cell_71965 ( .a(TIMEBOOST_net_23190), .b(g65402_sb), .o(TIMEBOOST_net_12597) );
in01f02 g57191_u0 ( .a(FE_OFN1382_n_8567), .o(g57191_sb) );
na04m06 TIMEBOOST_cell_67220 ( .a(n_4479), .b(FE_OFN682_n_4460), .c(g64820_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q), .o(n_4456) );
na02s01 TIMEBOOST_cell_52897 ( .a(parchk_pci_ad_out_in_1197), .b(configuration_wb_err_data_600), .o(TIMEBOOST_net_16666) );
in01f02 g57192_u0 ( .a(FE_OFN1387_n_8567), .o(g57192_sb) );
na03f02 TIMEBOOST_cell_72729 ( .a(TIMEBOOST_net_16207), .b(FE_OFN1797_n_2299), .c(g65970_sb), .o(n_2154) );
na03f02 TIMEBOOST_cell_47244 ( .a(FE_OFN1566_n_12502), .b(TIMEBOOST_net_13524), .c(n_12313), .o(n_12762) );
in01s02 TIMEBOOST_cell_67796 ( .a(TIMEBOOST_net_21223), .o(TIMEBOOST_net_21222) );
in01f02 g57193_u0 ( .a(FE_OFN1385_n_8567), .o(g57193_sb) );
na02s04 TIMEBOOST_cell_68102 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_94), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_21259) );
na04f03 TIMEBOOST_cell_24538 ( .a(n_337), .b(FE_OFN2185_n_8567), .c(n_8551), .d(g58610_sb), .o(n_9188) );
in01f02 g57194_u0 ( .a(FE_OFN2177_n_8567), .o(g57194_sb) );
na02f01 TIMEBOOST_cell_39434 ( .a(TIMEBOOST_net_8343), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_11329) );
na02s02 TIMEBOOST_cell_37249 ( .a(TIMEBOOST_net_10236), .b(g65700_sb), .o(n_2202) );
in01f02 g57195_u0 ( .a(FE_OFN1385_n_8567), .o(g57195_sb) );
na03f02 TIMEBOOST_cell_73599 ( .a(TIMEBOOST_net_17428), .b(FE_OFN1212_n_4151), .c(g62389_sb), .o(n_6821) );
na02f04 TIMEBOOST_cell_4397 ( .a(FE_OCP_RBN1983_FE_OFN1591_n_13741), .b(TIMEBOOST_net_758), .o(g53182_p) );
in01f02 g57196_u0 ( .a(FE_OFN1412_n_8567), .o(g57196_sb) );
na03f02 TIMEBOOST_cell_73812 ( .a(TIMEBOOST_net_13781), .b(FE_OFN1775_n_13800), .c(FE_OFN1768_n_14054), .o(n_14436) );
na02f04 TIMEBOOST_cell_4399 ( .a(FE_OCP_RBN1981_FE_OFN1591_n_13741), .b(TIMEBOOST_net_759), .o(g53170_p) );
in01f02 g57197_u0 ( .a(FE_OFN1401_n_8567), .o(g57197_sb) );
na02f04 TIMEBOOST_cell_4401 ( .a(FE_OCP_RBN1985_FE_OFN1591_n_13741), .b(TIMEBOOST_net_760), .o(g53158_p) );
in01f02 g57198_u0 ( .a(FE_OFN1373_n_8567), .o(g57198_sb) );
na02s01 TIMEBOOST_cell_70734 ( .a(FE_OFN1650_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q), .o(TIMEBOOST_net_22575) );
na02f02 TIMEBOOST_cell_70299 ( .a(TIMEBOOST_net_22357), .b(g54153_sb), .o(n_13658) );
in01f02 g57199_u0 ( .a(FE_OFN1427_n_8567), .o(g57199_sb) );
na02m02 TIMEBOOST_cell_63655 ( .a(TIMEBOOST_net_20813), .b(FE_OFN1011_n_4734), .o(TIMEBOOST_net_14428) );
na02s02 TIMEBOOST_cell_68191 ( .a(TIMEBOOST_net_21303), .b(g65810_sb), .o(n_2163) );
na02s02 TIMEBOOST_cell_37376 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(g65777_sb), .o(TIMEBOOST_net_10300) );
in01f02 g57200_u0 ( .a(FE_OFN1405_n_8567), .o(g57200_sb) );
na04f02 TIMEBOOST_cell_65842 ( .a(TIMEBOOST_net_7313), .b(g54318_sb), .c(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q), .d(FE_OCPN1909_n_16497), .o(n_13290) );
na02m01 TIMEBOOST_cell_48341 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_14388) );
na02f04 TIMEBOOST_cell_51449 ( .a(pci_target_unit_pcit_if_strd_addr_in_691), .b(g52650_sb), .o(TIMEBOOST_net_15942) );
in01f02 g57201_u0 ( .a(FE_OFN1402_n_8567), .o(g57201_sb) );
na02s02 TIMEBOOST_cell_71307 ( .a(TIMEBOOST_net_22861), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_11207) );
na02f02 TIMEBOOST_cell_4403 ( .a(FE_OCP_RBN1984_FE_OFN1591_n_13741), .b(TIMEBOOST_net_761), .o(g53211_p) );
in01f02 g57202_u0 ( .a(FE_OFN1399_n_8567), .o(g57202_sb) );
na03m04 TIMEBOOST_cell_73600 ( .a(g54195_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_414), .c(TIMEBOOST_net_655), .o(n_13423) );
na02f04 TIMEBOOST_cell_4405 ( .a(FE_OCP_RBN1985_FE_OFN1591_n_13741), .b(TIMEBOOST_net_762), .o(g74859_p) );
in01f01 g57203_u0 ( .a(FE_OFN1394_n_8567), .o(g57203_sb) );
na02m01 TIMEBOOST_cell_44065 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q), .o(TIMEBOOST_net_12927) );
in01f02 g57204_u0 ( .a(FE_OFN1384_n_8567), .o(g57204_sb) );
na03f02 TIMEBOOST_cell_35006 ( .a(TIMEBOOST_net_9574), .b(g57523_sb), .c(FE_OFN1376_n_8567), .o(n_11218) );
na02f02 TIMEBOOST_cell_4407 ( .a(FE_OCP_RBN1984_FE_OFN1591_n_13741), .b(TIMEBOOST_net_763), .o(g53230_p) );
in01f02 g57205_u0 ( .a(FE_OFN1412_n_8567), .o(g57205_sb) );
na04f04 TIMEBOOST_cell_35008 ( .a(n_9546), .b(g57390_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q), .d(FE_OFN1383_n_8567), .o(n_11353) );
na02f04 TIMEBOOST_cell_4409 ( .a(FE_OCP_RBN1985_FE_OFN1591_n_13741), .b(TIMEBOOST_net_764), .o(g53251_p) );
na02s06 TIMEBOOST_cell_68251 ( .a(TIMEBOOST_net_21333), .b(wbu_addr_in_260), .o(TIMEBOOST_net_10332) );
in01f02 g57206_u0 ( .a(FE_OFN1400_n_8567), .o(g57206_sb) );
na02s01 TIMEBOOST_cell_48157 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q), .o(TIMEBOOST_net_14296) );
in01f02 g57207_u0 ( .a(FE_OFN1427_n_8567), .o(g57207_sb) );
na02f02 TIMEBOOST_cell_51450 ( .a(TIMEBOOST_net_15942), .b(n_14837), .o(TIMEBOOST_net_11884) );
na02f08 TIMEBOOST_cell_37217 ( .a(TIMEBOOST_net_10220), .b(n_2428), .o(n_2429) );
na02s01 TIMEBOOST_cell_45375 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q), .o(TIMEBOOST_net_13582) );
in01f02 g57208_u0 ( .a(FE_OFN1425_n_8567), .o(g57208_sb) );
na02s02 TIMEBOOST_cell_68777 ( .a(TIMEBOOST_net_21596), .b(g65682_sb), .o(n_1955) );
na02s02 TIMEBOOST_cell_37607 ( .a(TIMEBOOST_net_10415), .b(g58051_db), .o(n_9737) );
na02s01 TIMEBOOST_cell_4414 ( .a(g52482_da), .b(FE_OFN8_n_11877), .o(TIMEBOOST_net_767) );
in01f02 g57209_u0 ( .a(FE_OFN1420_n_8567), .o(g57209_sb) );
na02m20 TIMEBOOST_cell_53191 ( .a(pci_target_unit_pcit_if_strd_addr_in_714), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78), .o(TIMEBOOST_net_16813) );
na02m02 TIMEBOOST_cell_63175 ( .a(TIMEBOOST_net_20534), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_15362) );
na03f06 TIMEBOOST_cell_66869 ( .a(n_12228), .b(FE_OFN1749_n_12004), .c(TIMEBOOST_net_21084), .o(n_15441) );
in01f02 g57210_u0 ( .a(FE_OFN1407_n_8567), .o(g57210_sb) );
na02f01 TIMEBOOST_cell_70058 ( .a(FE_OFN707_n_8119), .b(TIMEBOOST_net_14594), .o(TIMEBOOST_net_22237) );
na02s01 TIMEBOOST_cell_62448 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q), .o(TIMEBOOST_net_20171) );
na02m01 TIMEBOOST_cell_62596 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q), .b(n_3739), .o(TIMEBOOST_net_20245) );
in01f02 g57211_u0 ( .a(FE_OFN1422_n_8567), .o(g57211_sb) );
na03m02 TIMEBOOST_cell_72589 ( .a(TIMEBOOST_net_23148), .b(g64778_sb), .c(TIMEBOOST_net_21628), .o(TIMEBOOST_net_16773) );
na04f04 TIMEBOOST_cell_24667 ( .a(n_9501), .b(g57446_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q), .d(FE_OFN2188_n_8567), .o(n_11286) );
in01s08 TIMEBOOST_cell_67795 ( .a(TIMEBOOST_net_21222), .o(FE_OFN606_n_9904) );
in01f02 g57212_u0 ( .a(FE_OFN1397_n_8567), .o(g57212_sb) );
na03f02 TIMEBOOST_cell_73601 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_405), .b(g54186_sb), .c(TIMEBOOST_net_650), .o(n_13429) );
na02f02 TIMEBOOST_cell_4419 ( .a(TIMEBOOST_net_769), .b(n_8926), .o(n_9947) );
in01f02 g57213_u0 ( .a(FE_OFN1374_n_8567), .o(g57213_sb) );
na02s02 TIMEBOOST_cell_48630 ( .a(TIMEBOOST_net_14532), .b(g57986_sb), .o(TIMEBOOST_net_9568) );
na02s02 TIMEBOOST_cell_48109 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q), .b(FE_OFN1785_n_1699), .o(TIMEBOOST_net_14272) );
na03m06 TIMEBOOST_cell_67160 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q), .b(n_3749), .c(FE_OFN615_n_4501), .o(TIMEBOOST_net_10581) );
in01f02 g57214_u0 ( .a(FE_OFN2168_n_8567), .o(g57214_sb) );
na02s01 TIMEBOOST_cell_37448 ( .a(pci_target_unit_fifos_pcir_data_in), .b(g65761_sb), .o(TIMEBOOST_net_10336) );
na02m02 TIMEBOOST_cell_45133 ( .a(TIMEBOOST_net_8844), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_13461) );
in01f02 g57215_u0 ( .a(FE_OFN2168_n_8567), .o(g57215_sb) );
na02m10 TIMEBOOST_cell_52963 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q), .b(wishbone_slave_unit_pcim_sm_data_in_636), .o(TIMEBOOST_net_16699) );
na04f04 TIMEBOOST_cell_24656 ( .a(n_9086), .b(g57214_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q), .d(FE_OFN2168_n_8567), .o(n_10438) );
na02s01 TIMEBOOST_cell_4424 ( .a(FE_OFN1022_n_11877), .b(g52459_da), .o(TIMEBOOST_net_772) );
in01f02 g57216_u0 ( .a(FE_OFN1376_n_8567), .o(g57216_sb) );
na03f02 TIMEBOOST_cell_67032 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_13753), .c(FE_OFN1599_n_13995), .o(n_14437) );
na04f04 TIMEBOOST_cell_24658 ( .a(n_9232), .b(g57060_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q), .d(FE_OFN2174_n_8567), .o(n_10847) );
na02s01 TIMEBOOST_cell_4426 ( .a(FE_OFN1021_n_11877), .b(g52462_da), .o(TIMEBOOST_net_773) );
in01f02 g57217_u0 ( .a(FE_OFN1423_n_8567), .o(g57217_sb) );
na02s01 TIMEBOOST_cell_45377 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q), .o(TIMEBOOST_net_13583) );
na04f04 TIMEBOOST_cell_24660 ( .a(n_9733), .b(g57194_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q), .d(FE_OFN2177_n_8567), .o(n_11559) );
na02m02 TIMEBOOST_cell_54732 ( .a(TIMEBOOST_net_17583), .b(TIMEBOOST_net_12764), .o(TIMEBOOST_net_9447) );
in01f02 g57218_u0 ( .a(FE_OFN1389_n_8567), .o(g57218_sb) );
na03f02 TIMEBOOST_cell_65496 ( .a(FE_OFN712_n_8140), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q), .c(n_1905), .o(TIMEBOOST_net_14870) );
na02s01 TIMEBOOST_cell_4430 ( .a(g52456_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_775) );
in01f02 g57219_u0 ( .a(FE_OFN1349_n_8567), .o(g57219_sb) );
na03f02 TIMEBOOST_cell_66452 ( .a(TIMEBOOST_net_17109), .b(FE_OFN1312_n_6624), .c(g62912_sb), .o(n_6054) );
na02m02 TIMEBOOST_cell_68562 ( .a(FE_OFN634_n_4454), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_21489) );
na02m02 g61980_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61980_db) );
in01f02 g57220_u0 ( .a(FE_OFN1421_n_8567), .o(g57220_sb) );
in01s01 TIMEBOOST_cell_35490 ( .a(TIMEBOOST_net_10081), .o(wbs_dat_i_16_) );
na03f02 TIMEBOOST_cell_67010 ( .a(FE_OFN1586_n_13736), .b(n_13993), .c(TIMEBOOST_net_13720), .o(n_14422) );
na02s01 TIMEBOOST_cell_45437 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q), .o(TIMEBOOST_net_13613) );
in01f02 g57221_u0 ( .a(FE_OFN2177_n_8567), .o(g57221_sb) );
in01s04 TIMEBOOST_cell_67797 ( .a(TIMEBOOST_net_21224), .o(FE_OFN540_n_9690) );
na02f02 TIMEBOOST_cell_54670 ( .a(TIMEBOOST_net_17552), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_15480) );
in01f02 g57222_u0 ( .a(FE_OFN1390_n_8567), .o(g57222_sb) );
in01m02 TIMEBOOST_cell_45915 ( .a(TIMEBOOST_net_13925), .o(TIMEBOOST_net_13876) );
na02m04 TIMEBOOST_cell_72091 ( .a(TIMEBOOST_net_23253), .b(FE_OFN923_n_4740), .o(TIMEBOOST_net_22284) );
na02m02 TIMEBOOST_cell_63279 ( .a(TIMEBOOST_net_20586), .b(TIMEBOOST_net_12736), .o(TIMEBOOST_net_9392) );
in01f02 g57223_u0 ( .a(FE_OFN1407_n_8567), .o(g57223_sb) );
no02f02 TIMEBOOST_cell_4433 ( .a(TIMEBOOST_net_776), .b(n_13564), .o(g53012_p) );
na02s01 TIMEBOOST_cell_48905 ( .a(FE_OFN235_n_9834), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q), .o(TIMEBOOST_net_14670) );
in01f02 g57224_u0 ( .a(FE_OFN2187_n_8567), .o(g57224_sb) );
na02s01 TIMEBOOST_cell_48717 ( .a(FE_OFN554_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q), .o(TIMEBOOST_net_14576) );
na02m01 TIMEBOOST_cell_37041 ( .a(TIMEBOOST_net_10132), .b(n_574), .o(TIMEBOOST_net_535) );
in01f02 g57225_u0 ( .a(FE_OFN2189_n_8567), .o(g57225_sb) );
in01m02 TIMEBOOST_cell_45916 ( .a(TIMEBOOST_net_13876), .o(TIMEBOOST_net_13877) );
in01f02 g57226_u0 ( .a(FE_OFN1397_n_8567), .o(g57226_sb) );
na03m06 TIMEBOOST_cell_67165 ( .a(FE_OFN682_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q), .c(n_3792), .o(TIMEBOOST_net_14292) );
na02m01 TIMEBOOST_cell_4436 ( .a(g52478_da), .b(FE_OFN8_n_11877), .o(TIMEBOOST_net_778) );
in01f02 g57227_u0 ( .a(FE_OFN1387_n_8567), .o(g57227_sb) );
na02f02 TIMEBOOST_cell_4437 ( .a(n_10157), .b(TIMEBOOST_net_778), .o(n_11855) );
na02m01 TIMEBOOST_cell_4438 ( .a(g52477_da), .b(FE_OFN8_n_11877), .o(TIMEBOOST_net_779) );
in01f02 g57228_u0 ( .a(FE_OFN1385_n_8567), .o(g57228_sb) );
na02f02 TIMEBOOST_cell_70980 ( .a(TIMEBOOST_net_20526), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_22698) );
na02f02 TIMEBOOST_cell_4439 ( .a(n_10170), .b(TIMEBOOST_net_779), .o(n_11856) );
na02f02 TIMEBOOST_cell_30741 ( .a(n_9483), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q), .o(TIMEBOOST_net_9475) );
in01f02 g57229_u0 ( .a(FE_OFN2177_n_8567), .o(g57229_sb) );
na02f02 TIMEBOOST_cell_69873 ( .a(TIMEBOOST_net_22144), .b(g64263_sb), .o(n_3910) );
na02f02 TIMEBOOST_cell_26736 ( .a(TIMEBOOST_net_7472), .b(n_8757), .o(g52393_db) );
in01s01 TIMEBOOST_cell_35492 ( .a(TIMEBOOST_net_10083), .o(wbs_dat_i_13_) );
in01f02 g57230_u0 ( .a(FE_OFN2179_n_8567), .o(g57230_sb) );
na02f01 TIMEBOOST_cell_63249 ( .a(TIMEBOOST_net_20571), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_15557) );
na02f02 TIMEBOOST_cell_26738 ( .a(TIMEBOOST_net_7473), .b(n_8757), .o(g52446_db) );
na02m02 TIMEBOOST_cell_68857 ( .a(TIMEBOOST_net_21636), .b(TIMEBOOST_net_20282), .o(TIMEBOOST_net_13245) );
in01f02 g57231_u0 ( .a(FE_OFN1413_n_8567), .o(g57231_sb) );
in01s01 TIMEBOOST_cell_35493 ( .a(TIMEBOOST_net_10084), .o(TIMEBOOST_net_10083) );
na03f04 TIMEBOOST_cell_66441 ( .a(TIMEBOOST_net_17057), .b(n_6287), .c(g62632_sb), .o(n_6289) );
no03f40 TIMEBOOST_cell_64378 ( .a(n_15929), .b(n_15924), .c(n_15324), .o(n_15325) );
in01f02 g57232_u0 ( .a(FE_OFN2174_n_8567), .o(g57232_sb) );
in01s01 TIMEBOOST_cell_35497 ( .a(TIMEBOOST_net_10088), .o(TIMEBOOST_net_10087) );
in01f02 g57233_u0 ( .a(FE_OFN1401_n_8567), .o(g57233_sb) );
na03f02 TIMEBOOST_cell_72904 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q), .b(g64280_sb), .c(g64280_db), .o(TIMEBOOST_net_14950) );
na03f02 TIMEBOOST_cell_73194 ( .a(TIMEBOOST_net_23294), .b(FE_OFN1092_g64577_p), .c(g63574_sb), .o(n_4107) );
in01f02 g57234_u0 ( .a(FE_OFN2178_n_8567), .o(g57234_sb) );
na02m01 TIMEBOOST_cell_68779 ( .a(TIMEBOOST_net_21597), .b(g64752_db), .o(n_3791) );
na02m02 TIMEBOOST_cell_63278 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q), .b(g58396_sb), .o(TIMEBOOST_net_20586) );
in01f02 g57235_u0 ( .a(FE_OFN2174_n_8567), .o(g57235_sb) );
na03s02 TIMEBOOST_cell_70468 ( .a(FE_OFN219_n_9853), .b(FE_OFN526_n_9899), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q), .o(TIMEBOOST_net_22442) );
na02m04 TIMEBOOST_cell_52221 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q), .b(g65845_sb), .o(TIMEBOOST_net_16328) );
na04f04 TIMEBOOST_cell_36876 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q), .b(g58836_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q), .d(FE_OFN2156_n_16439), .o(n_8601) );
in01f02 g57236_u0 ( .a(FE_OFN1377_n_8567), .o(g57236_sb) );
na02s01 TIMEBOOST_cell_47773 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q), .o(TIMEBOOST_net_14104) );
na02s01 TIMEBOOST_cell_52383 ( .a(parchk_pci_ad_out_in_1174), .b(configuration_wb_err_data_577), .o(TIMEBOOST_net_16409) );
na04f04 TIMEBOOST_cell_24281 ( .a(n_9598), .b(g57328_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q), .d(FE_OFN1419_n_8567), .o(n_11421) );
in01f02 g57237_u0 ( .a(FE_OFN1399_n_8567), .o(g57237_sb) );
na04f04 TIMEBOOST_cell_24290 ( .a(n_9615), .b(g57314_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q), .d(FE_OFN1405_n_8567), .o(n_11437) );
na02m04 TIMEBOOST_cell_72093 ( .a(TIMEBOOST_net_23254), .b(FE_OFN1075_n_4740), .o(TIMEBOOST_net_22292) );
in01f02 g57238_u0 ( .a(FE_OFN1396_n_8567), .o(g57238_sb) );
na04f04 TIMEBOOST_cell_36875 ( .a(n_16842), .b(n_16843), .c(n_9328), .d(n_9325), .o(n_12163) );
na03f02 TIMEBOOST_cell_34898 ( .a(TIMEBOOST_net_9375), .b(FE_OFN1413_n_8567), .c(g57441_sb), .o(n_11295) );
na04f02 TIMEBOOST_cell_36878 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q), .b(g54491_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q), .d(n_13617), .o(n_13603) );
in01f02 g57239_u0 ( .a(FE_OFN2169_n_8567), .o(g57239_sb) );
na02s02 TIMEBOOST_cell_30493 ( .a(n_9776), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q), .o(TIMEBOOST_net_9351) );
in01f02 g57240_u0 ( .a(FE_OFN1382_n_8567), .o(g57240_sb) );
in01s01 TIMEBOOST_cell_35494 ( .a(TIMEBOOST_net_10085), .o(wbs_dat_i_26_) );
na03f04 TIMEBOOST_cell_73483 ( .a(wbm_adr_o_31_), .b(g59798_sb), .c(g52405_sb), .o(TIMEBOOST_net_674) );
in01f02 g57241_u0 ( .a(FE_OFN1397_n_8567), .o(g57241_sb) );
na03f02 TIMEBOOST_cell_66285 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q), .b(g62925_sb), .c(g62925_db), .o(n_6031) );
na02s02 TIMEBOOST_cell_43648 ( .a(TIMEBOOST_net_12718), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_11030) );
in01f02 g57242_u0 ( .a(FE_OFN2173_n_8567), .o(g57242_sb) );
na03m06 TIMEBOOST_cell_72430 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q), .b(n_4460), .c(g64813_sb), .o(TIMEBOOST_net_12342) );
na04f02 TIMEBOOST_cell_36877 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q), .b(g54492_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q), .d(n_13617), .o(n_13601) );
na04f02 TIMEBOOST_cell_36880 ( .a(n_829), .b(g54494_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q), .d(n_13617), .o(n_13597) );
in01f02 g57243_u0 ( .a(FE_OFN1408_n_8567), .o(g57243_sb) );
na03s01 TIMEBOOST_cell_72455 ( .a(pci_target_unit_del_sync_bc_in_203), .b(FE_OFN2094_n_2520), .c(g66413_db), .o(n_2521) );
na04m02 TIMEBOOST_cell_73049 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q), .b(FE_OFN2256_n_8060), .c(n_2193), .d(g61730_sb), .o(n_8360) );
in01f02 g57244_u0 ( .a(FE_OFN1420_n_8567), .o(g57244_sb) );
in01s01 TIMEBOOST_cell_35496 ( .a(TIMEBOOST_net_10087), .o(wbs_dat_i_27_) );
na02s01 TIMEBOOST_cell_37611 ( .a(TIMEBOOST_net_10417), .b(g58084_db), .o(n_9711) );
in01f02 g57245_u0 ( .a(FE_OFN2177_n_8567), .o(g57245_sb) );
na03m02 TIMEBOOST_cell_69874 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(FE_OFN1057_n_4727), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q), .o(TIMEBOOST_net_22145) );
na03f04 TIMEBOOST_cell_65933 ( .a(TIMEBOOST_net_17310), .b(FE_OFN1171_n_5592), .c(g62112_sb), .o(n_5585) );
na04f02 TIMEBOOST_cell_36882 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q), .b(g54490_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q), .d(n_13617), .o(n_13605) );
in01f02 g57246_u0 ( .a(FE_OFN1423_n_8567), .o(g57246_sb) );
na03m02 TIMEBOOST_cell_72751 ( .a(n_4442), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q), .c(TIMEBOOST_net_10632), .o(TIMEBOOST_net_17410) );
na03f02 TIMEBOOST_cell_67076 ( .a(FE_OFN1593_n_13741), .b(TIMEBOOST_net_13789), .c(n_13873), .o(n_14408) );
na02f01 TIMEBOOST_cell_54204 ( .a(TIMEBOOST_net_17319), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_15136) );
in01f02 g57247_u0 ( .a(FE_OFN1397_n_8567), .o(g57247_sb) );
na02f02 TIMEBOOST_cell_70421 ( .a(TIMEBOOST_net_22418), .b(FE_OFN1135_g64577_p), .o(n_5388) );
in01f02 g57248_u0 ( .a(FE_OFN1385_n_8567), .o(g57248_sb) );
na02m01 TIMEBOOST_cell_25487 ( .a(g57780_sb), .b(pci_target_unit_fifos_pcir_flush_in), .o(TIMEBOOST_net_6848) );
in01f02 g57249_u0 ( .a(FE_OFN2180_n_8567), .o(g57249_sb) );
na04f02 TIMEBOOST_cell_36881 ( .a(n_971), .b(g54493_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q), .d(n_13617), .o(n_13599) );
in01s01 TIMEBOOST_cell_45976 ( .a(TIMEBOOST_net_13936), .o(TIMEBOOST_net_13937) );
in01f02 g57250_u0 ( .a(FE_OFN1384_n_8567), .o(g57250_sb) );
na02m04 TIMEBOOST_cell_25511 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(g64122_sb), .o(TIMEBOOST_net_6860) );
na02f02 TIMEBOOST_cell_70974 ( .a(TIMEBOOST_net_17576), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_22695) );
in01f02 g57251_u0 ( .a(FE_OFN1376_n_8567), .o(g57251_sb) );
na03s02 TIMEBOOST_cell_65518 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q), .b(g58362_sb), .c(TIMEBOOST_net_11288), .o(TIMEBOOST_net_9525) );
na03f04 TIMEBOOST_cell_67932 ( .a(TIMEBOOST_net_14994), .b(g54134_sb), .c(TIMEBOOST_net_345), .o(n_13671) );
in01f02 g57252_u0 ( .a(FE_OFN1399_n_8567), .o(g57252_sb) );
na03s02 TIMEBOOST_cell_49485 ( .a(g58032_sb), .b(g58032_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q), .o(TIMEBOOST_net_14960) );
in01f02 g57253_u0 ( .a(FE_OFN1387_n_8567), .o(g57253_sb) );
na02f02 TIMEBOOST_cell_50428 ( .a(TIMEBOOST_net_15431), .b(g62760_sb), .o(n_6121) );
na02m02 TIMEBOOST_cell_62595 ( .a(TIMEBOOST_net_20244), .b(FE_OFN1657_n_9502), .o(TIMEBOOST_net_16924) );
na02s02 TIMEBOOST_cell_54177 ( .a(configuration_wb_err_addr_534), .b(TIMEBOOST_net_13839), .o(TIMEBOOST_net_17306) );
in01f02 g57254_u0 ( .a(FE_OFN1374_n_8567), .o(g57254_sb) );
na04s04 TIMEBOOST_cell_34358 ( .a(n_1907), .b(g61745_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q), .d(FE_OFN716_n_8176), .o(n_8327) );
na02m04 TIMEBOOST_cell_68538 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q), .b(n_3747), .o(TIMEBOOST_net_21477) );
na03f02 TIMEBOOST_cell_67352 ( .a(TIMEBOOST_net_16254), .b(g64118_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q), .o(TIMEBOOST_net_15058) );
in01f02 g57255_u0 ( .a(FE_OFN1421_n_8567), .o(g57255_sb) );
na03f02 TIMEBOOST_cell_72888 ( .a(n_1600), .b(g61816_db), .c(g61816_sb), .o(n_8159) );
na03f02 TIMEBOOST_cell_66792 ( .a(TIMEBOOST_net_16780), .b(FE_OFN1315_n_6624), .c(g62535_sb), .o(n_6501) );
in01f02 g57256_u0 ( .a(FE_OFN2177_n_8567), .o(g57256_sb) );
na03m06 TIMEBOOST_cell_64709 ( .a(n_3777), .b(FE_OFN681_n_4460), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q), .o(TIMEBOOST_net_16266) );
in01f02 g57257_u0 ( .a(FE_OFN1412_n_8567), .o(g57257_sb) );
na03m02 TIMEBOOST_cell_72506 ( .a(g64810_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q), .c(TIMEBOOST_net_16147), .o(TIMEBOOST_net_17460) );
na02m02 TIMEBOOST_cell_72156 ( .a(g64258_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q), .o(TIMEBOOST_net_23286) );
na02m02 TIMEBOOST_cell_68323 ( .a(TIMEBOOST_net_21369), .b(g65873_db), .o(TIMEBOOST_net_17010) );
in01f02 g57258_u0 ( .a(FE_OFN2179_n_8567), .o(g57258_sb) );
na03f02 TIMEBOOST_cell_70200 ( .a(TIMEBOOST_net_16638), .b(FE_OFN1150_n_13249), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_393), .o(TIMEBOOST_net_22308) );
na04f04 TIMEBOOST_cell_24589 ( .a(n_9485), .b(g57468_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q), .d(FE_OFN2167_n_8567), .o(n_11264) );
na04f02 TIMEBOOST_cell_36884 ( .a(FE_OCP_RBN2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .b(g54487_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q), .d(n_13617), .o(n_13611) );
in01f02 g57259_u0 ( .a(FE_OFN2187_n_8567), .o(g57259_sb) );
na04f02 TIMEBOOST_cell_36883 ( .a(n_13608), .b(g54488_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q), .d(n_13617), .o(n_13609) );
na04f02 TIMEBOOST_cell_36886 ( .a(n_1225), .b(g54471_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .d(n_13617), .o(n_13619) );
in01f02 g57260_u0 ( .a(FE_OFN1422_n_8567), .o(g57260_sb) );
na04f02 TIMEBOOST_cell_36885 ( .a(n_2269), .b(g54472_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q), .d(n_13617), .o(n_13618) );
na03m04 TIMEBOOST_cell_73144 ( .a(FE_OFN1076_n_4740), .b(TIMEBOOST_net_16352), .c(g64115_sb), .o(n_4045) );
na02m01 TIMEBOOST_cell_31099 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q), .o(TIMEBOOST_net_9654) );
in01f02 g57261_u0 ( .a(FE_OFN1397_n_8567), .o(g57261_sb) );
na03f02 TIMEBOOST_cell_66956 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_16501), .c(FE_OFN1568_n_11027), .o(n_12724) );
na03s04 TIMEBOOST_cell_70102 ( .a(TIMEBOOST_net_17237), .b(FE_OFN1043_n_2037), .c(g65924_sb), .o(TIMEBOOST_net_22259) );
in01f02 g57262_u0 ( .a(FE_OFN1386_n_8567), .o(g57262_sb) );
na03s01 TIMEBOOST_cell_41845 ( .a(g65781_da), .b(g65781_db), .c(TIMEBOOST_net_8289), .o(n_8255) );
in01f02 g57263_u0 ( .a(FE_OFN1374_n_8567), .o(g57263_sb) );
in01s01 TIMEBOOST_cell_67754 ( .a(TIMEBOOST_net_21180), .o(TIMEBOOST_net_21181) );
in01f02 g57264_u0 ( .a(FE_OFN1384_n_8567), .o(g57264_sb) );
na03f02 TIMEBOOST_cell_66796 ( .a(n_4069), .b(g62762_sb), .c(TIMEBOOST_net_7504), .o(n_5470) );
na02m04 TIMEBOOST_cell_68798 ( .a(g64894_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q), .o(TIMEBOOST_net_21607) );
in01f02 g57265_u0 ( .a(FE_OFN1407_n_8567), .o(g57265_sb) );
na04f04 TIMEBOOST_cell_42517 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_775), .c(FE_OFN2136_n_13124), .d(g54339_sb), .o(n_12978) );
na03f02 TIMEBOOST_cell_66287 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q), .b(g63154_sb), .c(g63154_db), .o(n_5833) );
na03f08 TIMEBOOST_cell_41835 ( .a(TIMEBOOST_net_8275), .b(n_5633), .c(g62095_sb), .o(n_5609) );
in01f02 g57266_u0 ( .a(FE_OFN1392_n_8567), .o(g57266_sb) );
na02s01 TIMEBOOST_cell_62594 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q), .o(TIMEBOOST_net_20244) );
na02f02 TIMEBOOST_cell_63953 ( .a(TIMEBOOST_net_20962), .b(FE_OFN1214_n_4151), .o(TIMEBOOST_net_15399) );
na02f02 TIMEBOOST_cell_70057 ( .a(TIMEBOOST_net_22236), .b(g62011_sb), .o(TIMEBOOST_net_20882) );
in01f02 g57267_u0 ( .a(FE_OFN1392_n_8567), .o(g57267_sb) );
na02f02 TIMEBOOST_cell_39455 ( .a(TIMEBOOST_net_11339), .b(g62802_sb), .o(n_5378) );
na04m02 TIMEBOOST_cell_67306 ( .a(TIMEBOOST_net_10398), .b(n_4488), .c(g64975_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q), .o(TIMEBOOST_net_21033) );
in01f02 g57268_u0 ( .a(FE_OFN2170_n_8567), .o(g57268_sb) );
na04f02 TIMEBOOST_cell_36879 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q), .b(g54495_sb), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q), .d(n_13617), .o(n_13595) );
na02m10 TIMEBOOST_cell_45791 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q), .o(TIMEBOOST_net_13790) );
in01f02 g57269_u0 ( .a(FE_OFN1399_n_8567), .o(g57269_sb) );
na02s01 g58434_u3 ( .a(g58434_db), .b(g58434_da), .o(n_9414) );
no02s02 TIMEBOOST_cell_68089 ( .a(TIMEBOOST_net_21252), .b(n_1666), .o(g64630_p) );
in01f02 g57270_u0 ( .a(FE_OFN1396_n_8567), .o(g57270_sb) );
na02m06 TIMEBOOST_cell_68859 ( .a(TIMEBOOST_net_21637), .b(FE_OFN654_n_4508), .o(TIMEBOOST_net_16626) );
na02s01 TIMEBOOST_cell_53221 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_771), .o(TIMEBOOST_net_16828) );
na03m02 TIMEBOOST_cell_72582 ( .a(TIMEBOOST_net_21440), .b(g64797_sb), .c(TIMEBOOST_net_21647), .o(TIMEBOOST_net_17466) );
in01f02 g57271_u0 ( .a(FE_OFN2170_n_8567), .o(g57271_sb) );
in01f02 g57272_u0 ( .a(FE_OFN1382_n_8567), .o(g57272_sb) );
na03f04 TIMEBOOST_cell_46661 ( .a(TIMEBOOST_net_12870), .b(FE_OFN2126_n_16497), .c(g54328_sb), .o(n_12988) );
in01s01 TIMEBOOST_cell_73915 ( .a(TIMEBOOST_net_23479), .o(TIMEBOOST_net_23480) );
in01f02 g57273_u0 ( .a(FE_OFN1399_n_8567), .o(g57273_sb) );
na02s01 g58421_u3 ( .a(g58421_da), .b(g58421_db), .o(n_9426) );
na02s01 TIMEBOOST_cell_48922 ( .a(TIMEBOOST_net_14678), .b(g58435_sb), .o(n_9413) );
na02m01 TIMEBOOST_cell_43025 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q), .o(TIMEBOOST_net_12407) );
in01f02 g57274_u0 ( .a(FE_OFN1420_n_8567), .o(g57274_sb) );
na02m02 TIMEBOOST_cell_47748 ( .a(TIMEBOOST_net_14091), .b(g65689_sb), .o(n_2207) );
na02s01 TIMEBOOST_cell_48325 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q), .b(g58444_sb), .o(TIMEBOOST_net_14380) );
in01f02 g57275_u0 ( .a(FE_OFN1423_n_8567), .o(g57275_sb) );
na02s01 TIMEBOOST_cell_25481 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q), .b(FE_OFN2054_n_8831), .o(TIMEBOOST_net_6845) );
na03f02 TIMEBOOST_cell_70310 ( .a(TIMEBOOST_net_17291), .b(FE_OFN1148_n_13249), .c(n_2103), .o(TIMEBOOST_net_22363) );
na03s02 TIMEBOOST_cell_41917 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q), .b(g58360_sb), .c(g58360_db), .o(n_9463) );
in01f02 g57276_u0 ( .a(FE_OFN1421_n_8567), .o(g57276_sb) );
in01s01 TIMEBOOST_cell_73930 ( .a(wbm_dat_i_16_), .o(TIMEBOOST_net_23495) );
na02f02 TIMEBOOST_cell_71119 ( .a(TIMEBOOST_net_22767), .b(g62761_sb), .o(n_6119) );
in01f02 g57277_u0 ( .a(FE_OFN1404_n_8567), .o(g57277_sb) );
na03f02 TIMEBOOST_cell_66776 ( .a(TIMEBOOST_net_17061), .b(n_6319), .c(g62992_sb), .o(n_5898) );
na02s01 TIMEBOOST_cell_47793 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q), .b(FE_OFN205_n_9140), .o(TIMEBOOST_net_14114) );
na02m02 TIMEBOOST_cell_69014 ( .a(g65340_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q), .o(TIMEBOOST_net_21715) );
in01f02 g57278_u0 ( .a(FE_OFN1425_n_8567), .o(g57278_sb) );
na02s02 TIMEBOOST_cell_48761 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q), .b(g65843_sb), .o(TIMEBOOST_net_14598) );
in01f02 g57279_u0 ( .a(FE_OFN1381_n_8567), .o(g57279_sb) );
no02f02 TIMEBOOST_cell_45227 ( .a(TIMEBOOST_net_7533), .b(FE_RN_545_0), .o(TIMEBOOST_net_13508) );
in01f02 g57280_u0 ( .a(FE_OFN1415_n_8567), .o(g57280_sb) );
na03f02 TIMEBOOST_cell_66539 ( .a(TIMEBOOST_net_16798), .b(FE_OFN1331_n_13547), .c(g53902_sb), .o(n_13539) );
na02m06 TIMEBOOST_cell_68991 ( .a(TIMEBOOST_net_21703), .b(g65320_sb), .o(TIMEBOOST_net_12544) );
in01f02 g57281_u0 ( .a(FE_OFN2169_n_8567), .o(g57281_sb) );
na02f01 TIMEBOOST_cell_43622 ( .a(TIMEBOOST_net_12705), .b(FE_OFN1046_n_16657), .o(TIMEBOOST_net_10958) );
na02s01 TIMEBOOST_cell_37311 ( .a(TIMEBOOST_net_10267), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_8225) );
na03m02 TIMEBOOST_cell_68674 ( .a(n_3741), .b(g64998_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_21545) );
in01f02 g57282_u0 ( .a(FE_OFN1405_n_8567), .o(g57282_sb) );
no02f08 TIMEBOOST_cell_62400 ( .a(n_15998), .b(n_15744), .o(TIMEBOOST_net_20147) );
in01s01 TIMEBOOST_cell_73926 ( .a(wbm_dat_i_14_), .o(TIMEBOOST_net_23491) );
na03m04 TIMEBOOST_cell_73133 ( .a(TIMEBOOST_net_22145), .b(g64257_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q), .o(TIMEBOOST_net_16669) );
in01f02 g57283_u0 ( .a(FE_OFN2182_n_8567), .o(g57283_sb) );
na02s01 TIMEBOOST_cell_27781 ( .a(g57790_sb), .b(TIMEBOOST_net_5307), .o(TIMEBOOST_net_7995) );
na02f02 TIMEBOOST_cell_70571 ( .a(TIMEBOOST_net_22493), .b(g62815_sb), .o(n_5347) );
in01f02 g57284_u0 ( .a(FE_OFN2188_n_8567), .o(g57284_sb) );
na04f10 TIMEBOOST_cell_72407 ( .a(FE_RN_598_0), .b(n_2841), .c(n_385), .d(FE_RN_597_0), .o(FE_RN_601_0) );
na02s01 TIMEBOOST_cell_49217 ( .a(g61879_sb), .b(g61879_db), .o(TIMEBOOST_net_14826) );
na03f02 TIMEBOOST_cell_67662 ( .a(TIMEBOOST_net_17005), .b(FE_OFN1224_n_6391), .c(g62428_sb), .o(n_6743) );
in01f02 g57285_u0 ( .a(FE_OFN1345_n_8567), .o(g57285_sb) );
na02s02 TIMEBOOST_cell_70266 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q), .o(TIMEBOOST_net_22341) );
na02m02 g61981_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61981_db) );
in01f02 g57286_u0 ( .a(FE_OFN1390_n_8567), .o(g57286_sb) );
na03f04 TIMEBOOST_cell_69582 ( .a(n_15262), .b(n_16763), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q), .o(TIMEBOOST_net_21999) );
in01f02 g57287_u0 ( .a(FE_OFN1411_n_8567), .o(g57287_sb) );
na02f02 TIMEBOOST_cell_71377 ( .a(TIMEBOOST_net_22896), .b(g62837_sb), .o(n_7128) );
na02m06 TIMEBOOST_cell_47973 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_143), .o(TIMEBOOST_net_14204) );
na03f02 TIMEBOOST_cell_66541 ( .a(g53924_sb), .b(FE_OFN1326_n_13547), .c(TIMEBOOST_net_16795), .o(n_13468) );
in01f02 g57288_u0 ( .a(FE_OFN1407_n_8567), .o(g57288_sb) );
na03f02 TIMEBOOST_cell_72959 ( .a(TIMEBOOST_net_23209), .b(g64281_sb), .c(FE_OFN1140_g64577_p), .o(TIMEBOOST_net_22467) );
na02m10 TIMEBOOST_cell_54279 ( .a(configuration_pci_err_cs_bit_466), .b(pci_target_unit_wishbone_master_bc_register_reg_3__Q), .o(TIMEBOOST_net_17357) );
in01f02 g57289_u0 ( .a(FE_OFN1368_n_8567), .o(g57289_sb) );
na02f01 TIMEBOOST_cell_49694 ( .a(TIMEBOOST_net_15064), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_13423) );
na02m10 TIMEBOOST_cell_45669 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_13729) );
in01f02 g57290_u0 ( .a(FE_OFN1345_n_8567), .o(g57290_sb) );
na02f02 TIMEBOOST_cell_70829 ( .a(TIMEBOOST_net_22622), .b(g62040_sb), .o(n_7774) );
na03f02 TIMEBOOST_cell_73358 ( .a(parchk_pci_cbe_out_in_1204), .b(FE_OFN1705_n_4868), .c(g52878_sb), .o(TIMEBOOST_net_7996) );
na02m01 g61985_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61985_db) );
in01f02 g57291_u0 ( .a(FE_OFN1422_n_8567), .o(g57291_sb) );
na02m02 TIMEBOOST_cell_72250 ( .a(n_3781), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q), .o(TIMEBOOST_net_23333) );
na03f02 TIMEBOOST_cell_66974 ( .a(FE_OFN1584_n_12306), .b(TIMEBOOST_net_16513), .c(FE_OFN1761_n_10780), .o(n_12504) );
in01f02 g57292_u0 ( .a(FE_OFN1424_n_8567), .o(g57292_sb) );
na02f02 TIMEBOOST_cell_70059 ( .a(TIMEBOOST_net_22237), .b(g61789_sb), .o(n_8223) );
na02m01 TIMEBOOST_cell_62592 ( .a(n_3752), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q), .o(TIMEBOOST_net_20243) );
in01f02 g57293_u0 ( .a(FE_OFN1380_n_8567), .o(g57293_sb) );
na02s01 TIMEBOOST_cell_25311 ( .a(pci_ad_i_29_), .b(parchk_pci_ad_reg_in_1233), .o(TIMEBOOST_net_6760) );
na02s01 TIMEBOOST_cell_53227 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_772), .o(TIMEBOOST_net_16831) );
in01s01 TIMEBOOST_cell_45950 ( .a(TIMEBOOST_net_13910), .o(TIMEBOOST_net_13911) );
in01f02 g57294_u0 ( .a(FE_OFN1383_n_8567), .o(g57294_sb) );
na04f04 TIMEBOOST_cell_24293 ( .a(n_9619), .b(g57310_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q), .d(FE_OFN1425_n_8567), .o(n_11440) );
na03s02 TIMEBOOST_cell_67819 ( .a(TIMEBOOST_net_14050), .b(g65951_db), .c(TIMEBOOST_net_20455), .o(n_7881) );
in01s01 TIMEBOOST_cell_45952 ( .a(TIMEBOOST_net_13913), .o(TIMEBOOST_net_13912) );
in01f02 g57295_u0 ( .a(FE_OFN1414_n_8567), .o(g57295_sb) );
na03f02 TIMEBOOST_cell_72960 ( .a(TIMEBOOST_net_21813), .b(g64270_sb), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_22461) );
in01s01 TIMEBOOST_cell_45951 ( .a(TIMEBOOST_net_13912), .o(TIMEBOOST_net_13901) );
in01f02 g57296_u0 ( .a(FE_OFN1419_n_8567), .o(g57296_sb) );
in01s03 TIMEBOOST_cell_45953 ( .a(pci_target_unit_fifos_pcir_data_in_167), .o(TIMEBOOST_net_13914) );
na02f10 TIMEBOOST_cell_37071 ( .a(TIMEBOOST_net_10147), .b(g54163_da), .o(n_13544) );
in01f02 g57297_u0 ( .a(FE_OFN1415_n_8567), .o(g57297_sb) );
in01f02 g57298_u0 ( .a(FE_OFN1368_n_8567), .o(g57298_sb) );
na02f10 TIMEBOOST_cell_37070 ( .a(n_236), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_10147) );
na02f01 TIMEBOOST_cell_37072 ( .a(n_1381), .b(n_3194), .o(TIMEBOOST_net_10148) );
in01f02 g57299_u0 ( .a(FE_OFN1417_n_8567), .o(g57299_sb) );
na02m02 TIMEBOOST_cell_37441 ( .a(TIMEBOOST_net_10332), .b(g58769_sb), .o(n_9860) );
na02s02 TIMEBOOST_cell_37074 ( .a(wbu_addr_in_273), .b(g58783_sb), .o(TIMEBOOST_net_10149) );
in01f02 g57300_u0 ( .a(FE_OFN1344_n_8567), .o(g57300_sb) );
na02s02 TIMEBOOST_cell_48508 ( .a(TIMEBOOST_net_14471), .b(g57971_sb), .o(TIMEBOOST_net_9423) );
na02m01 g61923_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61923_db) );
in01f02 g57301_u0 ( .a(FE_OFN1390_n_8567), .o(g57301_sb) );
na02s02 g58326_u3 ( .a(g58326_db), .b(g58326_da), .o(n_9488) );
na02f01 TIMEBOOST_cell_37073 ( .a(TIMEBOOST_net_10148), .b(n_3192), .o(TIMEBOOST_net_340) );
na02f01 TIMEBOOST_cell_26799 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_7504) );
in01f02 g57302_u0 ( .a(FE_OFN1401_n_8567), .o(g57302_sb) );
na02s02 TIMEBOOST_cell_37272 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(g65703_sb), .o(TIMEBOOST_net_10248) );
na02s02 TIMEBOOST_cell_37075 ( .a(TIMEBOOST_net_10149), .b(TIMEBOOST_net_5348), .o(n_9841) );
na02s02 TIMEBOOST_cell_48838 ( .a(TIMEBOOST_net_14636), .b(FE_OFN241_n_9830), .o(n_9756) );
in01f02 g57303_u0 ( .a(FE_OFN1416_n_8567), .o(g57303_sb) );
na02s02 TIMEBOOST_cell_63125 ( .a(TIMEBOOST_net_20509), .b(FE_OFN568_n_9528), .o(TIMEBOOST_net_13194) );
na02f02 TIMEBOOST_cell_49310 ( .a(TIMEBOOST_net_14872), .b(g61761_sb), .o(n_8291) );
in01f02 g57304_u0 ( .a(FE_OFN1380_n_8567), .o(g57304_sb) );
na02s03 TIMEBOOST_cell_37077 ( .a(TIMEBOOST_net_10150), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q), .o(n_9116) );
in01s01 TIMEBOOST_cell_45979 ( .a(TIMEBOOST_net_13940), .o(TIMEBOOST_net_13889) );
in01f02 g57305_u0 ( .a(FE_OFN1398_n_8567), .o(g57305_sb) );
na02m10 TIMEBOOST_cell_71964 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q), .b(FE_OFN1643_n_4671), .o(TIMEBOOST_net_23190) );
na02f01 TIMEBOOST_cell_26807 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_7508) );
in01f02 g57306_u0 ( .a(FE_OFN1420_n_8567), .o(g57306_sb) );
na02s01 g58309_u3 ( .a(g58309_da), .b(g58309_db), .o(n_9501) );
in01f02 g57307_u0 ( .a(FE_OFN1425_n_8567), .o(g57307_sb) );
na02m02 TIMEBOOST_cell_37425 ( .a(TIMEBOOST_net_10324), .b(g64138_sb), .o(n_4737) );
in01s01 TIMEBOOST_cell_45990 ( .a(TIMEBOOST_net_13951), .o(TIMEBOOST_net_13950) );
in01f02 g57308_u0 ( .a(FE_OFN1420_n_8567), .o(g57308_sb) );
na02s01 TIMEBOOST_cell_37082 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q), .o(TIMEBOOST_net_10153) );
in01f02 g57309_u0 ( .a(FE_OFN1404_n_8567), .o(g57309_sb) );
na03s02 TIMEBOOST_cell_41651 ( .a(FE_OFN227_n_9841), .b(g57930_sb), .c(g57930_db), .o(n_9879) );
in01s01 TIMEBOOST_cell_45991 ( .a(pci_target_unit_fifos_pcir_data_in_177), .o(TIMEBOOST_net_13952) );
na02s02 TIMEBOOST_cell_48834 ( .a(TIMEBOOST_net_14634), .b(g57995_sb), .o(TIMEBOOST_net_10841) );
in01f02 g57310_u0 ( .a(FE_OFN1425_n_8567), .o(g57310_sb) );
na02m02 TIMEBOOST_cell_54555 ( .a(n_3684), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q), .o(TIMEBOOST_net_17495) );
na03m20 TIMEBOOST_cell_46026 ( .a(n_1724), .b(pci_target_unit_pci_target_sm_rd_from_fifo), .c(n_1615), .o(TIMEBOOST_net_532) );
na02s01 TIMEBOOST_cell_37086 ( .a(TIMEBOOST_net_6755), .b(n_2373), .o(TIMEBOOST_net_10155) );
in01f02 g57311_u0 ( .a(FE_OFN1381_n_8567), .o(g57311_sb) );
na02s03 TIMEBOOST_cell_53229 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_766), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q), .o(TIMEBOOST_net_16832) );
in01f02 g57312_u0 ( .a(FE_OFN1415_n_8567), .o(g57312_sb) );
na02f02 TIMEBOOST_cell_71075 ( .a(TIMEBOOST_net_22745), .b(g62972_sb), .o(n_5938) );
na03f02 TIMEBOOST_cell_66466 ( .a(TIMEBOOST_net_17149), .b(FE_OFN1317_n_6624), .c(g62968_sb), .o(n_5946) );
in01f02 g57313_u0 ( .a(FE_OFN2169_n_8567), .o(g57313_sb) );
na03f02 TIMEBOOST_cell_73602 ( .a(TIMEBOOST_net_17019), .b(FE_OFN1272_n_4096), .c(g62650_sb), .o(n_6246) );
na02f02 TIMEBOOST_cell_37085 ( .a(TIMEBOOST_net_10154), .b(g67057_sb), .o(n_1474) );
na02s01 TIMEBOOST_cell_37088 ( .a(TIMEBOOST_net_6756), .b(n_2373), .o(TIMEBOOST_net_10156) );
in01f02 g57314_u0 ( .a(FE_OFN1405_n_8567), .o(g57314_sb) );
na02m80 TIMEBOOST_cell_72172 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .o(TIMEBOOST_net_23294) );
in01s01 TIMEBOOST_cell_45917 ( .a(TIMEBOOST_net_13927), .o(TIMEBOOST_net_13878) );
in01f02 g57315_u0 ( .a(FE_OFN2182_n_8567), .o(g57315_sb) );
na03f02 TIMEBOOST_cell_66167 ( .a(TIMEBOOST_net_16436), .b(FE_OFN1181_n_3476), .c(g60624_sb), .o(n_4830) );
na02f01 TIMEBOOST_cell_31103 ( .a(n_2705), .b(n_2243), .o(TIMEBOOST_net_9656) );
in01f02 g57316_u0 ( .a(FE_OFN2188_n_8567), .o(g57316_sb) );
na03m02 TIMEBOOST_cell_72497 ( .a(TIMEBOOST_net_21357), .b(n_3755), .c(TIMEBOOST_net_21395), .o(TIMEBOOST_net_17472) );
na03f02 TIMEBOOST_cell_67863 ( .a(TIMEBOOST_net_6915), .b(g52647_sb), .c(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(n_14738) );
na02s01 TIMEBOOST_cell_48835 ( .a(FE_OFN1794_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q), .o(TIMEBOOST_net_14635) );
in01f02 g57317_u0 ( .a(FE_OFN1388_n_8567), .o(g57317_sb) );
na02f02 TIMEBOOST_cell_71076 ( .a(TIMEBOOST_net_17402), .b(FE_OFN1226_n_6391), .o(TIMEBOOST_net_22746) );
na02f02 TIMEBOOST_cell_69971 ( .a(TIMEBOOST_net_22193), .b(g64314_db), .o(n_3861) );
in01f02 g57318_u0 ( .a(FE_OFN1411_n_8567), .o(g57318_sb) );
na02s01 TIMEBOOST_cell_53072 ( .a(TIMEBOOST_net_16753), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_10824) );
na03m02 TIMEBOOST_cell_72979 ( .a(g64954_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q), .c(TIMEBOOST_net_10726), .o(TIMEBOOST_net_20635) );
in01f02 g57319_u0 ( .a(FE_OFN1407_n_8567), .o(g57319_sb) );
na02s01 TIMEBOOST_cell_25337 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_85), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6773) );
na03s02 TIMEBOOST_cell_73026 ( .a(TIMEBOOST_net_7102), .b(FE_OFN775_n_15366), .c(g65893_sb), .o(n_2586) );
na02s01 TIMEBOOST_cell_45559 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q), .o(TIMEBOOST_net_13674) );
in01f02 g57320_u0 ( .a(FE_OFN1389_n_8567), .o(g57320_sb) );
na02m03 TIMEBOOST_cell_68090 ( .a(pci_target_unit_del_sync_sync_req_comp_pending), .b(g66433_sb), .o(TIMEBOOST_net_21253) );
na04f04 TIMEBOOST_cell_65489 ( .a(g61706_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q), .c(FE_OFN714_n_8140), .d(n_2211), .o(n_8415) );
na02s01 TIMEBOOST_cell_45561 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q), .o(TIMEBOOST_net_13675) );
in01f02 g57321_u0 ( .a(FE_OFN1368_n_8567), .o(g57321_sb) );
na02s01 TIMEBOOST_cell_45583 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q), .o(TIMEBOOST_net_13686) );
na02m08 TIMEBOOST_cell_45563 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q), .o(TIMEBOOST_net_13676) );
in01f02 g57322_u0 ( .a(FE_OFN1345_n_8567), .o(g57322_sb) );
na02s01 TIMEBOOST_cell_48339 ( .a(g58432_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q), .o(TIMEBOOST_net_14387) );
na02m01 g61968_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61968_db) );
in01f02 g57323_u0 ( .a(FE_OFN1422_n_8567), .o(g57323_sb) );
na02m02 TIMEBOOST_cell_69163 ( .a(TIMEBOOST_net_21789), .b(g64295_sb), .o(n_3879) );
na02m02 TIMEBOOST_cell_71844 ( .a(TIMEBOOST_net_17204), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q), .o(TIMEBOOST_net_23130) );
na04f04 TIMEBOOST_cell_24095 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q), .b(FE_OFN1349_n_8567), .c(n_9850), .d(g57079_sb), .o(n_11663) );
in01f02 g57324_u0 ( .a(FE_OFN1424_n_8567), .o(g57324_sb) );
na03f02 TIMEBOOST_cell_73771 ( .a(TIMEBOOST_net_16514), .b(FE_OFN1596_n_13741), .c(FE_OCPN1877_n_13903), .o(n_14414) );
na02m10 TIMEBOOST_cell_45565 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q), .o(TIMEBOOST_net_13677) );
na02f02 TIMEBOOST_cell_53119 ( .a(n_2029), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q), .o(TIMEBOOST_net_16777) );
in01f02 g57325_u0 ( .a(FE_OFN1381_n_8567), .o(g57325_sb) );
in01s01 TIMEBOOST_cell_73941 ( .a(TIMEBOOST_net_23505), .o(TIMEBOOST_net_23506) );
na02m10 TIMEBOOST_cell_45567 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q), .o(TIMEBOOST_net_13678) );
na02m02 TIMEBOOST_cell_69629 ( .a(TIMEBOOST_net_22022), .b(TIMEBOOST_net_14837), .o(TIMEBOOST_net_17011) );
in01f02 g57326_u0 ( .a(FE_OFN1383_n_8567), .o(g57326_sb) );
na02s01 TIMEBOOST_cell_45569 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q), .o(TIMEBOOST_net_13679) );
na04f04 TIMEBOOST_cell_24093 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN1349_n_8567), .c(n_9575), .d(g57353_sb), .o(n_11394) );
in01f02 g57327_u0 ( .a(FE_OFN1415_n_8567), .o(g57327_sb) );
na03s02 TIMEBOOST_cell_42120 ( .a(g58187_sb), .b(FE_OFN270_n_9836), .c(g58187_db), .o(n_9598) );
na04f04 TIMEBOOST_cell_24092 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q), .b(FE_OFN1349_n_8567), .c(n_9518), .d(g57421_sb), .o(n_11316) );
na02f01 TIMEBOOST_cell_26821 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .b(FE_OFN1117_g64577_p), .o(TIMEBOOST_net_7515) );
in01f02 g57328_u0 ( .a(FE_OFN1419_n_8567), .o(g57328_sb) );
na02m01 TIMEBOOST_cell_25351 ( .a(n_2967), .b(n_2681), .o(TIMEBOOST_net_6780) );
na02s02 TIMEBOOST_cell_37089 ( .a(TIMEBOOST_net_10156), .b(g67057_sb), .o(n_1640) );
na02s01 TIMEBOOST_cell_37092 ( .a(TIMEBOOST_net_6757), .b(n_2373), .o(TIMEBOOST_net_10158) );
in01f02 g57329_u0 ( .a(FE_OFN1415_n_8567), .o(g57329_sb) );
na02s03 TIMEBOOST_cell_25353 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q), .o(TIMEBOOST_net_6781) );
na03f02 TIMEBOOST_cell_73671 ( .a(TIMEBOOST_net_8332), .b(FE_OFN2106_g64577_p), .c(g63092_sb), .o(n_5068) );
na02s01 TIMEBOOST_cell_37094 ( .a(TIMEBOOST_net_6758), .b(n_2373), .o(TIMEBOOST_net_10159) );
in01f02 g57330_u0 ( .a(FE_OFN1368_n_8567), .o(g57330_sb) );
na02s02 TIMEBOOST_cell_37093 ( .a(TIMEBOOST_net_10158), .b(g67057_sb), .o(n_1652) );
na02s01 TIMEBOOST_cell_37096 ( .a(TIMEBOOST_net_6759), .b(n_2373), .o(TIMEBOOST_net_10160) );
in01f02 g57331_u0 ( .a(FE_OFN1344_n_8567), .o(g57331_sb) );
na02s02 TIMEBOOST_cell_48510 ( .a(TIMEBOOST_net_14472), .b(TIMEBOOST_net_10379), .o(TIMEBOOST_net_9485) );
na02m02 g61972_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61972_db) );
in01f02 g57332_u0 ( .a(FE_OFN1417_n_8567), .o(g57332_sb) );
na02s01 TIMEBOOST_cell_52778 ( .a(TIMEBOOST_net_16606), .b(TIMEBOOST_net_10923), .o(TIMEBOOST_net_9522) );
na02m02 TIMEBOOST_cell_37095 ( .a(TIMEBOOST_net_10159), .b(g67057_sb), .o(n_1614) );
na02f02 TIMEBOOST_cell_26829 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_7519) );
in01f02 g57333_u0 ( .a(FE_OFN1390_n_8567), .o(g57333_sb) );
na02f02 TIMEBOOST_cell_70523 ( .a(TIMEBOOST_net_22469), .b(g62742_sb), .o(n_5495) );
na02m02 TIMEBOOST_cell_37097 ( .a(TIMEBOOST_net_10160), .b(g67057_sb), .o(n_1683) );
in01s01 TIMEBOOST_cell_45997 ( .a(TIMEBOOST_net_13958), .o(TIMEBOOST_net_13857) );
in01f02 g57334_u0 ( .a(FE_OFN1401_n_8567), .o(g57334_sb) );
no02s01 TIMEBOOST_cell_25361 ( .a(n_1780), .b(n_2354), .o(TIMEBOOST_net_6785) );
na03f02 TIMEBOOST_cell_66639 ( .a(TIMEBOOST_net_16788), .b(FE_OFN1813_n_2919), .c(TIMEBOOST_net_15953), .o(n_13334) );
na02s01 TIMEBOOST_cell_37100 ( .a(parchk_pci_ad_reg_in_1213), .b(n_2503), .o(TIMEBOOST_net_10162) );
in01f02 g57335_u0 ( .a(FE_OFN1416_n_8567), .o(g57335_sb) );
na02s01 TIMEBOOST_cell_25363 ( .a(n_1117), .b(pci_target_unit_fifos_pcir_flush_in), .o(TIMEBOOST_net_6786) );
na03f02 TIMEBOOST_cell_66971 ( .a(n_11823), .b(TIMEBOOST_net_16040), .c(n_12099), .o(n_12506) );
na03f06 TIMEBOOST_cell_66871 ( .a(n_12228), .b(FE_OFN1749_n_12004), .c(TIMEBOOST_net_21082), .o(n_12759) );
in01f02 g57336_u0 ( .a(FE_OFN1380_n_8567), .o(g57336_sb) );
na03s02 TIMEBOOST_cell_67663 ( .a(TIMEBOOST_net_14924), .b(g57934_sb), .c(TIMEBOOST_net_16850), .o(TIMEBOOST_net_9571) );
na02s01 TIMEBOOST_cell_37101 ( .a(TIMEBOOST_net_10162), .b(n_2520), .o(TIMEBOOST_net_5393) );
na02f02 TIMEBOOST_cell_70959 ( .a(TIMEBOOST_net_22687), .b(g62685_sb), .o(n_6168) );
in01f02 g57337_u0 ( .a(FE_OFN1370_n_8567), .o(g57337_sb) );
na03m02 TIMEBOOST_cell_64665 ( .a(n_3739), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q), .c(FE_OFN687_n_4417), .o(TIMEBOOST_net_10536) );
na02m02 TIMEBOOST_cell_69771 ( .a(TIMEBOOST_net_22093), .b(TIMEBOOST_net_7027), .o(TIMEBOOST_net_20471) );
na02f02 TIMEBOOST_cell_70517 ( .a(TIMEBOOST_net_22466), .b(g62721_sb), .o(n_5541) );
in01f02 g57338_u0 ( .a(FE_OFN1420_n_8567), .o(g57338_sb) );
na02s01 TIMEBOOST_cell_62968 ( .a(conf_wb_err_addr_in_948), .b(configuration_wb_err_addr_539), .o(TIMEBOOST_net_20431) );
in01s01 TIMEBOOST_cell_45918 ( .a(TIMEBOOST_net_13878), .o(TIMEBOOST_net_13879) );
na02f02 TIMEBOOST_cell_49896 ( .a(TIMEBOOST_net_15165), .b(g63067_sb), .o(n_5116) );
in01f02 g57339_u0 ( .a(FE_OFN1425_n_8567), .o(g57339_sb) );
na02s01 TIMEBOOST_cell_25281 ( .a(pci_ad_i_10_), .b(parchk_pci_ad_reg_in_1214), .o(TIMEBOOST_net_6745) );
na02s01 TIMEBOOST_cell_48217 ( .a(n_3780), .b(g64977_sb), .o(TIMEBOOST_net_14326) );
na02m02 TIMEBOOST_cell_70061 ( .a(TIMEBOOST_net_22238), .b(g61773_sb), .o(n_8262) );
in01f02 g57340_u0 ( .a(FE_OFN1428_n_8567), .o(g57340_sb) );
na02s02 TIMEBOOST_cell_43106 ( .a(TIMEBOOST_net_12447), .b(g57990_sb), .o(TIMEBOOST_net_10423) );
na02f01 TIMEBOOST_cell_26839 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_7524) );
in01f02 g57341_u0 ( .a(FE_OFN2179_n_8567), .o(g57341_sb) );
na03m02 TIMEBOOST_cell_72854 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q), .b(g65403_sb), .c(TIMEBOOST_net_23237), .o(TIMEBOOST_net_17440) );
na02m02 TIMEBOOST_cell_37091 ( .a(TIMEBOOST_net_10157), .b(g67057_sb), .o(n_1654) );
na03f06 TIMEBOOST_cell_37102 ( .a(n_1209), .b(n_1167), .c(n_1080), .o(TIMEBOOST_net_10163) );
in01f02 g57342_u0 ( .a(FE_OFN1423_n_8567), .o(g57342_sb) );
na02s01 TIMEBOOST_cell_25293 ( .a(pci_ad_i_23_), .b(parchk_pci_ad_reg_in_1227), .o(TIMEBOOST_net_6751) );
na02s02 TIMEBOOST_cell_70464 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q), .b(FE_OFN219_n_9853), .o(TIMEBOOST_net_22440) );
na04m02 TIMEBOOST_cell_67337 ( .a(TIMEBOOST_net_20248), .b(FE_OFN651_n_4508), .c(g65426_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q), .o(TIMEBOOST_net_17107) );
in01f02 g57343_u0 ( .a(FE_OFN1376_n_8567), .o(g57343_sb) );
na02s01 TIMEBOOST_cell_25291 ( .a(pci_ad_i_3_), .b(parchk_pci_ad_reg_in_1207), .o(TIMEBOOST_net_6750) );
no02f02 TIMEBOOST_cell_45228 ( .a(TIMEBOOST_net_13508), .b(n_7702), .o(n_13571) );
in01f02 g57344_u0 ( .a(FE_OFN1398_n_8567), .o(g57344_sb) );
na02s01 TIMEBOOST_cell_25289 ( .a(pci_ad_i_20_), .b(parchk_pci_ad_reg_in_1224), .o(TIMEBOOST_net_6749) );
na02m04 TIMEBOOST_cell_72114 ( .a(FE_OFN1049_n_16657), .b(TIMEBOOST_net_17248), .o(TIMEBOOST_net_23265) );
na04m02 TIMEBOOST_cell_67865 ( .a(g64802_sb), .b(FE_OFN666_n_4495), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q), .d(n_4465), .o(n_4466) );
in01f02 g57345_u0 ( .a(FE_OFN2180_n_8567), .o(g57345_sb) );
na02s01 TIMEBOOST_cell_69702 ( .a(TIMEBOOST_net_20327), .b(FE_OFN1041_n_2037), .o(TIMEBOOST_net_22059) );
na02f02 TIMEBOOST_cell_54334 ( .a(TIMEBOOST_net_17384), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_15459) );
na02f01 TIMEBOOST_cell_26843 ( .a(n_504), .b(FE_RN_447_0), .o(TIMEBOOST_net_7526) );
in01f02 g57346_u0 ( .a(FE_OFN1384_n_8567), .o(g57346_sb) );
in01f02 g57347_u0 ( .a(FE_OFN1376_n_8567), .o(g57347_sb) );
na04f04 TIMEBOOST_cell_24094 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q), .b(FE_OFN1349_n_8567), .c(n_9741), .d(g57184_sb), .o(n_11570) );
na03s02 TIMEBOOST_cell_41922 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q), .b(g58287_sb), .c(g58287_db), .o(n_9516) );
in01f02 g57348_u0 ( .a(FE_OFN1399_n_8567), .o(g57348_sb) );
na02m08 TIMEBOOST_cell_52965 ( .a(wishbone_slave_unit_pcim_sm_data_in_656), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q), .o(TIMEBOOST_net_16700) );
na02f02 TIMEBOOST_cell_70508 ( .a(TIMEBOOST_net_8800), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_22462) );
na02m01 TIMEBOOST_cell_54007 ( .a(n_3764), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q), .o(TIMEBOOST_net_17221) );
in01f02 g57349_u0 ( .a(FE_OFN1389_n_8567), .o(g57349_sb) );
na02m02 TIMEBOOST_cell_44983 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_407), .b(FE_OFN2070_n_15978), .o(TIMEBOOST_net_13386) );
in01f02 g57350_u0 ( .a(FE_OFN1374_n_8567), .o(g57350_sb) );
na02s01 TIMEBOOST_cell_25285 ( .a(pci_ad_i_25_), .b(parchk_pci_ad_reg_in_1229), .o(TIMEBOOST_net_6747) );
na02m02 TIMEBOOST_cell_62770 ( .a(n_4677), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q), .o(TIMEBOOST_net_20332) );
in01f02 g57351_u0 ( .a(FE_OFN1421_n_8567), .o(g57351_sb) );
na02m08 TIMEBOOST_cell_52267 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_143), .o(TIMEBOOST_net_16351) );
na02m10 TIMEBOOST_cell_52679 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q), .o(TIMEBOOST_net_16557) );
in01f02 g57352_u0 ( .a(FE_OFN1376_n_8567), .o(g57352_sb) );
na02s01 TIMEBOOST_cell_25287 ( .a(pci_ad_i_2_), .b(parchk_pci_ad_reg_in_1206), .o(TIMEBOOST_net_6748) );
na03m02 TIMEBOOST_cell_69182 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(FE_OFN928_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q), .o(TIMEBOOST_net_21799) );
in01f02 g57353_u0 ( .a(FE_OFN1349_n_8567), .o(g57353_sb) );
na03f06 TIMEBOOST_cell_66767 ( .a(TIMEBOOST_net_16973), .b(FE_OFN1133_g64577_p), .c(g59372_sb), .o(n_7689) );
na02m02 g61973_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61973_db) );
in01f02 g57354_u0 ( .a(FE_OFN2179_n_8567), .o(g57354_sb) );
na04f20 TIMEBOOST_cell_20911 ( .a(FE_RN_508_0), .b(FE_RN_510_0), .c(FE_RN_512_0), .d(FE_RN_514_0), .o(n_16560) );
na02f02 TIMEBOOST_cell_39379 ( .a(TIMEBOOST_net_11301), .b(g63060_sb), .o(n_5130) );
na02s01 TIMEBOOST_cell_43127 ( .a(FE_OFN219_n_9853), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q), .o(TIMEBOOST_net_12458) );
in01f02 g57355_u0 ( .a(FE_OFN1390_n_8567), .o(g57355_sb) );
na03f03 TIMEBOOST_cell_66973 ( .a(n_16397), .b(TIMEBOOST_net_16048), .c(n_16395), .o(n_16398) );
na02f04 TIMEBOOST_cell_44985 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_390), .b(FE_OFN2070_n_15978), .o(TIMEBOOST_net_13387) );
in01f02 g57356_u0 ( .a(FE_OFN2190_n_8567), .o(g57356_sb) );
na02f02 TIMEBOOST_cell_51018 ( .a(TIMEBOOST_net_15726), .b(FE_OFN1100_g64577_p), .o(TIMEBOOST_net_11451) );
na02f04 TIMEBOOST_cell_37103 ( .a(TIMEBOOST_net_10163), .b(n_1207), .o(n_2232) );
no02m01 TIMEBOOST_cell_26857 ( .a(FE_RN_544_0), .b(n_13784), .o(TIMEBOOST_net_7533) );
in01f02 g57357_u0 ( .a(FE_OFN1397_n_8567), .o(g57357_sb) );
na02s01 TIMEBOOST_cell_25313 ( .a(n_15330), .b(n_2092), .o(TIMEBOOST_net_6761) );
na02f01 TIMEBOOST_cell_26845 ( .a(n_13447), .b(FE_RN_420_0), .o(TIMEBOOST_net_7527) );
in01f02 g57358_u0 ( .a(FE_OFN1388_n_8567), .o(g57358_sb) );
na02s01 TIMEBOOST_cell_25369 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q), .o(TIMEBOOST_net_6789) );
na02f02 TIMEBOOST_cell_26844 ( .a(TIMEBOOST_net_7526), .b(FE_RN_450_0), .o(FE_RN_452_0) );
no02f01 TIMEBOOST_cell_26847 ( .a(FE_RN_370_0), .b(n_13784), .o(TIMEBOOST_net_7528) );
in01f02 g57359_u0 ( .a(FE_OFN1374_n_8567), .o(g57359_sb) );
na03f02 TIMEBOOST_cell_73800 ( .a(TIMEBOOST_net_12145), .b(n_13997), .c(FE_OFN1601_n_13995), .o(g53302_p) );
na02f04 TIMEBOOST_cell_26846 ( .a(TIMEBOOST_net_7527), .b(FE_RN_423_0), .o(FE_RN_425_0) );
no02f01 TIMEBOOST_cell_26849 ( .a(FE_RN_376_0), .b(n_13784), .o(TIMEBOOST_net_7529) );
in01f02 g57360_u0 ( .a(FE_OFN1384_n_8567), .o(g57360_sb) );
in01s01 TIMEBOOST_cell_45954 ( .a(TIMEBOOST_net_13914), .o(TIMEBOOST_net_13915) );
na02s01 TIMEBOOST_cell_37604 ( .a(g58146_sb), .b(FE_OFN219_n_9853), .o(TIMEBOOST_net_10414) );
no02f01 TIMEBOOST_cell_26851 ( .a(FE_RN_710_0), .b(n_13784), .o(TIMEBOOST_net_7530) );
in01f02 g57361_u0 ( .a(FE_OFN1406_n_8567), .o(g57361_sb) );
na02s01 TIMEBOOST_cell_25375 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q), .o(TIMEBOOST_net_6792) );
na02s01 TIMEBOOST_cell_37606 ( .a(g58051_sb), .b(FE_OFN223_n_9844), .o(TIMEBOOST_net_10415) );
no02s01 TIMEBOOST_cell_26853 ( .a(FE_RN_373_0), .b(n_13784), .o(TIMEBOOST_net_7531) );
in01f02 g57362_u0 ( .a(FE_OFN1392_n_8567), .o(g57362_sb) );
na02s01 TIMEBOOST_cell_25377 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_6793) );
na02s01 TIMEBOOST_cell_37608 ( .a(g58154_sb), .b(FE_OFN227_n_9841), .o(TIMEBOOST_net_10416) );
no02s01 TIMEBOOST_cell_26855 ( .a(FE_RN_541_0), .b(n_13784), .o(TIMEBOOST_net_7532) );
in01f02 g57363_u0 ( .a(FE_OFN1392_n_8567), .o(g57363_sb) );
na02s01 TIMEBOOST_cell_25379 ( .a(wbs_ack_o), .b(n_16818), .o(TIMEBOOST_net_6794) );
na02s02 TIMEBOOST_cell_37610 ( .a(g58084_sb), .b(FE_OFN227_n_9841), .o(TIMEBOOST_net_10417) );
na02s01 TIMEBOOST_cell_26859 ( .a(FE_OFN606_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q), .o(TIMEBOOST_net_7534) );
in01f02 g57364_u0 ( .a(FE_OFN2170_n_8567), .o(g57364_sb) );
na04m20 TIMEBOOST_cell_67119 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q), .b(pci_target_unit_fifos_pcir_flush_in), .c(g57780_sb), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q), .o(TIMEBOOST_net_15865) );
no02f04 TIMEBOOST_cell_26856 ( .a(TIMEBOOST_net_7532), .b(FE_RN_542_0), .o(TIMEBOOST_net_736) );
in01f02 g57365_u0 ( .a(FE_OFN1399_n_8567), .o(g57365_sb) );
na02m01 TIMEBOOST_cell_53429 ( .a(TIMEBOOST_net_12677), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q), .o(TIMEBOOST_net_16932) );
na03f04 TIMEBOOST_cell_66564 ( .a(TIMEBOOST_net_17108), .b(FE_OFN1314_n_6624), .c(g62600_sb), .o(n_6350) );
in01f02 g57366_u0 ( .a(FE_OFN1396_n_8567), .o(g57366_sb) );
in01s01 TIMEBOOST_cell_46002 ( .a(TIMEBOOST_net_13962), .o(TIMEBOOST_net_13963) );
na02s01 TIMEBOOST_cell_54167 ( .a(FE_OFN258_n_9862), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q), .o(TIMEBOOST_net_17301) );
in01f02 g57367_u0 ( .a(FE_OFN2170_n_8567), .o(g57367_sb) );
na03m06 TIMEBOOST_cell_68344 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q), .b(FE_OFN906_n_4736), .c(TIMEBOOST_net_16572), .o(TIMEBOOST_net_21380) );
na02f02 TIMEBOOST_cell_69973 ( .a(TIMEBOOST_net_22194), .b(g64326_sb), .o(n_3850) );
na02f02 TIMEBOOST_cell_70448 ( .a(TIMEBOOST_net_609), .b(n_16452), .o(TIMEBOOST_net_22432) );
in01f02 g57368_u0 ( .a(FE_OFN1382_n_8567), .o(g57368_sb) );
na02f02 TIMEBOOST_cell_52287 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q), .b(g64349_sb), .o(TIMEBOOST_net_16361) );
na03m02 TIMEBOOST_cell_72852 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q), .b(g65299_sb), .c(TIMEBOOST_net_23238), .o(TIMEBOOST_net_17379) );
in01f02 g57369_u0 ( .a(FE_OFN1399_n_8567), .o(g57369_sb) );
na02s01 TIMEBOOST_cell_47755 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q), .o(TIMEBOOST_net_14095) );
na02s02 TIMEBOOST_cell_49735 ( .a(FE_OFN560_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q), .o(TIMEBOOST_net_15085) );
in01f02 g57370_u0 ( .a(FE_OFN1420_n_8567), .o(g57370_sb) );
na02s01 TIMEBOOST_cell_37104 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_10164) );
na03f02 TIMEBOOST_cell_25013 ( .a(FE_RN_188_0), .b(n_10890), .c(n_12566), .o(n_12828) );
na02f02 TIMEBOOST_cell_54400 ( .a(TIMEBOOST_net_17417), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_15524) );
in01f02 g57371_u0 ( .a(FE_OFN1423_n_8567), .o(g57371_sb) );
na03f02 TIMEBOOST_cell_66543 ( .a(TIMEBOOST_net_16811), .b(FE_OFN1333_n_13547), .c(g53901_sb), .o(n_13540) );
in01f02 g57372_u0 ( .a(FE_OFN1411_n_8567), .o(g57372_sb) );
na02s01 TIMEBOOST_cell_43071 ( .a(FE_OFN599_n_9687), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q), .o(TIMEBOOST_net_12430) );
in01f02 g57373_u0 ( .a(FE_OFN1419_n_8567), .o(g57373_sb) );
na02s01 TIMEBOOST_cell_52899 ( .a(parchk_pci_ad_out_in_1198), .b(configuration_wb_err_data_601), .o(TIMEBOOST_net_16667) );
na02m02 TIMEBOOST_cell_37754 ( .a(FE_OFN689_n_4438), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q), .o(TIMEBOOST_net_10489) );
in01f02 g57374_u0 ( .a(FE_OFN1422_n_8567), .o(g57374_sb) );
na02m01 TIMEBOOST_cell_25395 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q), .o(TIMEBOOST_net_6802) );
na03s02 TIMEBOOST_cell_49131 ( .a(n_1605), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q), .c(FE_OFN701_n_7845), .o(TIMEBOOST_net_14783) );
na02m01 TIMEBOOST_cell_71876 ( .a(n_3755), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q), .o(TIMEBOOST_net_23146) );
in01f02 g57375_u0 ( .a(FE_OFN1381_n_8567), .o(g57375_sb) );
na02m08 TIMEBOOST_cell_25397 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q), .o(TIMEBOOST_net_6803) );
in01f02 g57376_u0 ( .a(FE_OFN1414_n_8567), .o(g57376_sb) );
na02m02 TIMEBOOST_cell_44794 ( .a(TIMEBOOST_net_13291), .b(g60657_sb), .o(n_5664) );
in01f02 g57377_u0 ( .a(FE_OFN2169_n_8567), .o(g57377_sb) );
na04f02 TIMEBOOST_cell_36861 ( .a(g52594_sb), .b(n_10256), .c(TIMEBOOST_net_9584), .d(TIMEBOOST_net_775), .o(n_11876) );
na03f02 TIMEBOOST_cell_66806 ( .a(TIMEBOOST_net_16839), .b(FE_OFN1345_n_8567), .c(g57160_sb), .o(n_11589) );
in01f02 g57378_u0 ( .a(FE_OFN1384_n_8567), .o(g57378_sb) );
na02s01 TIMEBOOST_cell_25401 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_72), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6805) );
na02f02 TIMEBOOST_cell_69537 ( .a(TIMEBOOST_net_21976), .b(TIMEBOOST_net_14453), .o(TIMEBOOST_net_17119) );
in01f02 g57379_u0 ( .a(FE_OFN2185_n_8567), .o(g57379_sb) );
na02m01 TIMEBOOST_cell_54065 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_149), .o(TIMEBOOST_net_17250) );
na03m04 TIMEBOOST_cell_73120 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q), .b(g64262_sb), .c(TIMEBOOST_net_16958), .o(TIMEBOOST_net_14890) );
na02m02 TIMEBOOST_cell_68783 ( .a(TIMEBOOST_net_21599), .b(g64848_sb), .o(TIMEBOOST_net_16208) );
in01f02 g57380_u0 ( .a(FE_OFN1409_n_8567), .o(g57380_sb) );
na04f80 TIMEBOOST_cell_67116 ( .a(wbu_pciif_frame_out_in), .b(g74434_sb), .c(pci_frame_i), .d(parchk_pci_frame_en_in), .o(n_1551) );
in01f02 g57381_u0 ( .a(FE_OFN1383_n_8567), .o(g57381_sb) );
na02s01 TIMEBOOST_cell_25405 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_74), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6807) );
na03f02 TIMEBOOST_cell_73359 ( .a(parchk_pci_cbe_out_in), .b(FE_OFN1705_n_4868), .c(g52876_sb), .o(TIMEBOOST_net_7999) );
in01f02 g57382_u0 ( .a(FE_OFN1390_n_8567), .o(g57382_sb) );
na02s01 TIMEBOOST_cell_25407 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_77), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6808) );
na02f02 TIMEBOOST_cell_50632 ( .a(TIMEBOOST_net_15533), .b(g62951_sb), .o(n_5979) );
na02f02 TIMEBOOST_cell_50888 ( .a(TIMEBOOST_net_15661), .b(n_8529), .o(n_8531) );
in01f02 g57383_u0 ( .a(FE_OFN1411_n_8567), .o(g57383_sb) );
na03f06 TIMEBOOST_cell_72622 ( .a(FE_OFN1010_n_4734), .b(TIMEBOOST_net_20257), .c(g64155_sb), .o(n_4010) );
na03m02 TIMEBOOST_cell_65398 ( .a(wbs_sel_i_1_), .b(g63584_sb), .c(g63585_db), .o(n_4103) );
na02f02 TIMEBOOST_cell_50526 ( .a(TIMEBOOST_net_15480), .b(g62471_sb), .o(n_6649) );
in01f02 g57384_u0 ( .a(FE_OFN1419_n_8567), .o(g57384_sb) );
na02s01 TIMEBOOST_cell_25411 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q), .o(TIMEBOOST_net_6810) );
na02m02 TIMEBOOST_cell_37774 ( .a(g57940_sb), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_10499) );
na02m02 TIMEBOOST_cell_54082 ( .a(TIMEBOOST_net_17258), .b(FE_OFN1037_n_4732), .o(TIMEBOOST_net_14747) );
in01f02 g57385_u0 ( .a(FE_OFN1392_n_8567), .o(g57385_sb) );
na02s01 TIMEBOOST_cell_25413 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q), .o(TIMEBOOST_net_6811) );
na03f02 TIMEBOOST_cell_67046 ( .a(FE_OFN1606_n_13997), .b(TIMEBOOST_net_16537), .c(FE_OFN1599_n_13995), .o(n_16225) );
na03m02 TIMEBOOST_cell_73134 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(g64106_sb), .c(g64106_db), .o(n_4051) );
in01f02 g57386_u0 ( .a(FE_OFN1406_n_8567), .o(g57386_sb) );
na03s02 TIMEBOOST_cell_72545 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q), .b(FE_OFN587_n_9692), .c(TIMEBOOST_net_23165), .o(TIMEBOOST_net_14923) );
in01f02 g57387_u0 ( .a(FE_OFN2191_n_8567), .o(g57387_sb) );
na03m02 TIMEBOOST_cell_68358 ( .a(TIMEBOOST_net_20183), .b(FE_OFN905_n_4736), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q), .o(TIMEBOOST_net_21387) );
in01f02 g57388_u0 ( .a(FE_OFN1424_n_8567), .o(g57388_sb) );
na02m01 TIMEBOOST_cell_69578 ( .a(TIMEBOOST_net_14203), .b(FE_OFN952_n_2055), .o(TIMEBOOST_net_21997) );
na02f01 TIMEBOOST_cell_70572 ( .a(TIMEBOOST_net_13103), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_22494) );
in01f02 g57389_u0 ( .a(FE_OFN1381_n_8567), .o(g57389_sb) );
na03f02 TIMEBOOST_cell_42213 ( .a(n_4072), .b(g62811_sb), .c(g62811_db), .o(n_5356) );
na02m10 TIMEBOOST_cell_69612 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q), .o(TIMEBOOST_net_22014) );
na02s01 TIMEBOOST_cell_38182 ( .a(g58335_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q), .o(TIMEBOOST_net_10703) );
in01f02 g57390_u0 ( .a(FE_OFN1414_n_8567), .o(g57390_sb) );
na02f02 TIMEBOOST_cell_51184 ( .a(TIMEBOOST_net_15809), .b(g62887_sb), .o(n_6103) );
in01f02 g57391_u0 ( .a(FE_OFN1414_n_8567), .o(g57391_sb) );
na03m02 TIMEBOOST_cell_64600 ( .a(FE_OFN624_n_4409), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q), .c(n_3755), .o(TIMEBOOST_net_10397) );
na02s02 TIMEBOOST_cell_38183 ( .a(TIMEBOOST_net_10703), .b(g58335_db), .o(n_9021) );
na03f02 TIMEBOOST_cell_66998 ( .a(FE_OCPN1877_n_13903), .b(TIMEBOOST_net_16516), .c(FE_OCP_RBN1962_FE_OFN1591_n_13741), .o(n_14298) );
in01f02 g57392_u0 ( .a(FE_OFN1406_n_8567), .o(g57392_sb) );
na02s01 TIMEBOOST_cell_25425 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_6817) );
na02m02 TIMEBOOST_cell_38186 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q), .b(g65288_sb), .o(TIMEBOOST_net_10705) );
na02s01 TIMEBOOST_cell_37106 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_10165) );
in01f02 g57393_u0 ( .a(FE_OFN1404_n_8567), .o(g57393_sb) );
na02s02 TIMEBOOST_cell_68266 ( .a(g65698_sb), .b(TIMEBOOST_net_21139), .o(TIMEBOOST_net_21341) );
na03m02 TIMEBOOST_cell_72659 ( .a(g65309_da), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q), .c(TIMEBOOST_net_12439), .o(TIMEBOOST_net_17463) );
in01f02 g57394_u0 ( .a(FE_OFN1368_n_8567), .o(g57394_sb) );
na02s01 TIMEBOOST_cell_37107 ( .a(TIMEBOOST_net_10165), .b(g61943_sb), .o(TIMEBOOST_net_576) );
na02s02 TIMEBOOST_cell_48512 ( .a(TIMEBOOST_net_14473), .b(TIMEBOOST_net_10381), .o(TIMEBOOST_net_9575) );
na02f01 TIMEBOOST_cell_26989 ( .a(configuration_pci_err_addr_496), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_7599) );
in01f02 g57395_u0 ( .a(FE_OFN1344_n_8567), .o(g57395_sb) );
na02m02 TIMEBOOST_cell_43380 ( .a(g58313_db), .b(TIMEBOOST_net_12584), .o(n_9499) );
na02s01 TIMEBOOST_cell_4160 ( .a(n_9175), .b(n_1304), .o(TIMEBOOST_net_640) );
in01f02 g57396_u0 ( .a(FE_OFN1417_n_8567), .o(g57396_sb) );
na02s01 TIMEBOOST_cell_25427 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_6818) );
na02s01 TIMEBOOST_cell_48017 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_14226) );
in01f02 g57397_u0 ( .a(FE_OFN1390_n_8567), .o(g57397_sb) );
na02f02 TIMEBOOST_cell_70931 ( .a(TIMEBOOST_net_22673), .b(g62933_sb), .o(n_6015) );
na02s01 TIMEBOOST_cell_48019 ( .a(pci_target_unit_fifos_pciw_addr_data_in_142), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q), .o(TIMEBOOST_net_14227) );
na02m02 TIMEBOOST_cell_51917 ( .a(FE_OFN1632_n_9531), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q), .o(TIMEBOOST_net_16176) );
in01f02 g57398_u0 ( .a(FE_OFN1401_n_8567), .o(g57398_sb) );
na02s01 TIMEBOOST_cell_25429 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_6819) );
na02s02 TIMEBOOST_cell_48021 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q), .o(TIMEBOOST_net_14228) );
na02m01 TIMEBOOST_cell_51918 ( .a(TIMEBOOST_net_16176), .b(FE_OFN237_n_9118), .o(TIMEBOOST_net_12736) );
in01f02 g57399_u0 ( .a(FE_OFN1405_n_8567), .o(g57399_sb) );
na03m02 TIMEBOOST_cell_73040 ( .a(n_1893), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q), .c(FE_OFN707_n_8119), .o(TIMEBOOST_net_14796) );
na02m08 TIMEBOOST_cell_48023 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_125), .o(TIMEBOOST_net_14229) );
in01f02 g57400_u0 ( .a(FE_OFN1413_n_8567), .o(g57400_sb) );
na02f08 TIMEBOOST_cell_25431 ( .a(n_2427), .b(n_2237), .o(TIMEBOOST_net_6820) );
na02m01 TIMEBOOST_cell_48025 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q), .o(TIMEBOOST_net_14230) );
na03m04 TIMEBOOST_cell_72710 ( .a(g64817_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q), .c(TIMEBOOST_net_16205), .o(TIMEBOOST_net_17530) );
in01f02 g57401_u0 ( .a(FE_OFN1380_n_8567), .o(g57401_sb) );
na02s02 TIMEBOOST_cell_48027 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_14231) );
in01f02 g57402_u0 ( .a(FE_OFN2173_n_8567), .o(g57402_sb) );
na04m02 TIMEBOOST_cell_67328 ( .a(g64815_sb), .b(n_3774), .c(g64815_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q), .o(TIMEBOOST_net_17459) );
na02f04 TIMEBOOST_cell_50714 ( .a(TIMEBOOST_net_15574), .b(g54185_sb), .o(TIMEBOOST_net_13390) );
na02s02 TIMEBOOST_cell_70465 ( .a(TIMEBOOST_net_22440), .b(FE_OFN579_n_9531), .o(TIMEBOOST_net_20933) );
in01f02 g57403_u0 ( .a(FE_OFN1422_n_8567), .o(g57403_sb) );
na02s01 TIMEBOOST_cell_25435 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_91), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6822) );
na02m02 TIMEBOOST_cell_37775 ( .a(TIMEBOOST_net_10499), .b(g57940_db), .o(n_9130) );
na03f02 TIMEBOOST_cell_66370 ( .a(TIMEBOOST_net_13239), .b(FE_OFN1224_n_6391), .c(g62552_sb), .o(n_6461) );
in01f02 g57404_u0 ( .a(FE_OFN2175_n_8567), .o(g57404_sb) );
na02f01 TIMEBOOST_cell_26093 ( .a(pci_target_unit_pcit_if_strd_addr_in_707), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7151) );
no03f02 TIMEBOOST_cell_73360 ( .a(TIMEBOOST_net_7919), .b(FE_OFN1706_n_4868), .c(FE_RN_211_0), .o(TIMEBOOST_net_10029) );
in01f02 g57405_u0 ( .a(FE_OFN2184_n_8567), .o(g57405_sb) );
na03f02 TIMEBOOST_cell_66443 ( .a(TIMEBOOST_net_21035), .b(FE_OFN1316_n_6624), .c(g62427_sb), .o(n_7386) );
na04m02 TIMEBOOST_cell_46294 ( .a(g64845_sb), .b(FE_OFN1625_n_4438), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q), .d(n_4452), .o(n_4437) );
in01f02 g57406_u0 ( .a(FE_OFN2175_n_8567), .o(g57406_sb) );
na03m02 TIMEBOOST_cell_20799 ( .a(n_13766), .b(configuration_sync_command_bit8), .c(n_7396), .o(TIMEBOOST_net_98) );
na02m02 TIMEBOOST_cell_69122 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q), .b(FE_OFN1663_n_4490), .o(TIMEBOOST_net_21769) );
in01m01 TIMEBOOST_cell_67799 ( .a(TIMEBOOST_net_21226), .o(pci_target_unit_del_sync_sync_req_comp_pending) );
in01f02 g57407_u0 ( .a(FE_OFN1391_n_8567), .o(g57407_sb) );
na02m08 TIMEBOOST_cell_63782 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_), .o(TIMEBOOST_net_20877) );
na02f02 TIMEBOOST_cell_69133 ( .a(TIMEBOOST_net_21774), .b(n_1421), .o(TIMEBOOST_net_20665) );
in01f02 g57408_u0 ( .a(FE_OFN1411_n_8567), .o(g57408_sb) );
na03f02 TIMEBOOST_cell_73536 ( .a(TIMEBOOST_net_17515), .b(FE_OFN1232_n_6391), .c(g62461_sb), .o(n_6674) );
in01f02 g57409_u0 ( .a(FE_OFN1419_n_8567), .o(g57409_sb) );
na03s02 TIMEBOOST_cell_72439 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q), .b(FE_OFN603_n_9687), .c(TIMEBOOST_net_20180), .o(TIMEBOOST_net_14954) );
na02m02 TIMEBOOST_cell_52508 ( .a(TIMEBOOST_net_16471), .b(TIMEBOOST_net_12977), .o(TIMEBOOST_net_9555) );
na04f02 TIMEBOOST_cell_72615 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN1010_n_4734), .c(TIMEBOOST_net_14451), .d(g64154_sb), .o(TIMEBOOST_net_9970) );
in01f02 g57410_u0 ( .a(FE_OFN1422_n_8567), .o(g57410_sb) );
na02m10 TIMEBOOST_cell_71900 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q), .o(TIMEBOOST_net_23158) );
na03f02 TIMEBOOST_cell_70998 ( .a(TIMEBOOST_net_15240), .b(FE_OFN1207_n_6356), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q), .o(TIMEBOOST_net_22707) );
in01f02 g57411_u0 ( .a(FE_OFN1381_n_8567), .o(g57411_sb) );
na02s01 TIMEBOOST_cell_45379 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q), .o(TIMEBOOST_net_13584) );
na02s02 TIMEBOOST_cell_47895 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q), .b(FE_OFN938_n_2292), .o(TIMEBOOST_net_14165) );
in01f02 g57412_u0 ( .a(FE_OFN1414_n_8567), .o(g57412_sb) );
na03f02 TIMEBOOST_cell_66172 ( .a(TIMEBOOST_net_16746), .b(FE_OFN1181_n_3476), .c(g60625_sb), .o(n_4828) );
na02s01 TIMEBOOST_cell_54168 ( .a(TIMEBOOST_net_17301), .b(g57978_sb), .o(TIMEBOOST_net_14958) );
na04f02 TIMEBOOST_cell_67955 ( .a(n_14734), .b(n_14839), .c(TIMEBOOST_net_20562), .d(g52454_sb), .o(n_14836) );
in01f02 g57413_u0 ( .a(FE_OFN2169_n_8567), .o(g57413_sb) );
na02s01 TIMEBOOST_cell_47776 ( .a(TIMEBOOST_net_14105), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_414), .o(n_13167) );
na04f08 TIMEBOOST_cell_73284 ( .a(TIMEBOOST_net_22351), .b(g54161_sb), .c(n_13544), .d(n_692), .o(n_13554) );
na02f02 TIMEBOOST_cell_38246 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(g65709_sb), .o(TIMEBOOST_net_10735) );
in01f02 g57414_u0 ( .a(FE_OFN1384_n_8567), .o(g57414_sb) );
na02m10 TIMEBOOST_cell_52967 ( .a(wishbone_slave_unit_pcim_sm_data_in_657), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q), .o(TIMEBOOST_net_16701) );
na03m02 TIMEBOOST_cell_65399 ( .a(wbs_sel_i_0_), .b(g63584_sb), .c(g63584_db), .o(n_4104) );
na03m02 TIMEBOOST_cell_73152 ( .a(g64127_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q), .c(TIMEBOOST_net_14717), .o(TIMEBOOST_net_20920) );
in01f02 g57415_u0 ( .a(FE_OFN2185_n_8567), .o(g57415_sb) );
na04f04 TIMEBOOST_cell_73186 ( .a(FE_OFN709_n_8232), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q), .c(g61948_sb), .d(TIMEBOOST_net_22360), .o(n_7929) );
na03s01 TIMEBOOST_cell_46333 ( .a(TIMEBOOST_net_12401), .b(FE_OFN229_n_9120), .c(g58184_sb), .o(n_9059) );
na02m02 TIMEBOOST_cell_26987 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_413), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_7598) );
in01f02 g57416_u0 ( .a(FE_OFN1383_n_8567), .o(g57416_sb) );
na03f02 TIMEBOOST_cell_73285 ( .a(TIMEBOOST_net_16414), .b(FE_OFN1138_g64577_p), .c(FE_OFN1135_g64577_p), .o(n_5373) );
na02m02 TIMEBOOST_cell_69699 ( .a(TIMEBOOST_net_22057), .b(TIMEBOOST_net_20331), .o(TIMEBOOST_net_17457) );
in01f02 g57417_u0 ( .a(FE_OFN1409_n_8567), .o(g57417_sb) );
na03f02 TIMEBOOST_cell_72946 ( .a(pci_target_unit_del_sync_addr_in_223), .b(g65237_sb), .c(TIMEBOOST_net_7136), .o(n_2646) );
na03m04 TIMEBOOST_cell_73153 ( .a(g64179_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q), .c(TIMEBOOST_net_14722), .o(TIMEBOOST_net_13088) );
in01f02 g57418_u0 ( .a(FE_OFN1390_n_8567), .o(g57418_sb) );
na02s02 TIMEBOOST_cell_38544 ( .a(FE_OFN221_n_9846), .b(g58209_sb), .o(TIMEBOOST_net_10884) );
na03f02 TIMEBOOST_cell_66440 ( .a(TIMEBOOST_net_17101), .b(FE_OFN1316_n_6624), .c(g62520_sb), .o(n_6536) );
in01f02 g57419_u0 ( .a(FE_OFN1411_n_8567), .o(g57419_sb) );
na03f02 TIMEBOOST_cell_72973 ( .a(TIMEBOOST_net_21916), .b(FE_OFN1056_n_4727), .c(TIMEBOOST_net_23252), .o(TIMEBOOST_net_13095) );
na02s02 TIMEBOOST_cell_38546 ( .a(FE_OFN213_n_9124), .b(g58203_sb), .o(TIMEBOOST_net_10885) );
na02f01 TIMEBOOST_cell_71651 ( .a(TIMEBOOST_net_23033), .b(FE_OFN1579_n_12306), .o(n_12672) );
in01f02 g57420_u0 ( .a(FE_OFN1419_n_8567), .o(g57420_sb) );
na02s02 TIMEBOOST_cell_38548 ( .a(g58197_sb), .b(FE_OFN254_n_9825), .o(TIMEBOOST_net_10886) );
na03f02 TIMEBOOST_cell_34867 ( .a(TIMEBOOST_net_9342), .b(FE_OFN1387_n_8567), .c(g57570_sb), .o(n_11181) );
in01f02 g57421_u0 ( .a(FE_OFN1349_n_8567), .o(g57421_sb) );
na02m06 TIMEBOOST_cell_68663 ( .a(TIMEBOOST_net_21539), .b(g64890_sb), .o(TIMEBOOST_net_12513) );
na03f02 TIMEBOOST_cell_66072 ( .a(n_3204), .b(g63556_sb), .c(TIMEBOOST_net_7657), .o(n_4601) );
in01f02 g57422_u0 ( .a(FE_OFN1404_n_8567), .o(g57422_sb) );
na02s01 TIMEBOOST_cell_48870 ( .a(TIMEBOOST_net_14652), .b(FE_OFN526_n_9899), .o(TIMEBOOST_net_12816) );
na02s02 TIMEBOOST_cell_38550 ( .a(g57945_sb), .b(FE_OFN254_n_9825), .o(TIMEBOOST_net_10887) );
in01s01 TIMEBOOST_cell_67740 ( .a(TIMEBOOST_net_21166), .o(TIMEBOOST_net_21167) );
in01f02 g57423_u0 ( .a(FE_OFN1424_n_8567), .o(g57423_sb) );
na03f10 TIMEBOOST_cell_42529 ( .a(g75072_db), .b(n_16070), .c(g75072_sb), .o(n_16441) );
na02f06 TIMEBOOST_cell_26966 ( .a(TIMEBOOST_net_7587), .b(n_16165), .o(TIMEBOOST_net_421) );
in01s01 TIMEBOOST_cell_73874 ( .a(n_8105), .o(TIMEBOOST_net_23439) );
in01f02 g57424_u0 ( .a(FE_OFN1424_n_8567), .o(g57424_sb) );
na02m01 TIMEBOOST_cell_62590 ( .a(n_3755), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q), .o(TIMEBOOST_net_20242) );
na02m02 TIMEBOOST_cell_69050 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q), .b(FE_OFN1642_n_4671), .o(TIMEBOOST_net_21733) );
in01f02 g57425_u0 ( .a(FE_OFN1381_n_8567), .o(g57425_sb) );
na02f02 TIMEBOOST_cell_71487 ( .a(TIMEBOOST_net_22951), .b(g52402_db), .o(TIMEBOOST_net_20663) );
in01f02 g57426_u0 ( .a(FE_OFN2191_n_8567), .o(g57426_sb) );
na03f02 TIMEBOOST_cell_66641 ( .a(TIMEBOOST_net_8542), .b(FE_OCPN1847_n_14981), .c(g59118_sb), .o(n_8694) );
na02f20 TIMEBOOST_cell_53477 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_384), .o(TIMEBOOST_net_16956) );
na02s02 TIMEBOOST_cell_49276 ( .a(TIMEBOOST_net_14855), .b(TIMEBOOST_net_10852), .o(TIMEBOOST_net_9444) );
in01f02 g57427_u0 ( .a(FE_OFN1414_n_8567), .o(g57427_sb) );
na02s01 TIMEBOOST_cell_45381 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q), .o(TIMEBOOST_net_13585) );
na04f06 TIMEBOOST_cell_46041 ( .a(n_1164), .b(n_1073), .c(n_1159), .d(n_1166), .o(n_2231) );
in01f02 g57428_u0 ( .a(FE_OFN1384_n_8567), .o(g57428_sb) );
na04f04 TIMEBOOST_cell_42521 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_784), .c(FE_OFN2135_n_13124), .d(g54348_sb), .o(n_13094) );
in01s01 TIMEBOOST_cell_67768 ( .a(TIMEBOOST_net_21194), .o(TIMEBOOST_net_21195) );
na02m04 TIMEBOOST_cell_54067 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_130), .o(TIMEBOOST_net_17251) );
in01f02 g57429_u0 ( .a(FE_OFN1404_n_8567), .o(g57429_sb) );
in01f02 g57430_u0 ( .a(FE_OFN1368_n_8567), .o(g57430_sb) );
na03f04 TIMEBOOST_cell_46039 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q), .b(n_12595), .c(pci_target_unit_pcit_if_pcir_fifo_data_in_769), .o(TIMEBOOST_net_12850) );
in01f02 g57431_u0 ( .a(FE_OFN1401_n_8567), .o(g57431_sb) );
na02f01 TIMEBOOST_cell_39454 ( .a(TIMEBOOST_net_9309), .b(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_11339) );
na04m02 TIMEBOOST_cell_67224 ( .a(TIMEBOOST_net_14160), .b(FE_OFN667_n_4495), .c(g65091_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q), .o(TIMEBOOST_net_17470) );
in01f02 g57432_u0 ( .a(FE_OFN1417_n_8567), .o(g57432_sb) );
na02m06 TIMEBOOST_cell_68665 ( .a(TIMEBOOST_net_21540), .b(g64880_sb), .o(TIMEBOOST_net_12472) );
na03s01 TIMEBOOST_cell_72564 ( .a(pci_target_unit_del_sync_addr_in_221), .b(g66403_sb), .c(g66408_db), .o(n_2530) );
na02f02 TIMEBOOST_cell_70082 ( .a(g64869_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q), .o(TIMEBOOST_net_22249) );
in01f02 g57433_u0 ( .a(FE_OFN1377_n_8567), .o(g57433_sb) );
na02s01 TIMEBOOST_cell_47521 ( .a(parchk_pci_ad_reg_in_1235), .b(g67050_db), .o(TIMEBOOST_net_13978) );
na03f02 TIMEBOOST_cell_47360 ( .a(FE_OCPN1865_n_12377), .b(TIMEBOOST_net_13674), .c(FE_OFN1755_n_12681), .o(n_12610) );
na04s02 TIMEBOOST_cell_72878 ( .a(TIMEBOOST_net_12483), .b(g65746_sb), .c(g61796_sb), .d(g61796_db), .o(n_8205) );
in01f02 g57434_u0 ( .a(FE_OFN1416_n_8567), .o(g57434_sb) );
na02m01 TIMEBOOST_cell_52289 ( .a(pci_target_unit_pcit_if_strd_addr_in_698), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62), .o(TIMEBOOST_net_16362) );
na02s01 TIMEBOOST_cell_51591 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q), .o(TIMEBOOST_net_16013) );
in01f02 g57435_u0 ( .a(FE_OFN1377_n_8567), .o(g57435_sb) );
na04f04 TIMEBOOST_cell_24841 ( .a(wbs_dat_o_28_), .b(g52523_sb), .c(FE_OFN2241_g52675_p), .d(wbs_wbb3_2_wbb2_dat_o_i_127), .o(n_13697) );
na02f02 TIMEBOOST_cell_39399 ( .a(TIMEBOOST_net_11311), .b(g63133_sb), .o(n_4984) );
na02f02 TIMEBOOST_cell_72309 ( .a(TIMEBOOST_net_23362), .b(g54169_sb), .o(n_13502) );
in01f02 g57436_u0 ( .a(FE_OFN1402_n_8567), .o(g57436_sb) );
na02s01 TIMEBOOST_cell_47522 ( .a(TIMEBOOST_net_13978), .b(g67049_sb), .o(n_1470) );
na02f01 TIMEBOOST_cell_39411 ( .a(TIMEBOOST_net_11317), .b(g62801_sb), .o(n_5380) );
na02m02 TIMEBOOST_cell_68369 ( .a(TIMEBOOST_net_21392), .b(TIMEBOOST_net_16152), .o(TIMEBOOST_net_17473) );
in01f02 g57437_u0 ( .a(FE_OFN1382_n_8567), .o(g57437_sb) );
na03f02 TIMEBOOST_cell_73772 ( .a(TIMEBOOST_net_16515), .b(FE_OCP_RBN1962_FE_OFN1591_n_13741), .c(FE_OCPN1877_n_13903), .o(n_14284) );
na02f02 TIMEBOOST_cell_39413 ( .a(TIMEBOOST_net_11318), .b(g63433_sb), .o(n_4932) );
in01s01 TIMEBOOST_cell_73991 ( .a(TIMEBOOST_net_23555), .o(TIMEBOOST_net_23556) );
in01f02 g57438_u0 ( .a(FE_OFN1403_n_8567), .o(g57438_sb) );
na02m04 TIMEBOOST_cell_68566 ( .a(FE_OFN631_n_4454), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q), .o(TIMEBOOST_net_21491) );
in01f02 g57439_u0 ( .a(FE_OFN2170_n_8567), .o(g57439_sb) );
na03f10 TIMEBOOST_cell_20803 ( .a(n_15757), .b(n_15474), .c(n_16424), .o(n_16425) );
na03m02 TIMEBOOST_cell_69576 ( .a(n_3780), .b(g65051_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q), .o(TIMEBOOST_net_21996) );
na02m02 TIMEBOOST_cell_71077 ( .a(TIMEBOOST_net_22746), .b(g62920_sb), .o(n_6040) );
in01f02 g57440_u0 ( .a(FE_OFN1380_n_8567), .o(g57440_sb) );
na02f01 TIMEBOOST_cell_62827 ( .a(TIMEBOOST_net_20360), .b(FE_OFN1036_n_4732), .o(TIMEBOOST_net_16363) );
na02f02 TIMEBOOST_cell_39419 ( .a(TIMEBOOST_net_11321), .b(g63552_sb), .o(n_4605) );
na02s02 TIMEBOOST_cell_53190 ( .a(TIMEBOOST_net_16812), .b(TIMEBOOST_net_11485), .o(TIMEBOOST_net_9580) );
in01f02 g57441_u0 ( .a(FE_OFN1380_n_8567), .o(g57441_sb) );
na02m02 TIMEBOOST_cell_69413 ( .a(TIMEBOOST_net_21914), .b(TIMEBOOST_net_10725), .o(TIMEBOOST_net_20620) );
na04f04 TIMEBOOST_cell_24097 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q), .b(FE_OFN1349_n_8567), .c(n_9443), .d(g57529_sb), .o(n_11212) );
in01f02 g57442_u0 ( .a(FE_OFN2173_n_8567), .o(g57442_sb) );
na02m04 TIMEBOOST_cell_71980 ( .a(g64917_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q), .o(TIMEBOOST_net_23198) );
na02f02 TIMEBOOST_cell_26993 ( .a(configuration_pci_err_data_506), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_7601) );
in01f02 g57443_u0 ( .a(FE_OFN1422_n_8567), .o(g57443_sb) );
na02s01 TIMEBOOST_cell_47613 ( .a(g54167_db), .b(g54167_sb), .o(TIMEBOOST_net_14024) );
na04f04 TIMEBOOST_cell_24096 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q), .b(FE_OFN1349_n_8567), .c(n_9886), .d(g57044_sb), .o(n_11690) );
na04f04 TIMEBOOST_cell_34734 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q), .b(FE_OFN1373_n_8567), .c(n_9481), .d(g57478_sb), .o(n_11259) );
in01f02 g57444_u0 ( .a(FE_OFN1391_n_8567), .o(g57444_sb) );
in01s01 TIMEBOOST_cell_35495 ( .a(TIMEBOOST_net_10086), .o(TIMEBOOST_net_10085) );
na02f01 TIMEBOOST_cell_26991 ( .a(configuration_pci_err_cs_bit_465), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_7600) );
in01f02 g57445_u0 ( .a(FE_OFN1407_n_8567), .o(g57445_sb) );
no04f04 TIMEBOOST_cell_73361 ( .a(TIMEBOOST_net_7488), .b(FE_RN_584_0), .c(FE_OFN1710_n_4868), .d(FE_RN_577_0), .o(FE_RN_589_0) );
na04f02 TIMEBOOST_cell_73154 ( .a(n_3087), .b(FE_OFN1001_n_15978), .c(n_3391), .d(n_4681), .o(TIMEBOOST_net_9259) );
in01f02 g57446_u0 ( .a(FE_OFN2187_n_8567), .o(g57446_sb) );
na02s02 TIMEBOOST_cell_70886 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q), .o(TIMEBOOST_net_22651) );
na03m02 TIMEBOOST_cell_69134 ( .a(n_3792), .b(g64862_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q), .o(TIMEBOOST_net_21775) );
na02f01 TIMEBOOST_cell_70926 ( .a(TIMEBOOST_net_17383), .b(FE_OFN1208_n_6356), .o(TIMEBOOST_net_22671) );
in01f02 g57447_u0 ( .a(FE_OFN1370_n_8567), .o(g57447_sb) );
na02f02 TIMEBOOST_cell_44785 ( .a(n_3152), .b(FE_OFN1699_n_5751), .o(TIMEBOOST_net_13287) );
na04f04 TIMEBOOST_cell_24098 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q), .b(FE_OFN1349_n_8567), .c(n_9493), .d(g57457_sb), .o(n_11276) );
no04f06 TIMEBOOST_cell_24101 ( .a(FE_RN_154_0), .b(FE_RN_153_0), .c(n_2250), .d(n_3466), .o(n_4699) );
in01f02 g57448_u0 ( .a(FE_OFN1374_n_8567), .o(g57448_sb) );
na02m01 TIMEBOOST_cell_38219 ( .a(TIMEBOOST_net_10721), .b(TIMEBOOST_net_5438), .o(n_3031) );
na02s01 TIMEBOOST_cell_28007 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_8108) );
na02f02 TIMEBOOST_cell_71343 ( .a(TIMEBOOST_net_22879), .b(TIMEBOOST_net_597), .o(TIMEBOOST_net_15802) );
in01f02 g57449_u0 ( .a(FE_OFN2168_n_8567), .o(g57449_sb) );
na03m02 TIMEBOOST_cell_73155 ( .a(TIMEBOOST_net_22148), .b(g64850_sb), .c(TIMEBOOST_net_22271), .o(TIMEBOOST_net_20983) );
na02s01 TIMEBOOST_cell_26999 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_22__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_7604) );
in01f02 g57450_u0 ( .a(FE_OFN2180_n_8567), .o(g57450_sb) );
na02s02 TIMEBOOST_cell_53074 ( .a(TIMEBOOST_net_16754), .b(TIMEBOOST_net_12919), .o(TIMEBOOST_net_9539) );
na02m02 TIMEBOOST_cell_27003 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_23__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_7606) );
in01f01 g57451_u0 ( .a(FE_OFN1394_n_8567), .o(g57451_sb) );
na02m01 TIMEBOOST_cell_27000 ( .a(TIMEBOOST_net_7604), .b(FE_OFN1084_n_13221), .o(TIMEBOOST_net_650) );
no02f06 g74182_u0 ( .a(n_15457), .b(n_15456), .o(n_15458) );
na03s01 TIMEBOOST_cell_72409 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(n_2299), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q), .o(TIMEBOOST_net_14048) );
in01f02 g57452_u0 ( .a(FE_OFN1408_n_8567), .o(g57452_sb) );
in01s04 TIMEBOOST_cell_62386 ( .a(TIMEBOOST_net_20139), .o(FE_OFN532_n_9823) );
na02s01 TIMEBOOST_cell_68146 ( .a(g54219_sb), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q), .o(TIMEBOOST_net_21281) );
in01f02 g57453_u0 ( .a(FE_OFN1374_n_8567), .o(g57453_sb) );
na03f02 TIMEBOOST_cell_73444 ( .a(TIMEBOOST_net_17440), .b(FE_OFN1289_n_4098), .c(g62940_sb), .o(n_6001) );
na03f02 TIMEBOOST_cell_66150 ( .a(TIMEBOOST_net_16725), .b(FE_OFN1184_n_3476), .c(g60648_sb), .o(n_5678) );
in01f02 g57454_u0 ( .a(FE_OFN1386_n_8567), .o(g57454_sb) );
na04f04 TIMEBOOST_cell_73286 ( .a(n_2699), .b(FE_OFN1188_n_5742), .c(wishbone_slave_unit_wishbone_slave_img_hit_0_), .d(g59368_sb), .o(n_7541) );
na03f02 TIMEBOOST_cell_66566 ( .a(TIMEBOOST_net_17098), .b(FE_OFN1315_n_6624), .c(g62612_sb), .o(n_6333) );
in01f02 g57455_u0 ( .a(FE_OFN1391_n_8567), .o(g57455_sb) );
in01m06 TIMEBOOST_cell_45963 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .o(TIMEBOOST_net_13924) );
in01s01 TIMEBOOST_cell_63587 ( .a(TIMEBOOST_net_20767), .o(TIMEBOOST_net_20766) );
na03m02 TIMEBOOST_cell_70370 ( .a(FE_OFN2021_n_4778), .b(TIMEBOOST_net_16652), .c(TIMEBOOST_net_636), .o(TIMEBOOST_net_22393) );
in01f02 g57456_u0 ( .a(FE_OFN1376_n_8567), .o(g57456_sb) );
na02s01 TIMEBOOST_cell_47511 ( .a(parchk_pci_ad_reg_in_1212), .b(g67043_db), .o(TIMEBOOST_net_13973) );
na03f02 TIMEBOOST_cell_65939 ( .a(TIMEBOOST_net_16666), .b(FE_OFN1164_n_5615), .c(g62102_sb), .o(n_5600) );
in01f02 g57457_u0 ( .a(FE_OFN1349_n_8567), .o(g57457_sb) );
na02f06 g75192_u0 ( .a(n_15915), .b(n_16524), .o(n_16565) );
in01f02 g57458_u0 ( .a(FE_OFN1385_n_8567), .o(g57458_sb) );
na03f02 TIMEBOOST_cell_73156 ( .a(TIMEBOOST_net_14736), .b(g65848_sb), .c(TIMEBOOST_net_20405), .o(n_7979) );
na02s03 TIMEBOOST_cell_68476 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q), .b(TIMEBOOST_net_13869), .o(TIMEBOOST_net_21446) );
in01f02 g57459_u0 ( .a(FE_OFN1390_n_8567), .o(g57459_sb) );
na03f02 TIMEBOOST_cell_72894 ( .a(g61732_sb), .b(g61732_db), .c(n_1943), .o(n_8355) );
na03f02 TIMEBOOST_cell_66975 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_16052), .c(FE_OFN1581_n_12306), .o(n_12491) );
in01f02 g57460_u0 ( .a(FE_OFN1400_n_8567), .o(g57460_sb) );
na02m01 TIMEBOOST_cell_68640 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q), .b(FE_OFN666_n_4495), .o(TIMEBOOST_net_21528) );
na04f04 TIMEBOOST_cell_34735 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q), .b(FE_OFN1373_n_8567), .c(n_9433), .d(g57550_sb), .o(n_11194) );
in01f02 g57461_u0 ( .a(FE_OFN2187_n_8567), .o(g57461_sb) );
na03f02 TIMEBOOST_cell_73157 ( .a(TIMEBOOST_net_22157), .b(g64208_sb), .c(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_22554) );
na02m04 TIMEBOOST_cell_27005 ( .a(FE_OFN1000_n_15978), .b(wishbone_slave_unit_del_sync_addr_out_reg_13__Q), .o(TIMEBOOST_net_7607) );
in01f02 g57462_u0 ( .a(FE_OFN1388_n_8567), .o(g57462_sb) );
na03s02 TIMEBOOST_cell_70034 ( .a(n_1668), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q), .c(FE_OFN701_n_7845), .o(TIMEBOOST_net_22225) );
na02f01 TIMEBOOST_cell_70978 ( .a(TIMEBOOST_net_15339), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_22697) );
in01f02 g57463_u0 ( .a(FE_OFN1386_n_8567), .o(g57463_sb) );
na02f01 TIMEBOOST_cell_44002 ( .a(TIMEBOOST_net_12895), .b(FE_OFN1100_g64577_p), .o(TIMEBOOST_net_11301) );
na03m02 TIMEBOOST_cell_72738 ( .a(n_4482), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q), .c(TIMEBOOST_net_12508), .o(TIMEBOOST_net_20522) );
na03f02 TIMEBOOST_cell_34736 ( .a(TIMEBOOST_net_9503), .b(FE_OFN1422_n_8567), .c(g57410_sb), .o(n_11332) );
in01f02 g57464_u0 ( .a(FE_OFN2177_n_8567), .o(g57464_sb) );
na04f04 TIMEBOOST_cell_24953 ( .a(n_16849), .b(n_10163), .c(n_16848), .d(n_9309), .o(n_12159) );
na03f06 TIMEBOOST_cell_66868 ( .a(n_12228), .b(FE_OFN1749_n_12004), .c(TIMEBOOST_net_21085), .o(n_15439) );
na02f01 TIMEBOOST_cell_27007 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_18__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_7608) );
in01f02 g57465_u0 ( .a(FE_OFN1376_n_8567), .o(g57465_sb) );
na02f01 TIMEBOOST_cell_43038 ( .a(TIMEBOOST_net_12413), .b(FE_OFN1010_n_4734), .o(TIMEBOOST_net_10600) );
na04f04 TIMEBOOST_cell_24124 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q), .b(FE_OFN1403_n_8567), .c(n_8555), .d(g58593_sb), .o(n_8904) );
na02s02 TIMEBOOST_cell_48009 ( .a(FE_OFN1649_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q), .o(TIMEBOOST_net_14222) );
in01f02 g57466_u0 ( .a(FE_OFN1413_n_8567), .o(g57466_sb) );
no02s01 TIMEBOOST_cell_45295 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260), .b(FE_RN_237_0), .o(TIMEBOOST_net_13542) );
na03m06 TIMEBOOST_cell_68694 ( .a(g64994_sb), .b(FE_OFN661_n_4392), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q), .o(TIMEBOOST_net_21555) );
in01f02 g57467_u0 ( .a(FE_OFN1396_n_8567), .o(g57467_sb) );
na02f02 TIMEBOOST_cell_70986 ( .a(TIMEBOOST_net_17487), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_22701) );
na02f02 TIMEBOOST_cell_69631 ( .a(TIMEBOOST_net_22023), .b(TIMEBOOST_net_14381), .o(TIMEBOOST_net_17462) );
na04f02 TIMEBOOST_cell_67957 ( .a(conf_wb_err_addr_in_967), .b(g62127_sb), .c(configuration_wb_err_addr_558), .d(FE_OFN1174_n_5592), .o(n_5569) );
in01f02 g57468_u0 ( .a(FE_OFN2175_n_8567), .o(g57468_sb) );
na04f04 TIMEBOOST_cell_24955 ( .a(n_16850), .b(n_16851), .c(n_10564), .d(n_9982), .o(n_12134) );
na02m04 TIMEBOOST_cell_27009 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_27__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_7609) );
in01f02 g57469_u0 ( .a(FE_OFN2177_n_8567), .o(g57469_sb) );
na02m10 TIMEBOOST_cell_52799 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_151), .o(TIMEBOOST_net_16617) );
na02f04 TIMEBOOST_cell_27008 ( .a(TIMEBOOST_net_7608), .b(FE_OFN1085_n_13221), .o(TIMEBOOST_net_649) );
na02f01 TIMEBOOST_cell_27013 ( .a(FE_OFN2072_n_15978), .b(wishbone_slave_unit_del_sync_addr_out_reg_10__Q), .o(TIMEBOOST_net_7611) );
in01f02 g57470_u0 ( .a(FE_OFN1373_n_8567), .o(g57470_sb) );
in01f02 g57471_u0 ( .a(FE_OFN2184_n_8567), .o(g57471_sb) );
na04f04 TIMEBOOST_cell_24849 ( .a(wbs_dat_o_23_), .b(g52518_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_122), .d(FE_OFN2241_g52675_p), .o(n_13705) );
na03s02 TIMEBOOST_cell_67896 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q), .b(g65896_sb), .c(g65896_db), .o(n_1858) );
in01f02 g57472_u0 ( .a(FE_OFN2184_n_8567), .o(g57472_sb) );
na04m08 TIMEBOOST_cell_73078 ( .a(n_3774), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q), .c(FE_OFN1807_n_4501), .d(g64965_sb), .o(n_3655) );
na02m02 TIMEBOOST_cell_71347 ( .a(TIMEBOOST_net_22881), .b(g62025_sb), .o(n_7847) );
in01f02 g57473_u0 ( .a(FE_OFN1409_n_8567), .o(g57473_sb) );
na02s01 g66401_u2 ( .a(parchk_pci_ad_reg_in_1224), .b(FE_OFN2095_n_2520), .o(g66401_db) );
na02s01 TIMEBOOST_cell_71304 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q), .b(FE_OFN600_n_9687), .o(TIMEBOOST_net_22860) );
in01f02 g57474_u0 ( .a(FE_OFN1396_n_8567), .o(g57474_sb) );
na03f10 TIMEBOOST_cell_64280 ( .a(pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77), .b(n_532), .c(FE_OFN2125_n_16497), .o(TIMEBOOST_net_393) );
na02f02 TIMEBOOST_cell_39421 ( .a(TIMEBOOST_net_11322), .b(g63050_sb), .o(n_5151) );
na02f02 TIMEBOOST_cell_44502 ( .a(TIMEBOOST_net_13145), .b(g62792_sb), .o(n_5404) );
in01f02 g57475_u0 ( .a(FE_OFN2167_n_8567), .o(g57475_sb) );
na04f02 TIMEBOOST_cell_24851 ( .a(n_11716), .b(n_10527), .c(n_10859), .d(n_12560), .o(n_12822) );
na02f04 TIMEBOOST_cell_27014 ( .a(TIMEBOOST_net_7611), .b(FE_OFN1084_n_13221), .o(TIMEBOOST_net_658) );
na03f02 TIMEBOOST_cell_66188 ( .a(TIMEBOOST_net_16438), .b(FE_OFN1179_n_3476), .c(g60669_sb), .o(n_5649) );
in01f02 g57476_u0 ( .a(FE_OFN1382_n_8567), .o(g57476_sb) );
na03m04 TIMEBOOST_cell_72612 ( .a(TIMEBOOST_net_21477), .b(FE_OFN1663_n_4490), .c(TIMEBOOST_net_21743), .o(TIMEBOOST_net_17557) );
na02m01 TIMEBOOST_cell_47859 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q), .o(TIMEBOOST_net_14147) );
in01f02 g57477_u0 ( .a(FE_OFN1400_n_8567), .o(g57477_sb) );
in01s01 TIMEBOOST_cell_35498 ( .a(TIMEBOOST_net_10089), .o(wbs_dat_i_30_) );
na03m04 TIMEBOOST_cell_72148 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(FE_OFN1032_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_23282) );
na03m06 TIMEBOOST_cell_69866 ( .a(TIMEBOOST_net_16612), .b(FE_OFN1057_n_4727), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q), .o(TIMEBOOST_net_22141) );
in01f02 g57478_u0 ( .a(FE_OFN1373_n_8567), .o(g57478_sb) );
na03f02 TIMEBOOST_cell_73287 ( .a(wbm_adr_o_29_), .b(g52402_sb), .c(g59096_sb), .o(TIMEBOOST_net_22951) );
in01s01 TIMEBOOST_cell_67753 ( .a(pci_target_unit_fifos_pcir_data_in_179), .o(TIMEBOOST_net_21180) );
na02m06 TIMEBOOST_cell_27025 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_15__Q), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_7617) );
in01f02 g57479_u0 ( .a(FE_OFN1408_n_8567), .o(g57479_sb) );
na02m10 TIMEBOOST_cell_52995 ( .a(wishbone_slave_unit_pcim_sm_data_in_659), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q), .o(TIMEBOOST_net_16715) );
na02m02 TIMEBOOST_cell_39629 ( .a(TIMEBOOST_net_11426), .b(g62829_sb), .o(n_5318) );
na02m02 TIMEBOOST_cell_69633 ( .a(TIMEBOOST_net_22024), .b(g65346_da), .o(TIMEBOOST_net_17003) );
in01f02 g57480_u0 ( .a(FE_OFN1421_n_8567), .o(g57480_sb) );
in01s01 TIMEBOOST_cell_35499 ( .a(TIMEBOOST_net_10090), .o(TIMEBOOST_net_10089) );
in01s01 TIMEBOOST_cell_73875 ( .a(TIMEBOOST_net_23439), .o(TIMEBOOST_net_23440) );
na02m02 TIMEBOOST_cell_69634 ( .a(n_4442), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q), .o(TIMEBOOST_net_22025) );
in01f02 g57481_u0 ( .a(FE_OFN1419_n_8567), .o(g57481_sb) );
na02f01 TIMEBOOST_cell_54210 ( .a(TIMEBOOST_net_17322), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_15142) );
na02s01 TIMEBOOST_cell_47975 ( .a(FE_OFN527_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q), .o(TIMEBOOST_net_14205) );
na02s01 TIMEBOOST_cell_47889 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q), .b(FE_OFN938_n_2292), .o(TIMEBOOST_net_14162) );
in01f02 g57482_u0 ( .a(FE_OFN1422_n_8567), .o(g57482_sb) );
na03f02 TIMEBOOST_cell_73362 ( .a(TIMEBOOST_net_16703), .b(FE_OFN1299_n_5763), .c(g62051_sb), .o(n_7759) );
na02s04 TIMEBOOST_cell_68480 ( .a(g58778_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q), .o(TIMEBOOST_net_21448) );
in01f02 g57483_u0 ( .a(FE_OFN1370_n_8567), .o(g57483_sb) );
na04f04 TIMEBOOST_cell_46537 ( .a(n_2189), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q), .c(FE_OFN713_n_8140), .d(g61729_sb), .o(n_8362) );
na02s01 TIMEBOOST_cell_47993 ( .a(g57902_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q), .o(TIMEBOOST_net_14214) );
in01f02 g57484_u0 ( .a(FE_OFN1415_n_8567), .o(g57484_sb) );
na03f02 TIMEBOOST_cell_73363 ( .a(TIMEBOOST_net_16709), .b(FE_OFN1299_n_5763), .c(g62043_sb), .o(n_7769) );
in01f02 g57485_u0 ( .a(FE_OFN2167_n_8567), .o(g57485_sb) );
na04f04 TIMEBOOST_cell_24853 ( .a(wbs_dat_o_31_), .b(g52527_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_130), .d(FE_OFN1472_g52675_p), .o(n_13694) );
na03f02 TIMEBOOST_cell_34925 ( .a(TIMEBOOST_net_9495), .b(FE_OFN1412_n_8567), .c(g57205_sb), .o(n_10440) );
na02m02 TIMEBOOST_cell_27021 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_29__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_7615) );
in01f02 g57486_u0 ( .a(FE_OFN1405_n_8567), .o(g57486_sb) );
no02f06 TIMEBOOST_cell_48463 ( .a(FE_RN_582_0), .b(FE_RN_578_0), .o(TIMEBOOST_net_14449) );
na02f02 TIMEBOOST_cell_39467 ( .a(TIMEBOOST_net_11345), .b(g62778_sb), .o(n_5435) );
in01f02 g57487_u0 ( .a(FE_OFN2178_n_8567), .o(g57487_sb) );
in01s01 TIMEBOOST_cell_73876 ( .a(n_8044), .o(TIMEBOOST_net_23441) );
na02f02 TIMEBOOST_cell_27020 ( .a(TIMEBOOST_net_7614), .b(FE_OFN1082_n_13221), .o(TIMEBOOST_net_657) );
na02m02 TIMEBOOST_cell_27023 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_26__Q), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_7616) );
in01f02 g57488_u0 ( .a(FE_OFN1408_n_8567), .o(g57488_sb) );
na02f02 TIMEBOOST_cell_39501 ( .a(TIMEBOOST_net_11362), .b(g63063_sb), .o(n_5124) );
na03m04 TIMEBOOST_cell_73145 ( .a(TIMEBOOST_net_17274), .b(FE_OFN1077_n_4740), .c(g64112_sb), .o(n_4046) );
in01f02 g57489_u0 ( .a(FE_OFN1345_n_8567), .o(g57489_sb) );
na02m02 TIMEBOOST_cell_69472 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q), .o(TIMEBOOST_net_21944) );
na03s01 TIMEBOOST_cell_72536 ( .a(g58141_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q), .c(FE_OFN229_n_9120), .o(TIMEBOOST_net_14236) );
na02s01 TIMEBOOST_cell_68772 ( .a(TIMEBOOST_net_17218), .b(FE_OFN951_n_2055), .o(TIMEBOOST_net_21594) );
in01f02 g57490_u0 ( .a(FE_OFN1388_n_8567), .o(g57490_sb) );
na03f03 TIMEBOOST_cell_25115 ( .a(n_16411), .b(n_16410), .c(n_16409), .o(n_16412) );
in01f02 g57491_u0 ( .a(FE_OFN1421_n_8567), .o(g57491_sb) );
in01s02 TIMEBOOST_cell_45919 ( .a(TIMEBOOST_net_13929), .o(TIMEBOOST_net_13880) );
na02m02 TIMEBOOST_cell_70778 ( .a(n_14755), .b(n_14839), .o(TIMEBOOST_net_22597) );
na02f02 TIMEBOOST_cell_70577 ( .a(TIMEBOOST_net_22496), .b(g59379_sb), .o(n_7681) );
in01f02 g57492_u0 ( .a(FE_OFN1406_n_8567), .o(g57492_sb) );
in01s01 TIMEBOOST_cell_73837 ( .a(TIMEBOOST_net_23401), .o(TIMEBOOST_net_23402) );
na02f02 TIMEBOOST_cell_39577 ( .a(TIMEBOOST_net_11400), .b(g63040_sb), .o(n_5170) );
in01f02 g57493_u0 ( .a(FE_OFN1392_n_8567), .o(g57493_sb) );
na02m06 TIMEBOOST_cell_69105 ( .a(TIMEBOOST_net_21760), .b(g65416_sb), .o(TIMEBOOST_net_12546) );
na02f02 TIMEBOOST_cell_39597 ( .a(TIMEBOOST_net_11410), .b(g63022_sb), .o(n_5203) );
in01f02 g57494_u0 ( .a(FE_OFN1407_n_8567), .o(g57494_sb) );
na02s02 TIMEBOOST_cell_70467 ( .a(TIMEBOOST_net_22441), .b(FE_OFN209_n_9126), .o(TIMEBOOST_net_16984) );
na03f02 TIMEBOOST_cell_73499 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q), .b(g62450_sb), .c(g62450_db), .o(n_6697) );
in01f02 g57495_u0 ( .a(FE_OFN1424_n_8567), .o(g57495_sb) );
na02m02 TIMEBOOST_cell_68668 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN685_n_4417), .o(TIMEBOOST_net_21542) );
in01f02 g57496_u0 ( .a(FE_OFN1424_n_8567), .o(g57496_sb) );
na03f02 TIMEBOOST_cell_73681 ( .a(n_10680), .b(FE_RN_484_0), .c(n_9303), .o(n_15590) );
na02s02 TIMEBOOST_cell_44452 ( .a(TIMEBOOST_net_13120), .b(g58291_db), .o(n_9513) );
na03m02 TIMEBOOST_cell_72922 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q), .b(g65880_sb), .c(g65880_db), .o(TIMEBOOST_net_22354) );
in01f02 g57497_u0 ( .a(FE_OFN1413_n_8567), .o(g57497_sb) );
na02s01 TIMEBOOST_cell_68525 ( .a(TIMEBOOST_net_21470), .b(TIMEBOOST_net_14205), .o(TIMEBOOST_net_20561) );
in01f02 g57498_u0 ( .a(FE_OFN1383_n_8567), .o(g57498_sb) );
na03f02 TIMEBOOST_cell_70580 ( .a(n_3853), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q), .c(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_22498) );
in01f02 g57499_u0 ( .a(FE_OFN1414_n_8567), .o(g57499_sb) );
na03f02 TIMEBOOST_cell_70664 ( .a(n_4038), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q), .c(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_22540) );
na02s01 TIMEBOOST_cell_51427 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q), .o(TIMEBOOST_net_15931) );
in01f02 g57500_u0 ( .a(FE_OFN1419_n_8567), .o(g57500_sb) );
na03f02 TIMEBOOST_cell_70074 ( .a(g64973_sb), .b(n_4452), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q), .o(TIMEBOOST_net_22245) );
na04f04 TIMEBOOST_cell_73288 ( .a(n_2698), .b(FE_OFN1188_n_5742), .c(wishbone_slave_unit_wishbone_slave_img_hit_1_), .d(g59369_sb), .o(n_7540) );
in01f02 g57501_u0 ( .a(FE_OFN1415_n_8567), .o(g57501_sb) );
na03f04 TIMEBOOST_cell_66614 ( .a(TIMEBOOST_net_17122), .b(FE_OFN1323_n_6436), .c(g62444_sb), .o(n_6707) );
in01f02 g57502_u0 ( .a(FE_OFN1368_n_8567), .o(g57502_sb) );
na02s02 TIMEBOOST_cell_71157 ( .a(TIMEBOOST_net_22786), .b(FE_OFN554_n_9864), .o(TIMEBOOST_net_21070) );
na03f02 TIMEBOOST_cell_66043 ( .a(TIMEBOOST_net_8810), .b(n_7618), .c(g59808_sb), .o(n_7615) );
na02f04 TIMEBOOST_cell_51428 ( .a(TIMEBOOST_net_15931), .b(FE_OFN1485_n_15534), .o(TIMEBOOST_net_13485) );
in01f02 g57503_u0 ( .a(FE_OFN1401_n_8567), .o(g57503_sb) );
na02m02 TIMEBOOST_cell_62768 ( .a(n_3747), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q), .o(TIMEBOOST_net_20331) );
in01f02 g57504_u0 ( .a(FE_OFN1417_n_8567), .o(g57504_sb) );
na02m01 TIMEBOOST_cell_47969 ( .a(n_3744), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q), .o(TIMEBOOST_net_14202) );
in01f02 g57505_u0 ( .a(FE_OFN2184_n_8567), .o(g57505_sb) );
na03m02 TIMEBOOST_cell_72526 ( .a(TIMEBOOST_net_10317), .b(g64315_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q), .o(TIMEBOOST_net_22033) );
na02s01 TIMEBOOST_cell_27027 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_1__Q), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_7618) );
in01f02 g57506_u0 ( .a(FE_OFN1416_n_8567), .o(g57506_sb) );
na02m01 TIMEBOOST_cell_68926 ( .a(n_4498), .b(n_4396), .o(TIMEBOOST_net_21671) );
na02f02 TIMEBOOST_cell_39835 ( .a(TIMEBOOST_net_11529), .b(g52442_sb), .o(TIMEBOOST_net_6034) );
na03f02 TIMEBOOST_cell_70070 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN716_n_8176), .c(n_2213), .o(TIMEBOOST_net_22243) );
in01f02 g57507_u0 ( .a(FE_OFN1411_n_8567), .o(g57507_sb) );
na02s01 TIMEBOOST_cell_37147 ( .a(TIMEBOOST_net_10185), .b(g58042_sb), .o(TIMEBOOST_net_202) );
na02m02 TIMEBOOST_cell_68986 ( .a(n_3777), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q), .o(TIMEBOOST_net_21701) );
na02m02 TIMEBOOST_cell_70065 ( .a(TIMEBOOST_net_22240), .b(g61766_sb), .o(n_8279) );
in01f02 g57508_u0 ( .a(FE_OFN1402_n_8567), .o(g57508_sb) );
na02s01 TIMEBOOST_cell_37108 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_10166) );
na04f01 TIMEBOOST_cell_72450 ( .a(g57797_sb), .b(FE_OFN276_n_9941), .c(n_276), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_), .o(TIMEBOOST_net_21353) );
in01f02 g57509_u0 ( .a(FE_OFN1400_n_8567), .o(g57509_sb) );
na02f02 TIMEBOOST_cell_39533 ( .a(TIMEBOOST_net_11378), .b(g54316_sb), .o(n_13292) );
in01f02 g57510_u0 ( .a(FE_OFN1403_n_8567), .o(g57510_sb) );
na04f04 TIMEBOOST_cell_25009 ( .a(n_9276), .b(n_10930), .c(n_9277), .d(n_10078), .o(n_12439) );
in01f02 g57511_u0 ( .a(FE_OFN1405_n_8567), .o(g57511_sb) );
na02s01 TIMEBOOST_cell_37109 ( .a(TIMEBOOST_net_10166), .b(g61943_sb), .o(TIMEBOOST_net_577) );
na02m02 TIMEBOOST_cell_52283 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q), .b(g64325_sb), .o(TIMEBOOST_net_16359) );
na02f01 TIMEBOOST_cell_44522 ( .a(TIMEBOOST_net_13155), .b(FE_OFN1127_g64577_p), .o(n_6132) );
in01f02 g57512_u0 ( .a(FE_OFN1380_n_8567), .o(g57512_sb) );
na02f06 TIMEBOOST_cell_37110 ( .a(n_16940), .b(FE_RN_56_0), .o(TIMEBOOST_net_10167) );
na03m02 TIMEBOOST_cell_64823 ( .a(TIMEBOOST_net_16901), .b(FE_OFN908_n_4734), .c(g64185_sb), .o(TIMEBOOST_net_13045) );
in01f02 g57513_u0 ( .a(FE_OFN1409_n_8567), .o(g57513_sb) );
na02s02 TIMEBOOST_cell_70469 ( .a(TIMEBOOST_net_22442), .b(g58016_sb), .o(n_9776) );
na02f02 TIMEBOOST_cell_50606 ( .a(TIMEBOOST_net_15520), .b(g63156_sb), .o(n_5827) );
in01f02 g57514_u0 ( .a(FE_OFN1420_n_8567), .o(g57514_sb) );
na03f02 TIMEBOOST_cell_66045 ( .a(TIMEBOOST_net_20495), .b(n_7618), .c(g59804_sb), .o(n_7620) );
na02m08 TIMEBOOST_cell_52189 ( .a(configuration_wb_err_addr_563), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .o(TIMEBOOST_net_16312) );
in01f02 g57515_u0 ( .a(FE_OFN1425_n_8567), .o(g57515_sb) );
na03f02 TIMEBOOST_cell_68022 ( .a(TIMEBOOST_net_17367), .b(FE_OFN1260_n_4143), .c(g62952_sb), .o(n_5977) );
na02f02 TIMEBOOST_cell_52256 ( .a(TIMEBOOST_net_16345), .b(g64240_sb), .o(n_3932) );
na02f02 TIMEBOOST_cell_50620 ( .a(TIMEBOOST_net_15527), .b(g62615_sb), .o(n_6327) );
in01f02 g57517_u0 ( .a(FE_OFN1407_n_8567), .o(g57517_sb) );
na02s01 TIMEBOOST_cell_62760 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q), .b(TIMEBOOST_net_13829), .o(TIMEBOOST_net_20327) );
na02s02 TIMEBOOST_cell_39711 ( .a(TIMEBOOST_net_11467), .b(g58447_db), .o(n_9198) );
in01f02 g57518_u0 ( .a(FE_OFN2188_n_8567), .o(g57518_sb) );
na04f04 TIMEBOOST_cell_24855 ( .a(wbs_dat_o_18_), .b(g52512_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_117), .d(FE_OFN2243_g52675_p), .o(n_13815) );
na02m02 TIMEBOOST_cell_27029 ( .a(n_526), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_7619) );
in01f02 g57519_u0 ( .a(FE_OFN1370_n_8567), .o(g57519_sb) );
na02f02 TIMEBOOST_cell_70976 ( .a(TIMEBOOST_net_17399), .b(FE_OFN1247_n_4093), .o(TIMEBOOST_net_22696) );
na02m04 TIMEBOOST_cell_72334 ( .a(TIMEBOOST_net_15867), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_), .o(TIMEBOOST_net_23375) );
in01f02 g57520_u0 ( .a(FE_OFN1374_n_8567), .o(g57520_sb) );
na04f02 TIMEBOOST_cell_67867 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(g65804_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q), .d(FE_OFN952_n_2055), .o(n_1906) );
na03s02 TIMEBOOST_cell_72441 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN938_n_2292), .c(TIMEBOOST_net_21205), .o(TIMEBOOST_net_21350) );
in01f02 g57521_u0 ( .a(FE_OFN2168_n_8567), .o(g57521_sb) );
na04f04 TIMEBOOST_cell_24857 ( .a(wbs_dat_o_16_), .b(g52510_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_115), .d(FE_OFN2243_g52675_p), .o(n_13816) );
na02m01 TIMEBOOST_cell_27028 ( .a(TIMEBOOST_net_7618), .b(FE_OFN1082_n_13221), .o(TIMEBOOST_net_646) );
in01f02 g57522_u0 ( .a(FE_OFN2180_n_8567), .o(g57522_sb) );
na03m02 TIMEBOOST_cell_73027 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(FE_OFN1033_n_4732), .c(TIMEBOOST_net_22183), .o(TIMEBOOST_net_12981) );
na03m02 TIMEBOOST_cell_64589 ( .a(n_2199), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q), .c(FE_OFN1812_n_7845), .o(TIMEBOOST_net_15102) );
in01f01 g57523_u0 ( .a(FE_OFN1394_n_8567), .o(g57523_sb) );
na03f02 TIMEBOOST_cell_24139 ( .a(FE_OFN1398_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .c(n_9341), .o(n_9342) );
na02s01 TIMEBOOST_cell_39723 ( .a(TIMEBOOST_net_11473), .b(g58411_db), .o(n_9206) );
na03m02 TIMEBOOST_cell_68364 ( .a(TIMEBOOST_net_20169), .b(FE_OFN905_n_4736), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q), .o(TIMEBOOST_net_21390) );
in01f02 g57524_u0 ( .a(FE_OFN1399_n_8567), .o(g57524_sb) );
na02m04 TIMEBOOST_cell_52260 ( .a(TIMEBOOST_net_16347), .b(g64250_db), .o(n_3923) );
na02s01 TIMEBOOST_cell_39737 ( .a(TIMEBOOST_net_11480), .b(g57894_db), .o(n_9231) );
na03s01 TIMEBOOST_cell_33115 ( .a(FE_OFN235_n_9834), .b(g57997_sb), .c(g57997_db), .o(n_9796) );
in01f02 g57525_u0 ( .a(FE_OFN1374_n_8567), .o(g57525_sb) );
in01s01 TIMEBOOST_cell_73838 ( .a(n_8531), .o(TIMEBOOST_net_23403) );
na02s01 TIMEBOOST_cell_39743 ( .a(TIMEBOOST_net_11483), .b(TIMEBOOST_net_7534), .o(n_9223) );
na03s01 TIMEBOOST_cell_33116 ( .a(FE_OFN221_n_9846), .b(g57989_sb), .c(g57989_db), .o(n_9807) );
in01f02 g57526_u0 ( .a(FE_OFN1388_n_8567), .o(g57526_sb) );
na04s02 TIMEBOOST_cell_67437 ( .a(wbs_dat_i_12_), .b(TIMEBOOST_net_576), .c(g63599_sb), .d(g63599_db), .o(n_7191) );
na02f04 TIMEBOOST_cell_51582 ( .a(TIMEBOOST_net_16008), .b(FE_RN_365_0), .o(FE_RN_366_0) );
na03f02 TIMEBOOST_cell_73158 ( .a(n_4383), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q), .c(FE_OFN1284_n_4097), .o(TIMEBOOST_net_23339) );
in01f02 g57527_u0 ( .a(FE_OFN1391_n_8567), .o(g57527_sb) );
na03f02 TIMEBOOST_cell_24569 ( .a(n_3366), .b(n_3228), .c(n_3428), .o(n_4799) );
na04m08 TIMEBOOST_cell_67828 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q), .b(FE_OFN625_n_4409), .c(g64910_sb), .d(n_4442), .o(n_4402) );
in01f02 g57528_u0 ( .a(FE_OFN2182_n_8567), .o(g57528_sb) );
na03f02 TIMEBOOST_cell_24861 ( .a(FE_RN_140_0), .b(n_10961), .c(n_12580), .o(n_12842) );
na03f02 TIMEBOOST_cell_73215 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_0_), .b(g60407_sb), .c(TIMEBOOST_net_5466), .o(n_4861) );
na02m01 TIMEBOOST_cell_47979 ( .a(n_3792), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q), .o(TIMEBOOST_net_14207) );
in01f02 g57529_u0 ( .a(FE_OFN1349_n_8567), .o(g57529_sb) );
na03f02 TIMEBOOST_cell_47378 ( .a(FE_OFN1579_n_12306), .b(TIMEBOOST_net_13681), .c(FE_OFN1760_n_10780), .o(n_12658) );
na02m02 TIMEBOOST_cell_50616 ( .a(TIMEBOOST_net_15525), .b(g62640_sb), .o(n_6268) );
na03f06 TIMEBOOST_cell_1818 ( .a(n_16511), .b(n_16268), .c(n_15217), .o(FE_RN_302_0) );
in01f02 g57530_u0 ( .a(FE_OFN1385_n_8567), .o(g57530_sb) );
na02m02 TIMEBOOST_cell_53588 ( .a(TIMEBOOST_net_17011), .b(FE_OFN1244_n_4092), .o(TIMEBOOST_net_15498) );
na02m02 TIMEBOOST_cell_51162 ( .a(TIMEBOOST_net_15798), .b(g62674_sb), .o(n_6191) );
na03m02 TIMEBOOST_cell_68362 ( .a(TIMEBOOST_net_20178), .b(FE_OFN905_n_4736), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q), .o(TIMEBOOST_net_21389) );
in01f02 g57531_u0 ( .a(FE_OFN1390_n_8567), .o(g57531_sb) );
in01s01 TIMEBOOST_cell_35515 ( .a(TIMEBOOST_net_10106), .o(TIMEBOOST_net_10105) );
na02s02 TIMEBOOST_cell_47879 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN938_n_2292), .o(TIMEBOOST_net_14157) );
na03m02 TIMEBOOST_cell_33121 ( .a(TIMEBOOST_net_8262), .b(g64302_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q), .o(TIMEBOOST_net_9973) );
in01f02 g57532_u0 ( .a(FE_OFN2187_n_8567), .o(g57532_sb) );
na04f08 TIMEBOOST_cell_67869 ( .a(FE_OFN1797_n_2299), .b(pci_target_unit_fifos_pcir_data_in_163), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q), .d(g65971_sb), .o(n_2153) );
in01f02 g57533_u0 ( .a(FE_OFN1400_n_8567), .o(g57533_sb) );
na02s02 TIMEBOOST_cell_68270 ( .a(TIMEBOOST_net_17196), .b(FE_OFN938_n_2292), .o(TIMEBOOST_net_21343) );
na02s01 TIMEBOOST_cell_39713 ( .a(TIMEBOOST_net_11468), .b(g58415_db), .o(n_9203) );
na02s01 TIMEBOOST_cell_54015 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_135), .o(TIMEBOOST_net_17225) );
in01f02 g57534_u0 ( .a(FE_OFN1388_n_8567), .o(g57534_sb) );
na03f02 TIMEBOOST_cell_72980 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(FE_OFN1055_n_4727), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q), .o(TIMEBOOST_net_23308) );
na02s02 TIMEBOOST_cell_70184 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q), .b(FE_OFN2108_n_2047), .o(TIMEBOOST_net_22300) );
na02m01 TIMEBOOST_cell_52191 ( .a(configuration_wb_err_cs_bit_570), .b(parchk_pci_cbe_out_in_1204), .o(TIMEBOOST_net_16313) );
in01f02 g57535_u0 ( .a(FE_OFN1387_n_8567), .o(g57535_sb) );
na03s02 TIMEBOOST_cell_72947 ( .a(TIMEBOOST_net_14371), .b(g65876_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_22326) );
na02m02 TIMEBOOST_cell_50458 ( .a(TIMEBOOST_net_15446), .b(g62502_sb), .o(n_6578) );
in01f02 g57536_u0 ( .a(FE_OFN2177_n_8567), .o(g57536_sb) );
in01f02 g57537_u0 ( .a(FE_OFN1376_n_8567), .o(g57537_sb) );
na02f02 TIMEBOOST_cell_54378 ( .a(TIMEBOOST_net_17406), .b(FE_OFN1258_n_4143), .o(TIMEBOOST_net_16458) );
in01s01 TIMEBOOST_cell_67755 ( .a(pci_target_unit_fifos_pcir_data_in_165), .o(TIMEBOOST_net_21182) );
in01f02 g57538_u0 ( .a(FE_OFN1412_n_8567), .o(g57538_sb) );
na03f02 TIMEBOOST_cell_72948 ( .a(pci_target_unit_del_sync_addr_in_226), .b(g65223_sb), .c(TIMEBOOST_net_7164), .o(n_2664) );
na02f02 TIMEBOOST_cell_70984 ( .a(TIMEBOOST_net_20620), .b(FE_OFN1247_n_4093), .o(TIMEBOOST_net_22700) );
in01f02 g57539_u0 ( .a(FE_OFN1396_n_8567), .o(g57539_sb) );
na02m02 TIMEBOOST_cell_44534 ( .a(TIMEBOOST_net_13161), .b(g62819_sb), .o(n_5337) );
in01f02 g57540_u0 ( .a(FE_OFN2167_n_8567), .o(g57540_sb) );
na03f02 TIMEBOOST_cell_66873 ( .a(FE_OFN1565_n_12502), .b(TIMEBOOST_net_15989), .c(n_12313), .o(n_12700) );
na03f02 TIMEBOOST_cell_73364 ( .a(TIMEBOOST_net_16713), .b(FE_OFN1301_n_5763), .c(g62063_sb), .o(n_7746) );
in01f02 g57541_u0 ( .a(FE_OFN2177_n_8567), .o(g57541_sb) );
na02f02 TIMEBOOST_cell_70001 ( .a(TIMEBOOST_net_22208), .b(g61821_sb), .o(n_8147) );
in01f02 g57542_u0 ( .a(FE_OFN2175_n_8567), .o(g57542_sb) );
na04f02 TIMEBOOST_cell_24871 ( .a(g54486_sb), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_), .d(n_13617), .o(n_13613) );
na02f02 TIMEBOOST_cell_63445 ( .a(TIMEBOOST_net_20669), .b(n_15529), .o(n_15538) );
in01f02 g57543_u0 ( .a(FE_OFN1391_n_8567), .o(g57543_sb) );
na03m02 TIMEBOOST_cell_73037 ( .a(TIMEBOOST_net_21752), .b(FE_OFN666_n_4495), .c(TIMEBOOST_net_23372), .o(TIMEBOOST_net_20636) );
na03f02 TIMEBOOST_cell_66725 ( .a(TIMEBOOST_net_17570), .b(FE_OFN1284_n_4097), .c(g62900_sb), .o(n_6077) );
na02s02 TIMEBOOST_cell_49284 ( .a(TIMEBOOST_net_14859), .b(TIMEBOOST_net_10880), .o(TIMEBOOST_net_9337) );
in01f02 g57544_u0 ( .a(FE_OFN2185_n_8567), .o(g57544_sb) );
na04f02 TIMEBOOST_cell_24873 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q), .b(g54484_sb), .c(FE_OCP_RBN2265_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .d(n_13617), .o(n_13616) );
na02m04 TIMEBOOST_cell_68993 ( .a(TIMEBOOST_net_21704), .b(g65421_sb), .o(TIMEBOOST_net_10632) );
in01s01 TIMEBOOST_cell_73942 ( .a(wbm_dat_i_21_), .o(TIMEBOOST_net_23507) );
in01f02 g57545_u0 ( .a(FE_OFN1409_n_8567), .o(g57545_sb) );
na03f02 TIMEBOOST_cell_34771 ( .a(TIMEBOOST_net_9364), .b(FE_OFN1387_n_8567), .c(g57579_sb), .o(n_11173) );
na02m01 TIMEBOOST_cell_47957 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q), .o(TIMEBOOST_net_14196) );
na04s02 TIMEBOOST_cell_33127 ( .a(FE_OFN252_n_9868), .b(g58227_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q), .d(g58227_db), .o(TIMEBOOST_net_9582) );
in01f02 g57546_u0 ( .a(FE_OFN1396_n_8567), .o(g57546_sb) );
na03f02 TIMEBOOST_cell_25017 ( .a(n_11013), .b(FE_RN_98_0), .c(n_12591), .o(n_12853) );
in01f02 g57547_u0 ( .a(FE_OFN2167_n_8567), .o(g57547_sb) );
na02s01 TIMEBOOST_cell_44137 ( .a(FE_OFN1648_n_9428), .b(n_15567), .o(TIMEBOOST_net_12963) );
na02m02 TIMEBOOST_cell_63895 ( .a(TIMEBOOST_net_20933), .b(g58383_sb), .o(n_9448) );
na02m10 TIMEBOOST_cell_52969 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q), .b(wishbone_slave_unit_pcim_sm_data_in_635), .o(TIMEBOOST_net_16702) );
in01f02 g57548_u0 ( .a(FE_OFN1382_n_8567), .o(g57548_sb) );
na04s02 TIMEBOOST_cell_72893 ( .a(TIMEBOOST_net_10461), .b(g65725_sb), .c(g61771_sb), .d(g61771_db), .o(n_8267) );
na02f02 TIMEBOOST_cell_70961 ( .a(TIMEBOOST_net_22688), .b(g62930_sb), .o(n_6021) );
na02m02 TIMEBOOST_cell_68557 ( .a(TIMEBOOST_net_21486), .b(g64911_sb), .o(TIMEBOOST_net_12537) );
in01f02 g57549_u0 ( .a(FE_OFN1400_n_8567), .o(g57549_sb) );
na03f02 TIMEBOOST_cell_47245 ( .a(FE_OFN1566_n_12502), .b(TIMEBOOST_net_13525), .c(n_12313), .o(n_12748) );
in01f02 g57550_u0 ( .a(FE_OFN1373_n_8567), .o(g57550_sb) );
na02f01 TIMEBOOST_cell_63859 ( .a(TIMEBOOST_net_20915), .b(FE_OFN877_g64577_p), .o(TIMEBOOST_net_15165) );
na04f04 TIMEBOOST_cell_73773 ( .a(FE_RN_909_0), .b(n_11841), .c(n_16404), .d(FE_RN_910_0), .o(n_16406) );
in01f02 g57551_u0 ( .a(FE_OFN1408_n_8567), .o(g57551_sb) );
na03f02 TIMEBOOST_cell_25019 ( .a(n_10105), .b(FE_RN_191_0), .c(n_12442), .o(n_12775) );
na04m06 TIMEBOOST_cell_72831 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q), .b(FE_OFN1660_n_4490), .c(g64768_sb), .d(n_3780), .o(n_3781) );
na02f01 TIMEBOOST_cell_44536 ( .a(TIMEBOOST_net_13162), .b(g62795_sb), .o(n_5396) );
in01f02 g57552_u0 ( .a(FE_OFN1402_n_8567), .o(g57552_sb) );
na02s02 TIMEBOOST_cell_48768 ( .a(TIMEBOOST_net_14601), .b(TIMEBOOST_net_11289), .o(TIMEBOOST_net_9438) );
na02s02 TIMEBOOST_cell_68263 ( .a(TIMEBOOST_net_21339), .b(g65775_db), .o(n_2192) );
na03f02 TIMEBOOST_cell_73365 ( .a(TIMEBOOST_net_16711), .b(FE_OFN1300_n_5763), .c(g62061_sb), .o(n_7749) );
in01f02 g57553_u0 ( .a(FE_OFN1416_n_8567), .o(g57553_sb) );
na03f02 TIMEBOOST_cell_25021 ( .a(FE_RN_194_0), .b(n_10731), .c(n_12583), .o(n_12845) );
na02m02 TIMEBOOST_cell_48029 ( .a(FE_OFN1654_n_9502), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q), .o(TIMEBOOST_net_14232) );
na02f02 TIMEBOOST_cell_31820 ( .a(TIMEBOOST_net_10014), .b(n_2855), .o(n_4644) );
in01f02 g57554_u0 ( .a(FE_OFN1411_n_8567), .o(g57554_sb) );
na02m10 TIMEBOOST_cell_52997 ( .a(wishbone_slave_unit_pcim_sm_data_in_647), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q), .o(TIMEBOOST_net_16716) );
na03m04 TIMEBOOST_cell_73088 ( .a(g65364_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q), .c(TIMEBOOST_net_20367), .o(TIMEBOOST_net_17050) );
na03f02 TIMEBOOST_cell_73159 ( .a(TIMEBOOST_net_12867), .b(g52626_sb), .c(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_5471) );
in01f02 g57555_u0 ( .a(FE_OFN1402_n_8567), .o(g57555_sb) );
na03f02 TIMEBOOST_cell_73451 ( .a(TIMEBOOST_net_17539), .b(FE_OFN1253_n_4143), .c(g62604_sb), .o(n_6344) );
na02f02 TIMEBOOST_cell_39617 ( .a(TIMEBOOST_net_11420), .b(g62782_sb), .o(n_5427) );
na02s01 TIMEBOOST_cell_70130 ( .a(TIMEBOOST_net_12808), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q), .o(TIMEBOOST_net_22273) );
in01f02 g57556_u0 ( .a(FE_OFN1416_n_8567), .o(g57556_sb) );
na03f02 TIMEBOOST_cell_1124 ( .a(n_4005), .b(g62833_sb), .c(g62833_db), .o(n_5308) );
in01f02 g57557_u0 ( .a(FE_OFN1377_n_8567), .o(g57557_sb) );
na03f02 TIMEBOOST_cell_66977 ( .a(FE_OFN1593_n_13741), .b(n_13901), .c(TIMEBOOST_net_13695), .o(n_16169) );
na02s02 TIMEBOOST_cell_47815 ( .a(g58270_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q), .o(TIMEBOOST_net_14125) );
na02m01 TIMEBOOST_cell_44542 ( .a(TIMEBOOST_net_13165), .b(g62865_sb), .o(n_5235) );
in01f02 g57558_u0 ( .a(FE_OFN2182_n_8567), .o(g57558_sb) );
na02s01 TIMEBOOST_cell_47630 ( .a(TIMEBOOST_net_14032), .b(TIMEBOOST_net_9651), .o(TIMEBOOST_net_12835) );
na03m04 TIMEBOOST_cell_72747 ( .a(n_4447), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q), .c(TIMEBOOST_net_9763), .o(TIMEBOOST_net_17505) );
na04f01 TIMEBOOST_cell_72417 ( .a(FE_OFN276_n_9941), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q), .c(g57797_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_), .o(TIMEBOOST_net_21316) );
in01f02 g57559_u0 ( .a(FE_OFN2175_n_8567), .o(g57559_sb) );
no03f02 TIMEBOOST_cell_72662 ( .a(FE_RN_741_0), .b(FE_RN_740_0), .c(n_14532), .o(n_14622) );
na02s01 TIMEBOOST_cell_68082 ( .a(parchk_pci_ad_reg_in_1216), .b(FE_OFN988_n_574), .o(TIMEBOOST_net_21249) );
na02f01 g64324_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(FE_OFN1034_n_4732), .o(g64324_db) );
in01f02 g57560_u0 ( .a(FE_OFN1391_n_8567), .o(g57560_sb) );
na03f02 TIMEBOOST_cell_25023 ( .a(n_10986), .b(FE_RN_32_0), .c(n_12588), .o(n_12850) );
na04f04 TIMEBOOST_cell_24563 ( .a(n_9205), .b(g57555_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q), .d(FE_OFN1402_n_8567), .o(n_10806) );
in01f02 g57561_u0 ( .a(FE_OFN1428_n_8567), .o(g57561_sb) );
na02f02 TIMEBOOST_cell_47591 ( .a(n_1998), .b(n_2390), .o(TIMEBOOST_net_14013) );
in01f02 g57562_u0 ( .a(FE_OFN2180_n_8567), .o(g57562_sb) );
na02m01 TIMEBOOST_cell_47925 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q), .o(TIMEBOOST_net_14180) );
na03f02 TIMEBOOST_cell_66545 ( .a(g53905_sb), .b(FE_OFN1332_n_13547), .c(TIMEBOOST_net_16794), .o(n_13536) );
na02s02 TIMEBOOST_cell_68421 ( .a(TIMEBOOST_net_21418), .b(FE_OFN952_n_2055), .o(TIMEBOOST_net_20823) );
in01f02 g57563_u0 ( .a(FE_OFN2188_n_8567), .o(g57563_sb) );
na02m02 TIMEBOOST_cell_48467 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q), .o(TIMEBOOST_net_14451) );
na04s03 TIMEBOOST_cell_73079 ( .a(g61887_sb), .b(TIMEBOOST_net_10779), .c(g65824_sb), .d(g61887_db), .o(n_8056) );
in01f02 g57564_u0 ( .a(FE_OFN1370_n_8567), .o(g57564_sb) );
na03f02 TIMEBOOST_cell_1123 ( .a(n_3969), .b(g62803_sb), .c(g62803_db), .o(n_5376) );
na02m04 TIMEBOOST_cell_39795 ( .a(g58331_db), .b(TIMEBOOST_net_11509), .o(n_9214) );
na02f02 TIMEBOOST_cell_44544 ( .a(TIMEBOOST_net_13166), .b(g63555_sb), .o(n_4922) );
in01f02 g57565_u0 ( .a(FE_OFN1345_n_8567), .o(g57565_sb) );
na03f02 TIMEBOOST_cell_47380 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_13688), .c(FE_OFN1581_n_12306), .o(n_12516) );
in01f02 g57566_u0 ( .a(FE_OFN2177_n_8567), .o(g57566_sb) );
na03f02 TIMEBOOST_cell_73567 ( .a(TIMEBOOST_net_17501), .b(FE_OFN1230_n_6391), .c(g62679_sb), .o(n_6181) );
na02m10 TIMEBOOST_cell_51643 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q), .o(TIMEBOOST_net_16039) );
in01f02 g57567_u0 ( .a(FE_OFN1384_n_8567), .o(g57567_sb) );
na03f02 TIMEBOOST_cell_25011 ( .a(FE_RN_230_0), .b(n_10885), .c(n_12565), .o(n_12827) );
in01f01 g57568_u0 ( .a(FE_OFN1394_n_8567), .o(g57568_sb) );
na03m04 TIMEBOOST_cell_68404 ( .a(g64216_sb), .b(pci_target_unit_fifos_pciw_addr_data_in_151), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q), .o(TIMEBOOST_net_21410) );
in01f02 g57569_u0 ( .a(FE_OFN1408_n_8567), .o(g57569_sb) );
na03m02 TIMEBOOST_cell_72949 ( .a(TIMEBOOST_net_17244), .b(g65727_sb), .c(FE_OFN699_n_7845), .o(TIMEBOOST_net_16953) );
na02s01 TIMEBOOST_cell_47951 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q), .b(pci_target_unit_fifos_pcir_data_in_174), .o(TIMEBOOST_net_14193) );
na02f02 TIMEBOOST_cell_44546 ( .a(TIMEBOOST_net_13167), .b(g63059_sb), .o(n_5132) );
in01f02 g57570_u0 ( .a(FE_OFN1387_n_8567), .o(g57570_sb) );
na02s01 TIMEBOOST_cell_49427 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q), .o(TIMEBOOST_net_14931) );
na02s02 TIMEBOOST_cell_47909 ( .a(TIMEBOOST_net_13873), .b(g65770_sb), .o(TIMEBOOST_net_14172) );
na03f02 TIMEBOOST_cell_73366 ( .a(TIMEBOOST_net_16714), .b(FE_OFN1299_n_5763), .c(g62059_sb), .o(n_7751) );
in01f02 g57571_u0 ( .a(FE_OFN1349_n_8567), .o(g57571_sb) );
na04f04 TIMEBOOST_cell_35194 ( .a(n_9334), .b(n_16986), .c(n_9335), .d(n_16987), .o(n_12166) );
in01f02 g57572_u0 ( .a(FE_OFN1391_n_8567), .o(g57572_sb) );
na02s01 TIMEBOOST_cell_44138 ( .a(TIMEBOOST_net_12963), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_11189) );
in01f02 g57573_u0 ( .a(FE_OFN2180_n_8567), .o(g57573_sb) );
na02f02 TIMEBOOST_cell_70838 ( .a(TIMEBOOST_net_16719), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_22627) );
na03f02 TIMEBOOST_cell_72823 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q), .b(g65338_sb), .c(TIMEBOOST_net_22254), .o(TIMEBOOST_net_17437) );
in01f02 g57574_u0 ( .a(FE_OFN1412_n_8567), .o(g57574_sb) );
na02s01 TIMEBOOST_cell_47623 ( .a(TIMEBOOST_net_6773), .b(g54205_sb), .o(TIMEBOOST_net_14029) );
na02s01 TIMEBOOST_cell_47769 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_14102) );
na02f01 TIMEBOOST_cell_69636 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q), .o(TIMEBOOST_net_22026) );
in01f02 g57575_u0 ( .a(FE_OFN1389_n_8567), .o(g57575_sb) );
na02m02 TIMEBOOST_cell_71899 ( .a(TIMEBOOST_net_23157), .b(g64833_sb), .o(TIMEBOOST_net_17388) );
in01f02 g57576_u0 ( .a(FE_OFN1387_n_8567), .o(g57576_sb) );
na02m02 TIMEBOOST_cell_53829 ( .a(TIMEBOOST_net_7630), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q), .o(TIMEBOOST_net_17132) );
na02m02 TIMEBOOST_cell_69954 ( .a(pci_target_unit_pcit_if_strd_addr_in_709), .b(g52638_sb), .o(TIMEBOOST_net_22185) );
in01f02 g57577_u0 ( .a(FE_OFN1387_n_8567), .o(g57577_sb) );
na02m01 TIMEBOOST_cell_52387 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q), .b(FE_OFN1076_n_4740), .o(TIMEBOOST_net_16411) );
na03m02 TIMEBOOST_cell_65438 ( .a(TIMEBOOST_net_10568), .b(g64777_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q), .o(TIMEBOOST_net_20957) );
in01f02 g57578_u0 ( .a(FE_OFN1382_n_8567), .o(g57578_sb) );
na04f04 TIMEBOOST_cell_67810 ( .a(FE_RN_622_0), .b(n_3404), .c(n_290), .d(FE_RN_623_0), .o(FE_RN_626_0) );
na03f02 TIMEBOOST_cell_73367 ( .a(TIMEBOOST_net_15225), .b(FE_OFN1300_n_5763), .c(g62064_sb), .o(n_7745) );
in01f02 g57579_u0 ( .a(FE_OFN1387_n_8567), .o(g57579_sb) );
na02m02 TIMEBOOST_cell_31743 ( .a(n_982), .b(TIMEBOOST_net_681), .o(TIMEBOOST_net_9976) );
na02f02 TIMEBOOST_cell_39473 ( .a(TIMEBOOST_net_11348), .b(g62850_sb), .o(n_5269) );
na02m01 TIMEBOOST_cell_69752 ( .a(pci_target_unit_del_sync_bc_in_203), .b(g65940_sb), .o(TIMEBOOST_net_22084) );
in01f02 g57580_u0 ( .a(FE_OFN1389_n_8567), .o(g57580_sb) );
na03f02 TIMEBOOST_cell_66914 ( .a(FE_OFN1735_n_16317), .b(TIMEBOOST_net_16490), .c(FE_OFN1741_n_11019), .o(n_12683) );
na02m02 TIMEBOOST_cell_38190 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q), .b(g65276_sb), .o(TIMEBOOST_net_10707) );
in01f02 g57581_u0 ( .a(FE_OFN2177_n_8567), .o(g57581_sb) );
na02m01 TIMEBOOST_cell_48055 ( .a(FE_OFN631_n_4454), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q), .o(TIMEBOOST_net_14245) );
na03f02 TIMEBOOST_cell_73289 ( .a(TIMEBOOST_net_16412), .b(FE_OFN1189_n_5742), .c(n_5732), .o(n_7721) );
na02f02 TIMEBOOST_cell_70263 ( .a(TIMEBOOST_net_22339), .b(g61842_sb), .o(n_6967) );
in01f02 g57582_u0 ( .a(FE_OFN2179_n_8567), .o(g57582_sb) );
na04m02 TIMEBOOST_cell_67297 ( .a(TIMEBOOST_net_20818), .b(g65097_sb), .c(n_4444), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_20597) );
na03f02 TIMEBOOST_cell_73603 ( .a(TIMEBOOST_net_17550), .b(FE_OFN2064_n_6391), .c(g62534_sb), .o(n_6504) );
na02f01 TIMEBOOST_cell_54440 ( .a(TIMEBOOST_net_17437), .b(FE_OFN1242_n_4092), .o(TIMEBOOST_net_15485) );
in01f02 g57583_u0 ( .a(FE_OFN1412_n_8567), .o(g57583_sb) );
na02s02 TIMEBOOST_cell_44454 ( .a(TIMEBOOST_net_13121), .b(TIMEBOOST_net_11217), .o(TIMEBOOST_net_9352) );
na03m02 TIMEBOOST_cell_69136 ( .a(g65429_sb), .b(n_4447), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q), .o(TIMEBOOST_net_21776) );
na02s01 TIMEBOOST_cell_63134 ( .a(FE_OFN533_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q), .o(TIMEBOOST_net_20514) );
in01f02 g57584_u0 ( .a(FE_OFN1396_n_8567), .o(g57584_sb) );
na02s01 TIMEBOOST_cell_47778 ( .a(TIMEBOOST_net_14106), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_399), .o(n_13179) );
na02f01 g64314_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(FE_OFN1034_n_4732), .o(g64314_db) );
no03f04 TIMEBOOST_cell_47135 ( .a(TIMEBOOST_net_13381), .b(n_4703), .c(FE_RN_285_0), .o(n_7094) );
in01f02 g57586_u0 ( .a(FE_OFN2170_n_8567), .o(g57586_sb) );
na04f04 TIMEBOOST_cell_24845 ( .a(wbs_dat_o_29_), .b(g52524_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_128), .d(FE_OFN2242_g52675_p), .o(n_13696) );
na02s02 TIMEBOOST_cell_39191 ( .a(TIMEBOOST_net_11207), .b(g57952_sb), .o(n_9837) );
in01f02 g57587_u0 ( .a(FE_OFN1391_n_8567), .o(g57587_sb) );
na03f02 TIMEBOOST_cell_67871 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q), .b(g64352_sb), .c(g64352_db), .o(TIMEBOOST_net_12961) );
na04f02 TIMEBOOST_cell_73216 ( .a(FE_OFN2022_n_4778), .b(TIMEBOOST_net_16650), .c(TIMEBOOST_net_633), .d(g63608_sb), .o(n_7159) );
in01f02 g57588_u0 ( .a(FE_OFN2184_n_8567), .o(g57588_sb) );
na02s01 TIMEBOOST_cell_39193 ( .a(TIMEBOOST_net_11208), .b(g57961_db), .o(n_9843) );
na03f02 TIMEBOOST_cell_71162 ( .a(TIMEBOOST_net_13387), .b(wishbone_slave_unit_del_sync_addr_out_reg_7__Q), .c(n_13221), .o(TIMEBOOST_net_22789) );
in01f02 g57589_u0 ( .a(FE_OFN1409_n_8567), .o(g57589_sb) );
na03f02 TIMEBOOST_cell_73710 ( .a(n_12010), .b(TIMEBOOST_net_13565), .c(FE_OFN1747_n_12004), .o(n_12727) );
na02s01 TIMEBOOST_cell_39195 ( .a(TIMEBOOST_net_11209), .b(g57948_db), .o(n_9861) );
in01f02 g57590_u0 ( .a(FE_OFN1374_n_8567), .o(g57590_sb) );
na02s01 TIMEBOOST_cell_52912 ( .a(TIMEBOOST_net_16673), .b(TIMEBOOST_net_10554), .o(TIMEBOOST_net_9414) );
na02s02 TIMEBOOST_cell_39197 ( .a(TIMEBOOST_net_11210), .b(g57956_db), .o(n_9850) );
na03m10 TIMEBOOST_cell_72730 ( .a(g64345_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q), .c(TIMEBOOST_net_21998), .o(TIMEBOOST_net_20926) );
in01f02 g57591_u0 ( .a(FE_OFN2170_n_8567), .o(g57591_sb) );
na02f02 TIMEBOOST_cell_71159 ( .a(TIMEBOOST_net_22787), .b(g54198_sb), .o(n_13420) );
na02s01 TIMEBOOST_cell_39189 ( .a(TIMEBOOST_net_11206), .b(g57979_db), .o(n_9820) );
in01f02 g57592_u0 ( .a(FE_OFN1412_n_8567), .o(g57592_sb) );
in01f02 g57593_u0 ( .a(FE_OFN1399_n_8567), .o(g57593_sb) );
na02f02 TIMEBOOST_cell_49306 ( .a(TIMEBOOST_net_14870), .b(g61747_sb), .o(n_8323) );
na02s02 TIMEBOOST_cell_68348 ( .a(TIMEBOOST_net_13909), .b(g65713_sb), .o(TIMEBOOST_net_21382) );
in01f02 g57594_u0 ( .a(FE_OFN1427_n_8567), .o(g57594_sb) );
na03f02 TIMEBOOST_cell_66809 ( .a(TIMEBOOST_net_16848), .b(FE_OFN1344_n_8567), .c(g57331_sb), .o(n_11419) );
in01f02 g57595_u0 ( .a(FE_OFN1425_n_8567), .o(g57595_sb) );
na02s01 TIMEBOOST_cell_49407 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_14921) );
na02s01 TIMEBOOST_cell_43163 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q), .o(TIMEBOOST_net_12476) );
in01f02 g57596_u0 ( .a(FE_OFN1402_n_8567), .o(g57596_sb) );
na03f02 TIMEBOOST_cell_34805 ( .a(TIMEBOOST_net_9554), .b(FE_OFN1381_n_8567), .c(g57411_sb), .o(n_10365) );
na03s02 TIMEBOOST_cell_72731 ( .a(TIMEBOOST_net_13883), .b(g65705_sb), .c(g65705_db), .o(n_1948) );
na03m06 TIMEBOOST_cell_72468 ( .a(TIMEBOOST_net_20181), .b(FE_OFN904_n_4736), .c(g64123_sb), .o(n_4038) );
in01f02 g57597_u0 ( .a(FE_OFN1416_n_8567), .o(g57597_sb) );
na02s01 TIMEBOOST_cell_71152 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q), .b(FE_OFN241_n_9830), .o(TIMEBOOST_net_22784) );
na02s01 TIMEBOOST_cell_47526 ( .a(TIMEBOOST_net_13980), .b(pci_target_unit_del_sync_comp_rty_exp_reg), .o(TIMEBOOST_net_10130) );
in01f02 g57598_u0 ( .a(FE_OFN1377_n_8567), .o(g57598_sb) );
na02f02 TIMEBOOST_cell_49182 ( .a(TIMEBOOST_net_14808), .b(g61886_sb), .o(n_8059) );
na02f01 TIMEBOOST_cell_27111 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q), .b(FE_OFN1128_g64577_p), .o(TIMEBOOST_net_7660) );
na02f02 g57641_u0 ( .a(n_8842), .b(FE_OFN276_n_9941), .o(n_9160) );
in01f04 g57644_u0 ( .a(n_8800), .o(n_8801) );
no02s01 g57646_u0 ( .a(n_3330), .b(FE_OFN778_n_4152), .o(n_4153) );
na02f02 g57648_u0 ( .a(n_8794), .b(pci_target_unit_fifos_pcir_flush_in), .o(n_8871) );
no02f02 g57649_u0 ( .a(n_3329), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8662) );
na02f04 g57654_u0 ( .a(n_16535), .b(n_8866), .o(n_16888) );
in01f08 g57667_u0 ( .a(n_8932), .o(n_10588) );
na02f06 g57668_u0 ( .a(n_16535), .b(n_16105), .o(n_8932) );
in01f08 g57671_u0 ( .a(n_15589), .o(n_10680) );
in01f06 g57676_u0 ( .a(n_16572), .o(n_9991) );
in01f08 g57698_u0 ( .a(n_8864), .o(n_10566) );
na02f06 g57699_u0 ( .a(n_8863), .b(n_8866), .o(n_8864) );
in01f06 g57700_u0 ( .a(n_8928), .o(n_9320) );
na02f06 g57710_u0 ( .a(n_16535), .b(n_16579), .o(n_8928) );
in01f06 g57725_u0 ( .a(n_8861), .o(n_9975) );
na02f06 g57726_u0 ( .a(n_16566), .b(n_8866), .o(n_8861) );
in01f10 g57734_u0 ( .a(FE_OCPN1905_n_8927), .o(n_11728) );
in01f04 g57735_u0 ( .a(FE_OCPN1905_n_8927), .o(n_10185) );
in01f03 g57736_u0 ( .a(FE_OCPN1905_n_8927), .o(n_10141) );
in01f04 g57737_u0 ( .a(FE_OCPN1905_n_8927), .o(n_10232) );
in01f01 g57738_u0 ( .a(n_8927), .o(n_10195) );
na02f03 g57739_u0 ( .a(n_8860), .b(n_16535), .o(n_8927) );
in01f08 g57747_u0 ( .a(n_9155), .o(n_10143) );
na02f08 g57751_u0 ( .a(n_8863), .b(n_15453), .o(n_9155) );
in01f08 g57755_u0 ( .a(n_8859), .o(n_10853) );
na02f06 g57756_u0 ( .a(n_8863), .b(n_8860), .o(n_8859) );
in01f02 g57759_u0 ( .a(n_15560), .o(n_10693) );
in01f04 g57770_u0 ( .a(n_8857), .o(n_10892) );
na02f06 g57771_u0 ( .a(n_8867), .b(n_8860), .o(n_8857) );
na02m10 TIMEBOOST_cell_52645 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_16540) );
na02f02 TIMEBOOST_cell_71049 ( .a(TIMEBOOST_net_22732), .b(g62387_sb), .o(n_6826) );
in01f20 g57780_u0 ( .a(pci_target_unit_fifos_pcir_flush_in), .o(g57780_sb) );
na02s01 TIMEBOOST_cell_44045 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q), .o(TIMEBOOST_net_12917) );
na02m01 TIMEBOOST_cell_69150 ( .a(n_4470), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q), .o(TIMEBOOST_net_21783) );
na03f02 TIMEBOOST_cell_73290 ( .a(TIMEBOOST_net_12981), .b(g63091_sb), .c(g63091_db), .o(n_5071) );
na04f04 TIMEBOOST_cell_24620 ( .a(n_9804), .b(g57119_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q), .d(FE_OFN2191_n_8567), .o(n_11626) );
na03m02 TIMEBOOST_cell_72575 ( .a(TIMEBOOST_net_21412), .b(FE_OFN664_n_4495), .c(TIMEBOOST_net_21536), .o(TIMEBOOST_net_20965) );
na04f02 TIMEBOOST_cell_67961 ( .a(n_4026), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q), .c(FE_OFN1134_g64577_p), .d(g62728_sb), .o(n_5523) );
na03f02 TIMEBOOST_cell_34909 ( .a(TIMEBOOST_net_9451), .b(FE_OFN1420_n_8567), .c(g57308_sb), .o(n_11442) );
na03m02 TIMEBOOST_cell_69124 ( .a(FE_OFN1640_n_4671), .b(g65369_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q), .o(TIMEBOOST_net_21770) );
na03m02 TIMEBOOST_cell_65889 ( .a(n_4737), .b(g62783_sb), .c(g62783_db), .o(n_7132) );
na02s01 TIMEBOOST_cell_28245 ( .a(FE_OFN243_n_9116), .b(g58033_sb), .o(TIMEBOOST_net_8227) );
na02s01 TIMEBOOST_cell_30969 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_18__Q), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_9589) );
na02m02 TIMEBOOST_cell_68423 ( .a(TIMEBOOST_net_21419), .b(TIMEBOOST_net_16165), .o(TIMEBOOST_net_17487) );
no02f06 TIMEBOOST_cell_4067 ( .a(TIMEBOOST_net_593), .b(FE_RN_838_0), .o(n_16511) );
no02f01 TIMEBOOST_cell_4068 ( .a(n_15645), .b(n_7114), .o(TIMEBOOST_net_594) );
na02m04 TIMEBOOST_cell_68634 ( .a(g65060_sb), .b(n_83), .o(TIMEBOOST_net_21525) );
na04f04 TIMEBOOST_cell_33807 ( .a(n_2201), .b(g61721_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q), .d(FE_OFN717_n_8176), .o(n_8382) );
na03f02 TIMEBOOST_cell_35049 ( .a(TIMEBOOST_net_9599), .b(FE_OFN1436_n_9372), .c(g58479_sb), .o(n_9358) );
na02m01 g57787_u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .b(g56933_sb), .o(g57787_da) );
na02f02 TIMEBOOST_cell_40361 ( .a(TIMEBOOST_net_11792), .b(n_4154), .o(n_13556) );
na02m01 g57788_u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .b(g56933_sb), .o(g57788_da) );
na02s01 TIMEBOOST_cell_68147 ( .a(TIMEBOOST_net_21281), .b(TIMEBOOST_net_6808), .o(TIMEBOOST_net_17194) );
na04m02 TIMEBOOST_cell_67301 ( .a(n_4476), .b(g64789_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q), .d(FE_OFN666_n_4495), .o(n_4477) );
na02s02 TIMEBOOST_cell_49087 ( .a(g58263_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q), .o(TIMEBOOST_net_14761) );
na02f02 TIMEBOOST_cell_47871 ( .a(g65851_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q), .o(TIMEBOOST_net_14153) );
na02m10 TIMEBOOST_cell_52865 ( .a(wbs_dat_i_5_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q), .o(TIMEBOOST_net_16650) );
in01f01 g57790_u0 ( .a(parchk_pci_cbe_en_in), .o(g57790_sb) );
na03f02 TIMEBOOST_cell_66549 ( .a(TIMEBOOST_net_21040), .b(FE_OFN1330_n_13547), .c(g53899_sb), .o(n_13546) );
na03f02 TIMEBOOST_cell_73537 ( .a(TIMEBOOST_net_17494), .b(FE_OFN1231_n_6391), .c(g62662_sb), .o(n_6216) );
na04f06 TIMEBOOST_cell_73179 ( .a(TIMEBOOST_net_20391), .b(FE_OFN1150_n_13249), .c(n_2114), .d(g54133_sb), .o(n_13672) );
na02s01 TIMEBOOST_cell_49408 ( .a(TIMEBOOST_net_14921), .b(FE_OFN563_n_9895), .o(TIMEBOOST_net_12969) );
na02m01 TIMEBOOST_cell_3982 ( .a(n_3395), .b(n_188), .o(TIMEBOOST_net_551) );
in01f08 g57792_u0 ( .a(n_9173), .o(n_9152) );
in01f10 g57794_u0 ( .a(n_8747), .o(g57794_sb) );
na02s01 TIMEBOOST_cell_48099 ( .a(pci_target_unit_pcit_if_strd_addr_in), .b(n_2671), .o(TIMEBOOST_net_14267) );
na02f20 g57794_u2 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q), .b(n_8747), .o(g57794_db) );
in01f04 g57795_u0 ( .a(FE_OFN276_n_9941), .o(g57795_sb) );
na03m02 TIMEBOOST_cell_69804 ( .a(n_4476), .b(g65392_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q), .o(TIMEBOOST_net_22110) );
na02m02 TIMEBOOST_cell_3983 ( .a(TIMEBOOST_net_551), .b(FE_OFN2121_n_2687), .o(TIMEBOOST_net_287) );
na03f02 TIMEBOOST_cell_73604 ( .a(TIMEBOOST_net_17486), .b(n_6645), .c(g63029_sb), .o(n_5860) );
na02f02 TIMEBOOST_cell_4051 ( .a(TIMEBOOST_net_585), .b(n_16452), .o(TIMEBOOST_net_403) );
no02s01 TIMEBOOST_cell_45297 ( .a(FE_RN_243_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236), .o(TIMEBOOST_net_13543) );
in01f02 g57797_u0 ( .a(FE_OFN276_n_9941), .o(g57797_sb) );
na04f02 TIMEBOOST_cell_73217 ( .a(FE_OFN2022_n_4778), .b(TIMEBOOST_net_16656), .c(TIMEBOOST_net_630), .d(g63620_sb), .o(n_7139) );
na03f02 TIMEBOOST_cell_66551 ( .a(TIMEBOOST_net_17568), .b(FE_OFN1330_n_13547), .c(g53919_sb), .o(n_13627) );
na02s02 TIMEBOOST_cell_48326 ( .a(TIMEBOOST_net_14380), .b(TIMEBOOST_net_10774), .o(TIMEBOOST_net_9474) );
na02s01 TIMEBOOST_cell_3712 ( .a(g57798_da), .b(FE_OFN276_n_9941), .o(TIMEBOOST_net_416) );
in01s01 TIMEBOOST_cell_73943 ( .a(TIMEBOOST_net_23507), .o(TIMEBOOST_net_23508) );
na02m01 TIMEBOOST_cell_3986 ( .a(n_188), .b(n_1459), .o(TIMEBOOST_net_553) );
na03f02 TIMEBOOST_cell_34787 ( .a(TIMEBOOST_net_9539), .b(FE_OFN1420_n_8567), .c(g57102_sb), .o(n_11644) );
na02f04 TIMEBOOST_cell_71928 ( .a(g64343_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q), .o(TIMEBOOST_net_23172) );
na02m10 TIMEBOOST_cell_52971 ( .a(wishbone_slave_unit_pcim_sm_data_in_660), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q), .o(TIMEBOOST_net_16703) );
no02s02 TIMEBOOST_cell_3990 ( .a(n_1667), .b(n_1995), .o(TIMEBOOST_net_555) );
no02f02 TIMEBOOST_cell_3991 ( .a(TIMEBOOST_net_555), .b(FE_OFN1024_n_11877), .o(n_3453) );
na02s02 TIMEBOOST_cell_49409 ( .a(FE_OFN1654_n_9502), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q), .o(TIMEBOOST_net_14922) );
na02s01 TIMEBOOST_cell_49461 ( .a(FE_OFN262_n_9851), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q), .o(TIMEBOOST_net_14948) );
na03m04 TIMEBOOST_cell_72798 ( .a(n_4452), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q), .c(TIMEBOOST_net_9706), .o(TIMEBOOST_net_20603) );
na02s01 TIMEBOOST_cell_3994 ( .a(wbs_adr_i_1_), .b(g52466_sb), .o(TIMEBOOST_net_557) );
in01f02 g57803_u0 ( .a(n_16368), .o(n_8926) );
na02s02 TIMEBOOST_cell_39188 ( .a(g57979_sb), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11206) );
na02f02 g57850_u0 ( .a(n_8571), .b(n_3363), .o(n_8688) );
na02s01 TIMEBOOST_cell_3197 ( .a(TIMEBOOST_net_158), .b(n_15390), .o(n_8746) );
na03f02 TIMEBOOST_cell_71350 ( .a(TIMEBOOST_net_660), .b(TIMEBOOST_net_657), .c(g54200_da), .o(TIMEBOOST_net_22883) );
na02f08 g57856_u0 ( .a(n_15515), .b(n_15517), .o(g57856_p) );
in01f08 g57856_u1 ( .a(g57856_p), .o(n_8939) );
in01f06 g57857_u0 ( .a(n_8924), .o(n_16605) );
na02f08 g57858_u0 ( .a(n_8790), .b(n_8792), .o(n_8924) );
na02f08 g57863_u0 ( .a(n_16537), .b(n_16534), .o(g57863_p) );
in01f08 g57863_u1 ( .a(g57863_p), .o(n_8863) );
na02f08 g57864_u0 ( .a(n_8686), .b(n_16533), .o(g57864_p) );
in01f08 g57864_u1 ( .a(g57864_p), .o(n_8867) );
no02f08 g57865_u0 ( .a(n_8790), .b(n_15517), .o(n_9171) );
in01f04 g57867_u0 ( .a(n_15581), .o(n_10258) );
oa12f02 g57871_u0 ( .a(n_9143), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .c(n_9144), .o(n_9146) );
oa12f02 g57872_u0 ( .a(n_8575), .b(pci_target_unit_pci_target_sm_rd_request), .c(FE_OFN2093_n_2301), .o(n_8687) );
na02s02 TIMEBOOST_cell_47893 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q), .b(FE_OFN937_n_2292), .o(TIMEBOOST_net_14164) );
oa12f02 g57874_u0 ( .a(n_9143), .b(wishbone_slave_unit_fifos_inGreyCount_0_), .c(n_9144), .o(n_9145) );
in01f01 g57875_u0 ( .a(n_9144), .o(g57875_sb) );
na02f02 TIMEBOOST_cell_37112 ( .a(n_692), .b(g53892_sb), .o(TIMEBOOST_net_10168) );
no02f01 g57876_u0 ( .a(n_3024), .b(pci_target_unit_del_sync_comp_cycle_count_12_), .o(g57876_p) );
ao12f01 g57876_u1 ( .a(g57876_p), .b(pci_target_unit_del_sync_comp_cycle_count_12_), .c(n_3024), .o(n_3330) );
ao12f02 g57877_u0 ( .a(n_5754), .b(conf_wb_err_addr_in_971), .c(FE_OFN1145_n_15261), .o(n_7362) );
no02m02 g57878_u0 ( .a(n_3073), .b(n_206), .o(g57878_p) );
ao12m02 g57878_u1 ( .a(g57878_p), .b(n_206), .c(n_3073), .o(n_3329) );
ao12s01 g57879_u0 ( .a(n_8971), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q), .c(FE_OFN601_n_9687), .o(n_9928) );
ao12s01 g57880_u0 ( .a(n_8970), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q), .c(FE_OFN562_n_9895), .o(n_9926) );
ao12s01 g57881_u0 ( .a(n_8968), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q), .c(FE_OFN554_n_9864), .o(n_9924) );
ao12s01 g57882_u0 ( .a(n_8967), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q), .c(FE_OFN519_n_9697), .o(n_9922) );
ao12s01 g57883_u0 ( .a(n_8966), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q), .c(FE_OFN587_n_9692), .o(n_9920) );
ao12s01 g57884_u0 ( .a(n_8965), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q), .c(FE_OFN532_n_9823), .o(n_9918) );
ao12s01 g57885_u0 ( .a(n_8964), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q), .c(FE_OFN595_n_9694), .o(n_9916) );
ao12s01 g57886_u0 ( .a(n_8963), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q), .c(FE_OFN529_n_9899), .o(n_9914) );
ao12s01 g57887_u0 ( .a(n_8962), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q), .c(FE_OFN606_n_9904), .o(n_9912) );
ao12s01 g57888_u0 ( .a(n_8961), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q), .c(FE_OFN1803_n_9690), .o(n_9910) );
ao12s01 g57889_u0 ( .a(n_8960), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q), .c(FE_OFN577_n_9902), .o(n_9908) );
in01m02 g57890_u0 ( .a(FE_OFN576_n_9902), .o(g57890_sb) );
in01s01 TIMEBOOST_cell_63577 ( .a(TIMEBOOST_net_20757), .o(TIMEBOOST_net_20756) );
in01s01 g57891_u0 ( .a(FE_OFN562_n_9895), .o(g57891_sb) );
na02s01 g57891_u2 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q), .o(g57891_db) );
na02s02 TIMEBOOST_cell_63888 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q), .b(FE_OFN229_n_9120), .o(TIMEBOOST_net_20930) );
in01s01 g57892_u0 ( .a(FE_OFN564_n_9895), .o(g57892_sb) );
na02f02 TIMEBOOST_cell_40060 ( .a(wbm_adr_o_16_), .b(g60691_sb), .o(TIMEBOOST_net_11642) );
na02s01 g57892_u2 ( .a(FE_OFN564_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q), .o(g57892_db) );
in01m01 g57893_u0 ( .a(FE_OFN562_n_9895), .o(g57893_sb) );
na02s01 g57893_u2 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q), .o(g57893_db) );
na02f02 TIMEBOOST_cell_70525 ( .a(TIMEBOOST_net_22470), .b(g62826_sb), .o(n_5325) );
in01s01 g57894_u0 ( .a(FE_OFN554_n_9864), .o(g57894_sb) );
na03m02 TIMEBOOST_cell_68670 ( .a(n_3747), .b(g64843_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q), .o(TIMEBOOST_net_21543) );
na02s01 g57894_u2 ( .a(FE_OFN554_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q), .o(g57894_db) );
na02f04 TIMEBOOST_cell_27798 ( .a(TIMEBOOST_net_8003), .b(n_3403), .o(n_4807) );
in01s01 g57895_u0 ( .a(FE_OFN556_n_9864), .o(g57895_sb) );
na02f02 TIMEBOOST_cell_71973 ( .a(TIMEBOOST_net_23194), .b(TIMEBOOST_net_12603), .o(TIMEBOOST_net_17404) );
na02s01 g57895_u2 ( .a(FE_OFN556_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q), .o(g57895_db) );
in01s01 g57896_u0 ( .a(FE_OFN554_n_9864), .o(g57896_sb) );
na03f03 TIMEBOOST_cell_35013 ( .a(TIMEBOOST_net_7995), .b(n_7095), .c(n_7724), .o(n_8576) );
na03m04 TIMEBOOST_cell_73089 ( .a(g65389_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q), .c(TIMEBOOST_net_16329), .o(TIMEBOOST_net_17398) );
na02s03 TIMEBOOST_cell_53231 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_789), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q), .o(TIMEBOOST_net_16833) );
in01s01 g57897_u0 ( .a(FE_OFN532_n_9823), .o(g57897_sb) );
na02s01 g57897_u2 ( .a(FE_OFN532_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q), .o(g57897_db) );
na03f02 TIMEBOOST_cell_66690 ( .a(TIMEBOOST_net_17564), .b(FE_OFN1278_n_4097), .c(g62526_sb), .o(n_6523) );
in01s01 g57898_u0 ( .a(FE_OFN534_n_9823), .o(g57898_sb) );
na02s01 g57898_u2 ( .a(FE_OFN534_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q), .o(g57898_db) );
in01s01 g57899_u0 ( .a(FE_OFN532_n_9823), .o(g57899_sb) );
na02s02 g57899_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q), .b(FE_OFN532_n_9823), .o(g57899_db) );
na02f04 TIMEBOOST_cell_70383 ( .a(TIMEBOOST_net_22399), .b(n_2795), .o(n_8448) );
in01s01 g57900_u0 ( .a(FE_OFN529_n_9899), .o(g57900_sb) );
na03s02 TIMEBOOST_cell_65773 ( .a(TIMEBOOST_net_10838), .b(n_8272), .c(g61865_sb), .o(n_8107) );
na02f02 TIMEBOOST_cell_47872 ( .a(TIMEBOOST_net_14153), .b(g65851_db), .o(n_2184) );
na02s02 TIMEBOOST_cell_69304 ( .a(TIMEBOOST_net_17226), .b(FE_OFN956_n_1699), .o(TIMEBOOST_net_21860) );
in01s01 g57901_u0 ( .a(FE_OFN528_n_9899), .o(g57901_sb) );
na02m02 TIMEBOOST_cell_68671 ( .a(TIMEBOOST_net_21543), .b(g64843_db), .o(TIMEBOOST_net_17529) );
na02s01 g57901_u2 ( .a(FE_OFN528_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q), .o(g57901_db) );
na03f01 TIMEBOOST_cell_65128 ( .a(n_3777), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q), .c(FE_OFN660_n_4392), .o(TIMEBOOST_net_14418) );
in01s01 g57902_u0 ( .a(FE_OFN529_n_9899), .o(g57902_sb) );
na03f02 TIMEBOOST_cell_64586 ( .a(n_2212), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q), .c(FE_OFN720_n_8060), .o(TIMEBOOST_net_15047) );
na03f02 TIMEBOOST_cell_71690 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q), .c(n_13997), .o(TIMEBOOST_net_23053) );
in01s01 g57903_u0 ( .a(FE_OFN606_n_9904), .o(g57903_sb) );
na02f02 TIMEBOOST_cell_72257 ( .a(TIMEBOOST_net_23336), .b(g60656_sb), .o(n_5666) );
na02m04 TIMEBOOST_cell_71879 ( .a(TIMEBOOST_net_23147), .b(n_3741), .o(TIMEBOOST_net_16205) );
na03f10 TIMEBOOST_cell_72385 ( .a(n_2426), .b(n_2433), .c(n_2441), .o(n_2434) );
in01s01 g57904_u0 ( .a(FE_OFN606_n_9904), .o(g57904_sb) );
na02f02 TIMEBOOST_cell_51375 ( .a(FE_OFN1186_n_3476), .b(configuration_pci_err_cs_bit10), .o(TIMEBOOST_net_15905) );
na02s01 g57904_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q), .b(FE_OFN606_n_9904), .o(g57904_db) );
in01s01 g57905_u0 ( .a(FE_OFN606_n_9904), .o(g57905_sb) );
na02f02 TIMEBOOST_cell_70197 ( .a(TIMEBOOST_net_22306), .b(FE_OFN2126_n_16497), .o(n_13027) );
na02s02 TIMEBOOST_cell_70887 ( .a(TIMEBOOST_net_22651), .b(TIMEBOOST_net_12918), .o(TIMEBOOST_net_21004) );
in01s01 g57906_u0 ( .a(FE_OFN576_n_9902), .o(g57906_sb) );
in01s01 TIMEBOOST_cell_73931 ( .a(TIMEBOOST_net_23495), .o(TIMEBOOST_net_23496) );
na02s01 g57906_u2 ( .a(FE_OFN576_n_9902), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q), .o(g57906_db) );
in01s01 g57907_u0 ( .a(FE_OFN576_n_9902), .o(g57907_sb) );
na03f02 TIMEBOOST_cell_70046 ( .a(n_4523), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q), .c(FE_OFN706_n_8119), .o(TIMEBOOST_net_22231) );
na02s01 g57907_u2 ( .a(FE_OFN576_n_9902), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q), .o(g57907_db) );
in01s01 TIMEBOOST_cell_73961 ( .a(TIMEBOOST_net_23525), .o(TIMEBOOST_net_23526) );
in01f01 g57908_u0 ( .a(n_9144), .o(g57908_sb) );
na03s02 TIMEBOOST_cell_72714 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q), .b(g64328_sb), .c(g64328_db), .o(n_3848) );
na03m02 TIMEBOOST_cell_73121 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q), .b(g64347_sb), .c(TIMEBOOST_net_12933), .o(n_3830) );
in01s02 g57909_u0 ( .a(FE_OFN1795_n_9904), .o(g57909_sb) );
na02s01 g57909_u2 ( .a(FE_OFN1795_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q), .o(g57909_db) );
na02f02 TIMEBOOST_cell_70960 ( .a(TIMEBOOST_net_17390), .b(FE_OFN1264_n_4095), .o(TIMEBOOST_net_22688) );
in01m02 g57910_u0 ( .a(FE_OFN576_n_9902), .o(g57910_sb) );
na02f02 TIMEBOOST_cell_51912 ( .a(TIMEBOOST_net_16173), .b(g67040_sb), .o(n_2471) );
na02m01 TIMEBOOST_cell_62588 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q), .b(n_3792), .o(TIMEBOOST_net_20241) );
na03f02 TIMEBOOST_cell_65188 ( .a(TIMEBOOST_net_12615), .b(g64291_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q), .o(TIMEBOOST_net_15067) );
in01s01 g57911_u0 ( .a(FE_OFN527_n_9899), .o(g57911_sb) );
na03f02 TIMEBOOST_cell_35014 ( .a(TIMEBOOST_net_10015), .b(FE_OFN2180_n_8567), .c(g57567_sb), .o(n_11186) );
na02s01 g57911_u2 ( .a(FE_OFN527_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q), .o(g57911_db) );
na03f06 TIMEBOOST_cell_35015 ( .a(TIMEBOOST_net_9578), .b(FE_OFN2179_n_8567), .c(g57445_sb), .o(n_11287) );
in01s01 g57912_u0 ( .a(FE_OFN576_n_9902), .o(g57912_sb) );
na02s01 TIMEBOOST_cell_37780 ( .a(g57954_sb), .b(FE_OFN219_n_9853), .o(TIMEBOOST_net_10502) );
na02s01 g57912_u2 ( .a(FE_OFN576_n_9902), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q), .o(g57912_db) );
in01s01 g57913_u0 ( .a(FE_OFN1794_n_9904), .o(g57913_sb) );
na02s01 TIMEBOOST_cell_44455 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q), .o(TIMEBOOST_net_13122) );
na02m02 TIMEBOOST_cell_68867 ( .a(TIMEBOOST_net_21641), .b(g64980_db), .o(TIMEBOOST_net_17538) );
na02s01 TIMEBOOST_cell_38397 ( .a(TIMEBOOST_net_10810), .b(g58130_db), .o(n_9663) );
in01s01 g57914_u0 ( .a(FE_OFN562_n_9895), .o(g57914_sb) );
in01s01 TIMEBOOST_cell_63580 ( .a(TIMEBOOST_net_20759), .o(TIMEBOOST_net_20760) );
na02m01 TIMEBOOST_cell_68190 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q), .b(g65959_db), .o(TIMEBOOST_net_21303) );
in01s01 g57915_u0 ( .a(FE_OFN563_n_9895), .o(g57915_sb) );
na03f02 TIMEBOOST_cell_35016 ( .a(TIMEBOOST_net_9579), .b(FE_OFN2179_n_8567), .c(g57537_sb), .o(n_11205) );
na04m08 TIMEBOOST_cell_67173 ( .a(n_3755), .b(FE_OFN672_n_4505), .c(g64782_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q), .o(n_3768) );
na03f02 TIMEBOOST_cell_35017 ( .a(TIMEBOOST_net_9580), .b(FE_OFN1428_n_8567), .c(g57444_sb), .o(n_11289) );
in01m01 g57916_u0 ( .a(FE_OFN561_n_9895), .o(g57916_sb) );
na03m08 TIMEBOOST_cell_64755 ( .a(g65316_sb), .b(FE_OFN1642_n_4671), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q), .o(TIMEBOOST_net_16339) );
na02f02 TIMEBOOST_cell_50540 ( .a(TIMEBOOST_net_15487), .b(g62335_sb), .o(n_6929) );
in01s01 g57917_u0 ( .a(FE_OFN560_n_9895), .o(g57917_sb) );
na02f01 TIMEBOOST_cell_31104 ( .a(TIMEBOOST_net_9656), .b(n_1096), .o(TIMEBOOST_net_286) );
na03f02 TIMEBOOST_cell_66553 ( .a(FE_OFN1327_n_13547), .b(g53917_sb), .c(TIMEBOOST_net_16805), .o(n_13525) );
in01s01 g57918_u0 ( .a(FE_OFN562_n_9895), .o(g57918_sb) );
na02m02 TIMEBOOST_cell_69885 ( .a(TIMEBOOST_net_22150), .b(g64200_db), .o(n_3969) );
na03f02 TIMEBOOST_cell_66875 ( .a(FE_OFN1565_n_12502), .b(TIMEBOOST_net_15988), .c(n_12313), .o(n_12620) );
in01s01 g57919_u0 ( .a(FE_OFN564_n_9895), .o(g57919_sb) );
na02s01 TIMEBOOST_cell_42796 ( .a(TIMEBOOST_net_12292), .b(FE_OFN935_n_2292), .o(TIMEBOOST_net_10231) );
na02s01 g57919_u2 ( .a(FE_OFN564_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q), .o(g57919_db) );
na03m02 TIMEBOOST_cell_72600 ( .a(TIMEBOOST_net_23154), .b(FE_OFN615_n_4501), .c(TIMEBOOST_net_21705), .o(TIMEBOOST_net_17026) );
in01s01 g57920_u0 ( .a(FE_OFN564_n_9895), .o(g57920_sb) );
na02s01 g57920_u2 ( .a(FE_OFN564_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q), .o(g57920_db) );
in01s01 g57921_u0 ( .a(FE_OFN562_n_9895), .o(g57921_sb) );
na02s01 TIMEBOOST_cell_31130 ( .a(TIMEBOOST_net_9669), .b(g65760_db), .o(n_1603) );
in01s01 g57922_u0 ( .a(FE_OFN561_n_9895), .o(g57922_sb) );
na04s02 TIMEBOOST_cell_72900 ( .a(g61736_sb), .b(g61736_db), .c(g65753_db), .d(TIMEBOOST_net_10347), .o(n_8346) );
na02s01 g57922_u2 ( .a(FE_OFN561_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q), .o(g57922_db) );
na03m02 TIMEBOOST_cell_72748 ( .a(TIMEBOOST_net_14334), .b(g65740_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q), .o(TIMEBOOST_net_22034) );
in01s02 g57923_u0 ( .a(FE_OFN563_n_9895), .o(g57923_sb) );
na02s01 g57923_u2 ( .a(FE_OFN563_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q), .o(g57923_db) );
na03f02 TIMEBOOST_cell_73793 ( .a(TIMEBOOST_net_16529), .b(FE_OFN1599_n_13995), .c(FE_OFN1606_n_13997), .o(g53159_p) );
in01s01 g57924_u0 ( .a(FE_OFN562_n_9895), .o(g57924_sb) );
na02f02 TIMEBOOST_cell_28291 ( .a(n_2675), .b(n_1251), .o(TIMEBOOST_net_8250) );
na02s01 g57924_u2 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q), .o(g57924_db) );
na02f04 TIMEBOOST_cell_28292 ( .a(TIMEBOOST_net_8250), .b(TIMEBOOST_net_193), .o(n_15292) );
in01m01 g57925_u0 ( .a(FE_OFN562_n_9895), .o(g57925_sb) );
na03f02 TIMEBOOST_cell_66047 ( .a(TIMEBOOST_net_16674), .b(n_7618), .c(g59809_sb), .o(n_7614) );
na02s01 TIMEBOOST_cell_53954 ( .a(TIMEBOOST_net_17194), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_390), .o(TIMEBOOST_net_9190) );
in01s01 g57926_u0 ( .a(FE_OFN563_n_9895), .o(g57926_sb) );
na03f02 TIMEBOOST_cell_66594 ( .a(TIMEBOOST_net_16781), .b(FE_OFN1317_n_6624), .c(g62519_sb), .o(n_6538) );
na02s01 g57926_u2 ( .a(FE_OFN563_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q), .o(g57926_db) );
na03f02 TIMEBOOST_cell_66555 ( .a(TIMEBOOST_net_21042), .b(FE_OFN1330_n_13547), .c(g53898_sb), .o(n_13550) );
in01m02 g57927_u0 ( .a(FE_OFN562_n_9895), .o(g57927_sb) );
na02m01 TIMEBOOST_cell_48074 ( .a(TIMEBOOST_net_14254), .b(FE_OFN927_n_4730), .o(TIMEBOOST_net_12634) );
na02m02 g57927_u2 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q), .o(g57927_db) );
na02f02 TIMEBOOST_cell_70243 ( .a(TIMEBOOST_net_22329), .b(g63165_sb), .o(n_4957) );
in01s01 g57928_u0 ( .a(FE_OFN563_n_9895), .o(g57928_sb) );
na04f04 TIMEBOOST_cell_67696 ( .a(TIMEBOOST_net_16856), .b(FE_OFN2200_n_10256), .c(g52612_sb), .d(TIMEBOOST_net_706), .o(n_11859) );
in01s01 g57929_u0 ( .a(FE_OFN561_n_9895), .o(g57929_sb) );
na04m02 TIMEBOOST_cell_67898 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(FE_OFN1041_n_2037), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q), .d(g65840_sb), .o(n_2017) );
na02s01 g57929_u2 ( .a(FE_OFN561_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q), .o(g57929_db) );
na02s01 TIMEBOOST_cell_25307 ( .a(pci_ad_i_7_), .b(parchk_pci_ad_reg_in_1211), .o(TIMEBOOST_net_6758) );
in01s01 g57930_u0 ( .a(FE_OFN561_n_9895), .o(g57930_sb) );
na03s02 TIMEBOOST_cell_67830 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q), .b(FE_OFN539_n_9690), .c(g58230_sb), .o(TIMEBOOST_net_14470) );
na02s01 g57930_u2 ( .a(FE_OFN561_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q), .o(g57930_db) );
na02s01 TIMEBOOST_cell_30985 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_11__Q), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_9597) );
in01s02 g57931_u0 ( .a(FE_OFN560_n_9895), .o(g57931_sb) );
na02f01 TIMEBOOST_cell_48076 ( .a(TIMEBOOST_net_14255), .b(FE_OFN929_n_4730), .o(TIMEBOOST_net_12615) );
na02s03 TIMEBOOST_cell_62980 ( .a(TIMEBOOST_net_13841), .b(configuration_wb_err_addr_540), .o(TIMEBOOST_net_20437) );
na02s01 TIMEBOOST_cell_30987 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_7__Q), .b(FE_OFN250_n_9789), .o(TIMEBOOST_net_9598) );
in01m02 g57932_u0 ( .a(FE_OFN561_n_9895), .o(g57932_sb) );
na02s02 TIMEBOOST_cell_37241 ( .a(TIMEBOOST_net_10232), .b(g65776_sb), .o(n_2191) );
na02f01 TIMEBOOST_cell_45058 ( .a(TIMEBOOST_net_13423), .b(g63191_sb), .o(n_4941) );
na03m04 TIMEBOOST_cell_69162 ( .a(FE_OFN927_n_4730), .b(pci_target_unit_fifos_pciw_cbe_in_153), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q), .o(TIMEBOOST_net_21789) );
in01s01 g57933_u0 ( .a(FE_OFN563_n_9895), .o(g57933_sb) );
na03f02 TIMEBOOST_cell_72516 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q), .b(g65934_sb), .c(g65934_db), .o(n_2170) );
na02f01 TIMEBOOST_cell_69718 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q), .b(FE_OFN1676_n_4655), .o(TIMEBOOST_net_22067) );
na03f02 TIMEBOOST_cell_66906 ( .a(FE_OFN1734_n_16317), .b(TIMEBOOST_net_16489), .c(FE_OFN1740_n_11019), .o(n_12500) );
in01s01 g57934_u0 ( .a(FE_OFN564_n_9895), .o(g57934_sb) );
na04f04 TIMEBOOST_cell_35196 ( .a(n_9956), .b(n_16838), .c(n_16839), .d(n_10533), .o(n_12129) );
na02s01 TIMEBOOST_cell_50729 ( .a(g58436_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q), .o(TIMEBOOST_net_15582) );
na02m01 TIMEBOOST_cell_53233 ( .a(n_13145), .b(pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77), .o(TIMEBOOST_net_16834) );
in01m01 g57935_u0 ( .a(FE_OFN563_n_9895), .o(g57935_sb) );
na02s01 TIMEBOOST_cell_42800 ( .a(TIMEBOOST_net_12294), .b(FE_OFN937_n_2292), .o(TIMEBOOST_net_10233) );
na02s01 g57935_u2 ( .a(FE_OFN563_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q), .o(g57935_db) );
na02m04 TIMEBOOST_cell_69066 ( .a(n_3785), .b(n_15), .o(TIMEBOOST_net_21741) );
in01m01 g57936_u0 ( .a(FE_OFN562_n_9895), .o(g57936_sb) );
na03f02 TIMEBOOST_cell_66578 ( .a(TIMEBOOST_net_17434), .b(FE_OFN1249_n_4093), .c(g62497_sb), .o(n_6589) );
na02s01 TIMEBOOST_cell_48849 ( .a(FE_OFN239_n_9832), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q), .o(TIMEBOOST_net_14642) );
in01s01 g57937_u0 ( .a(FE_OFN562_n_9895), .o(g57937_sb) );
na02m02 g52471_u1 ( .a(wbs_adr_i_25_), .b(g52459_sb), .o(g52471_da) );
na03f02 TIMEBOOST_cell_66557 ( .a(g53926_sb), .b(FE_OFN1327_n_13547), .c(TIMEBOOST_net_16808), .o(n_13519) );
na02s01 TIMEBOOST_cell_71132 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q), .b(FE_OFN554_n_9864), .o(TIMEBOOST_net_22774) );
in01s01 g57938_u0 ( .a(FE_OFN564_n_9895), .o(g57938_sb) );
na02m01 TIMEBOOST_cell_62452 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_146), .o(TIMEBOOST_net_20173) );
na02s01 g57938_u2 ( .a(FE_OFN564_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q), .o(g57938_db) );
in01s02 g57939_u0 ( .a(FE_OFN560_n_9895), .o(g57939_sb) );
na02m01 TIMEBOOST_cell_54069 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_125), .o(TIMEBOOST_net_17252) );
in01m02 g57940_u0 ( .a(FE_OFN562_n_9895), .o(g57940_sb) );
na02s01 g57940_u2 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q), .o(g57940_db) );
na02m04 TIMEBOOST_cell_69038 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q), .b(FE_OFN1640_n_4671), .o(TIMEBOOST_net_21727) );
in01s01 g57941_u0 ( .a(FE_OFN564_n_9895), .o(g57941_sb) );
na02s01 TIMEBOOST_cell_30989 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_31__Q), .b(FE_OFN241_n_9830), .o(TIMEBOOST_net_9599) );
na02s01 g57941_u2 ( .a(FE_OFN564_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q), .o(g57941_db) );
in01s02 g57942_u0 ( .a(FE_OFN559_n_9895), .o(g57942_sb) );
na03f02 TIMEBOOST_cell_73032 ( .a(TIMEBOOST_net_21740), .b(g64927_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q), .o(TIMEBOOST_net_17053) );
na02s02 TIMEBOOST_cell_53913 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q), .b(g58315_sb), .o(TIMEBOOST_net_17174) );
na03m02 TIMEBOOST_cell_72833 ( .a(g65307_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q), .c(TIMEBOOST_net_16251), .o(TIMEBOOST_net_13368) );
na02m01 TIMEBOOST_cell_63690 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q), .o(TIMEBOOST_net_20831) );
na02m02 TIMEBOOST_cell_68817 ( .a(TIMEBOOST_net_21616), .b(n_4476), .o(TIMEBOOST_net_16268) );
in01s01 g57944_u0 ( .a(FE_OFN564_n_9895), .o(g57944_sb) );
in01s01 TIMEBOOST_cell_73992 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .o(TIMEBOOST_net_23557) );
na02s01 g57944_u2 ( .a(FE_OFN564_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q), .o(g57944_db) );
na03f02 TIMEBOOST_cell_66728 ( .a(TIMEBOOST_net_16823), .b(FE_OFN1305_n_13124), .c(g54362_sb), .o(n_13080) );
in01m01 g57945_u0 ( .a(FE_OFN561_n_9895), .o(g57945_sb) );
na02s01 g57945_u2 ( .a(FE_OFN561_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q), .o(g57945_db) );
na03s02 TIMEBOOST_cell_48757 ( .a(TIMEBOOST_net_10300), .b(g65777_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q), .o(TIMEBOOST_net_14596) );
in01s01 g57946_u0 ( .a(FE_OFN554_n_9864), .o(g57946_sb) );
na03m02 TIMEBOOST_cell_65129 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q), .b(n_3770), .c(FE_OFN649_n_4497), .o(TIMEBOOST_net_10726) );
na03f02 TIMEBOOST_cell_66560 ( .a(g53918_sb), .b(FE_OFN1327_n_13547), .c(TIMEBOOST_net_16804), .o(n_13469) );
in01s01 g57947_u0 ( .a(FE_OFN555_n_9864), .o(g57947_sb) );
na04m08 TIMEBOOST_cell_67912 ( .a(FE_OFN1648_n_9428), .b(FE_OFN211_n_9858), .c(TIMEBOOST_net_12910), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q), .o(TIMEBOOST_net_16843) );
in01s01 g57948_u0 ( .a(FE_OFN553_n_9864), .o(g57948_sb) );
na03f04 TIMEBOOST_cell_73484 ( .a(wbm_adr_o_20_), .b(g61855_sb), .c(g52396_sb), .o(TIMEBOOST_net_23348) );
na02s01 g57948_u2 ( .a(FE_OFN553_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q), .o(g57948_db) );
na02s01 TIMEBOOST_cell_43647 ( .a(pci_target_unit_del_sync_addr_in_217), .b(parchk_pci_ad_reg_in_1218), .o(TIMEBOOST_net_12718) );
in01s01 g57949_u0 ( .a(FE_OFN551_n_9864), .o(g57949_sb) );
na03f02 TIMEBOOST_cell_73605 ( .a(TIMEBOOST_net_17566), .b(FE_OFN1259_n_4143), .c(g62342_sb), .o(n_6915) );
na03f02 TIMEBOOST_cell_66231 ( .a(TIMEBOOST_net_20955), .b(FE_OFN1264_n_4095), .c(g62698_sb), .o(n_6158) );
na02m02 TIMEBOOST_cell_69422 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q), .b(FE_OFN649_n_4497), .o(TIMEBOOST_net_21919) );
na02s01 g57950_u2 ( .a(FE_OFN555_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q), .o(g57950_db) );
na02f02 TIMEBOOST_cell_50308 ( .a(TIMEBOOST_net_15371), .b(g62672_sb), .o(n_6195) );
in01s01 g57951_u0 ( .a(FE_OFN556_n_9864), .o(g57951_sb) );
na04f08 TIMEBOOST_cell_73218 ( .a(TIMEBOOST_net_14987), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q), .c(FE_OFN1147_n_13249), .d(g54158_sb), .o(g53891_da) );
na02s01 g57951_u2 ( .a(FE_OFN556_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q), .o(g57951_db) );
in01s01 g57952_u0 ( .a(FE_OFN556_n_9864), .o(g57952_sb) );
na02s01 g57952_u2 ( .a(FE_OFN556_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q), .o(g57952_db) );
na03m06 TIMEBOOST_cell_67820 ( .a(n_3780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q), .c(FE_OFN652_n_4508), .o(TIMEBOOST_net_14413) );
in01s01 g57953_u0 ( .a(FE_OFN554_n_9864), .o(g57953_sb) );
na03f02 TIMEBOOST_cell_35019 ( .a(TIMEBOOST_net_9582), .b(FE_OFN1428_n_8567), .c(g57370_sb), .o(n_11380) );
na02s01 g57953_u2 ( .a(FE_OFN554_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q), .o(g57953_db) );
na03f02 TIMEBOOST_cell_35018 ( .a(TIMEBOOST_net_9581), .b(FE_OFN2179_n_8567), .c(g57210_sb), .o(n_11546) );
in01s01 g57954_u0 ( .a(FE_OFN553_n_9864), .o(g57954_sb) );
na02s01 g57954_u2 ( .a(FE_OFN553_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q), .o(g57954_db) );
na03f02 TIMEBOOST_cell_34738 ( .a(TIMEBOOST_net_9504), .b(FE_OFN1377_n_8567), .c(g57061_sb), .o(n_10506) );
na02m10 g57955_u2 ( .a(FE_OFN555_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q), .o(g57955_db) );
na03f02 TIMEBOOST_cell_34739 ( .a(TIMEBOOST_net_9505), .b(FE_OFN1413_n_8567), .c(g57231_sb), .o(n_10433) );
in01s02 g57956_u0 ( .a(FE_OFN554_n_9864), .o(g57956_sb) );
na03f02 TIMEBOOST_cell_34740 ( .a(TIMEBOOST_net_9506), .b(FE_OFN1397_n_8567), .c(g57212_sb), .o(n_10439) );
na02s02 g57956_u2 ( .a(FE_OFN554_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q), .o(g57956_db) );
na03f02 TIMEBOOST_cell_34741 ( .a(TIMEBOOST_net_9558), .b(FE_OFN1383_n_8567), .c(g57294_sb), .o(n_11458) );
in01s01 g57957_u0 ( .a(FE_OFN554_n_9864), .o(g57957_sb) );
na04s04 TIMEBOOST_cell_41376 ( .a(g58116_sb), .b(g58116_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q), .d(FE_OFN264_n_9849), .o(TIMEBOOST_net_9393) );
na02s02 g57957_u2 ( .a(FE_OFN554_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q), .o(g57957_db) );
na03f02 TIMEBOOST_cell_34831 ( .a(TIMEBOOST_net_9444), .b(FE_OFN1392_n_8567), .c(g57267_sb), .o(n_11485) );
in01s01 g57958_u0 ( .a(FE_OFN555_n_9864), .o(g57958_sb) );
na02f01 TIMEBOOST_cell_54214 ( .a(TIMEBOOST_net_17324), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_15144) );
na02s01 g57958_u2 ( .a(FE_OFN555_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q), .o(g57958_db) );
in01s02 g57959_u0 ( .a(FE_OFN554_n_9864), .o(g57959_sb) );
na02m01 TIMEBOOST_cell_49400 ( .a(TIMEBOOST_net_14917), .b(TIMEBOOST_net_566), .o(n_2588) );
na03f02 TIMEBOOST_cell_66727 ( .a(TIMEBOOST_net_16834), .b(FE_OFN1306_n_13124), .c(g54244_sb), .o(n_13146) );
na03f02 TIMEBOOST_cell_72871 ( .a(configuration_wb_err_addr_558), .b(n_15445), .c(n_2768), .o(TIMEBOOST_net_20658) );
na02s02 TIMEBOOST_cell_49088 ( .a(TIMEBOOST_net_14761), .b(TIMEBOOST_net_11001), .o(TIMEBOOST_net_9383) );
na02s01 g57960_u2 ( .a(FE_OFN555_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q), .o(g57960_db) );
in01s01 g57961_u0 ( .a(FE_OFN553_n_9864), .o(g57961_sb) );
na02m10 TIMEBOOST_cell_53567 ( .a(configuration_pci_err_cs_bit_464), .b(pci_target_unit_wishbone_master_bc_register_reg_1__Q), .o(TIMEBOOST_net_17001) );
na02s01 g57961_u2 ( .a(FE_OFN553_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q), .o(g57961_db) );
na03m02 TIMEBOOST_cell_65270 ( .a(g64243_sb), .b(FE_OFN1056_n_4727), .c(TIMEBOOST_net_16931), .o(n_3929) );
na02s02 TIMEBOOST_cell_43654 ( .a(TIMEBOOST_net_12721), .b(FE_OFN1801_n_9690), .o(TIMEBOOST_net_11001) );
na02s01 g57962_u2 ( .a(FE_OFN553_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q), .o(g57962_db) );
na02s10 TIMEBOOST_cell_62660 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q), .b(TIMEBOOST_net_13865), .o(TIMEBOOST_net_20277) );
na03f02 TIMEBOOST_cell_70694 ( .a(n_3947), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q), .c(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_22555) );
na04m06 TIMEBOOST_cell_72695 ( .a(FE_OFN682_n_4460), .b(g65080_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q), .d(n_4645), .o(n_4307) );
na03m04 TIMEBOOST_cell_72594 ( .a(TIMEBOOST_net_21435), .b(g64804_sb), .c(TIMEBOOST_net_21640), .o(TIMEBOOST_net_17485) );
in01f06 g57964_u0 ( .a(FE_OFN555_n_9864), .o(g57964_sb) );
na02f02 TIMEBOOST_cell_68999 ( .a(TIMEBOOST_net_21707), .b(TIMEBOOST_net_20293), .o(TIMEBOOST_net_17055) );
na02m02 TIMEBOOST_cell_53914 ( .a(TIMEBOOST_net_17174), .b(TIMEBOOST_net_11192), .o(TIMEBOOST_net_9406) );
na03f02 TIMEBOOST_cell_73538 ( .a(TIMEBOOST_net_17517), .b(FE_OFN1233_n_6391), .c(g62606_sb), .o(n_6340) );
in01s01 g57965_u0 ( .a(FE_OFN555_n_9864), .o(g57965_sb) );
na02f02 TIMEBOOST_cell_70515 ( .a(TIMEBOOST_net_22465), .b(g62776_sb), .o(n_5441) );
na02s01 g57965_u2 ( .a(FE_OFN555_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q), .o(g57965_db) );
na04m02 TIMEBOOST_cell_64841 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q), .b(TIMEBOOST_net_10389), .c(g64904_sb), .d(n_4450), .o(TIMEBOOST_net_8844) );
na02s01 TIMEBOOST_cell_62476 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_101), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_20185) );
na03f02 TIMEBOOST_cell_65891 ( .a(n_3972), .b(g62843_sb), .c(g62843_db), .o(n_5285) );
na02f02 TIMEBOOST_cell_37810 ( .a(FE_OFN223_n_9844), .b(g57927_sb), .o(TIMEBOOST_net_10517) );
na03m02 TIMEBOOST_cell_72702 ( .a(g65018_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q), .c(TIMEBOOST_net_14284), .o(TIMEBOOST_net_13234) );
na02f02 TIMEBOOST_cell_37811 ( .a(TIMEBOOST_net_10517), .b(g57927_db), .o(n_9882) );
in01s01 g57968_u0 ( .a(FE_OFN552_n_9864), .o(g57968_sb) );
na03m04 TIMEBOOST_cell_72842 ( .a(g65296_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q), .c(TIMEBOOST_net_14436), .o(TIMEBOOST_net_13376) );
na02s01 g57968_u2 ( .a(FE_OFN552_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q), .o(g57968_db) );
na02f02 TIMEBOOST_cell_51313 ( .a(n_7329), .b(n_14618), .o(TIMEBOOST_net_15874) );
in01s01 g57969_u0 ( .a(FE_OFN554_n_9864), .o(g57969_sb) );
na02m04 TIMEBOOST_cell_69887 ( .a(TIMEBOOST_net_22151), .b(g64213_sb), .o(TIMEBOOST_net_16972) );
na02m02 TIMEBOOST_cell_54035 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q), .o(TIMEBOOST_net_17235) );
in01s01 g57970_u0 ( .a(FE_OFN556_n_9864), .o(g57970_sb) );
na03f06 TIMEBOOST_cell_65402 ( .a(n_2922), .b(n_3004), .c(n_3079), .o(n_4145) );
na02s01 g57970_u2 ( .a(FE_OFN556_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q), .o(g57970_db) );
na02f02 TIMEBOOST_cell_54460 ( .a(TIMEBOOST_net_17447), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_15657) );
in01s01 g57971_u0 ( .a(FE_OFN551_n_9864), .o(g57971_sb) );
na03m02 TIMEBOOST_cell_66335 ( .a(n_1934), .b(g61741_sb), .c(g61741_db), .o(n_8335) );
in01s01 g57972_u0 ( .a(FE_OFN554_n_9864), .o(g57972_sb) );
na03f02 TIMEBOOST_cell_35020 ( .a(TIMEBOOST_net_9577), .b(FE_OFN2180_n_8567), .c(g57186_sb), .o(n_11566) );
in01s01 g57973_u0 ( .a(FE_OFN556_n_9864), .o(g57973_sb) );
na02s01 g57973_u2 ( .a(FE_OFN556_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q), .o(g57973_db) );
na02m02 TIMEBOOST_cell_44007 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q), .b(g65335_sb), .o(TIMEBOOST_net_12898) );
na03f02 TIMEBOOST_cell_66880 ( .a(FE_OFN1566_n_12502), .b(FE_OCPN1825_n_12030), .c(TIMEBOOST_net_13539), .o(n_12488) );
na03m04 TIMEBOOST_cell_69886 ( .a(TIMEBOOST_net_16616), .b(FE_OFN1051_n_16657), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q), .o(TIMEBOOST_net_22151) );
in01s02 g57975_u0 ( .a(FE_OFN554_n_9864), .o(g57975_sb) );
na02s03 TIMEBOOST_cell_53957 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q), .o(TIMEBOOST_net_17196) );
na03f02 TIMEBOOST_cell_73291 ( .a(n_3885), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q), .c(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_15183) );
na02s02 TIMEBOOST_cell_30655 ( .a(n_9410), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q), .o(TIMEBOOST_net_9432) );
na02s01 g57976_u2 ( .a(FE_OFN553_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q), .o(g57976_db) );
na02m01 TIMEBOOST_cell_54085 ( .a(n_4498), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q), .o(TIMEBOOST_net_17260) );
in01s01 g57977_u0 ( .a(FE_OFN532_n_9823), .o(g57977_sb) );
na03s02 TIMEBOOST_cell_67818 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q), .b(g65866_sb), .c(g65866_db), .o(n_1709) );
na02s01 TIMEBOOST_cell_63056 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q), .o(TIMEBOOST_net_20475) );
na02s02 TIMEBOOST_cell_63218 ( .a(FE_OFN1793_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q), .o(TIMEBOOST_net_20556) );
in01s01 g57978_u0 ( .a(FE_OFN535_n_9823), .o(g57978_sb) );
na02m02 TIMEBOOST_cell_69639 ( .a(TIMEBOOST_net_22027), .b(TIMEBOOST_net_10650), .o(TIMEBOOST_net_17004) );
in01s01 g57979_u0 ( .a(FE_OFN533_n_9823), .o(g57979_sb) );
na02m02 TIMEBOOST_cell_28315 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q), .b(g64302_sb), .o(TIMEBOOST_net_8262) );
na02s01 g57979_u2 ( .a(FE_OFN533_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q), .o(g57979_db) );
in01s01 g57980_u0 ( .a(FE_OFN1789_n_9823), .o(g57980_sb) );
na03s02 TIMEBOOST_cell_32075 ( .a(g58126_sb), .b(g58126_db), .c(FE_OFN270_n_9836), .o(n_9667) );
na02f20 TIMEBOOST_cell_54127 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_776), .o(TIMEBOOST_net_17281) );
in01s01 g57981_u0 ( .a(FE_OFN535_n_9823), .o(g57981_sb) );
na02s01 g57981_u2 ( .a(FE_OFN535_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q), .o(g57981_db) );
na02f02 TIMEBOOST_cell_70003 ( .a(TIMEBOOST_net_22209), .b(g61793_sb), .o(n_8213) );
in01s01 g57982_u0 ( .a(FE_OFN534_n_9823), .o(g57982_sb) );
na03m02 TIMEBOOST_cell_72653 ( .a(TIMEBOOST_net_21498), .b(g64836_sb), .c(TIMEBOOST_net_21673), .o(TIMEBOOST_net_17091) );
na02s01 g57982_u2 ( .a(FE_OFN534_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q), .o(g57982_db) );
in01s01 TIMEBOOST_cell_73877 ( .a(TIMEBOOST_net_23441), .o(TIMEBOOST_net_23442) );
in01s01 g57983_u0 ( .a(FE_OFN534_n_9823), .o(g57983_sb) );
in01s01 TIMEBOOST_cell_63562 ( .a(TIMEBOOST_net_20742), .o(wbs_adr_i_9_) );
na02s01 g57983_u2 ( .a(FE_OFN534_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q), .o(g57983_db) );
in01s01 g57984_u0 ( .a(FE_OFN531_n_9823), .o(g57984_sb) );
na02s01 g57984_u2 ( .a(FE_OFN531_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q), .o(g57984_db) );
na02f02 TIMEBOOST_cell_54508 ( .a(TIMEBOOST_net_17471), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_15353) );
in01m08 g57985_u0 ( .a(FE_OFN535_n_9823), .o(g57985_sb) );
in01s01 TIMEBOOST_cell_35500 ( .a(TIMEBOOST_net_10091), .o(wbs_dat_i_10_) );
na02m10 g57985_u2 ( .a(FE_OFN535_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q), .o(g57985_db) );
in01s01 TIMEBOOST_cell_35501 ( .a(TIMEBOOST_net_10092), .o(TIMEBOOST_net_10091) );
in01s01 g57986_u0 ( .a(FE_OFN533_n_9823), .o(g57986_sb) );
na02s02 TIMEBOOST_cell_49420 ( .a(TIMEBOOST_net_14927), .b(g58108_sb), .o(n_9685) );
na02f06 TIMEBOOST_cell_63683 ( .a(TIMEBOOST_net_20827), .b(n_2397), .o(n_2398) );
in01s01 g57987_u0 ( .a(FE_OFN531_n_9823), .o(g57987_sb) );
in01s01 TIMEBOOST_cell_35502 ( .a(TIMEBOOST_net_10093), .o(wbs_dat_i_22_) );
na02s02 g57987_u2 ( .a(FE_OFN531_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q), .o(g57987_db) );
in01s01 TIMEBOOST_cell_35503 ( .a(TIMEBOOST_net_10094), .o(TIMEBOOST_net_10093) );
in01s01 g57988_u0 ( .a(FE_OFN532_n_9823), .o(g57988_sb) );
in01s01 TIMEBOOST_cell_35504 ( .a(TIMEBOOST_net_10095), .o(TIMEBOOST_net_10074) );
in01s01 TIMEBOOST_cell_35505 ( .a(TIMEBOOST_net_10096), .o(TIMEBOOST_net_10095) );
in01s01 g57989_u0 ( .a(FE_OFN535_n_9823), .o(g57989_sb) );
na02s01 TIMEBOOST_cell_42960 ( .a(TIMEBOOST_net_12374), .b(FE_OFN953_n_2055), .o(TIMEBOOST_net_10534) );
na02s01 g57989_u2 ( .a(FE_OFN535_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q), .o(g57989_db) );
na03m04 TIMEBOOST_cell_73090 ( .a(g65397_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q), .c(TIMEBOOST_net_12757), .o(TIMEBOOST_net_17080) );
in01s02 g57990_u0 ( .a(FE_OFN531_n_9823), .o(g57990_sb) );
na02f02 TIMEBOOST_cell_70828 ( .a(TIMEBOOST_net_16691), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_22622) );
na03f02 TIMEBOOST_cell_46328 ( .a(TIMEBOOST_net_12496), .b(g64227_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q), .o(TIMEBOOST_net_13100) );
in01m08 g57991_u0 ( .a(FE_OFN535_n_9823), .o(g57991_sb) );
na03f01 TIMEBOOST_cell_68078 ( .a(pci_ad_i_27_), .b(n_574), .c(parchk_pci_ad_reg_in_1231), .o(TIMEBOOST_net_21247) );
na03s02 TIMEBOOST_cell_73500 ( .a(FE_OFN554_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q), .c(TIMEBOOST_net_12470), .o(TIMEBOOST_net_14324) );
in01s01 g57992_u0 ( .a(FE_OFN533_n_9823), .o(g57992_sb) );
in01s01 TIMEBOOST_cell_35506 ( .a(TIMEBOOST_net_10097), .o(TIMEBOOST_net_10080) );
na02s01 g57992_u2 ( .a(FE_OFN533_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q), .o(g57992_db) );
in01s01 TIMEBOOST_cell_35507 ( .a(TIMEBOOST_net_10098), .o(TIMEBOOST_net_10097) );
in01s01 g57993_u0 ( .a(FE_OFN533_n_9823), .o(g57993_sb) );
na02s01 TIMEBOOST_cell_30995 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_6__Q), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_9602) );
na02s01 g57993_u2 ( .a(FE_OFN533_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q), .o(g57993_db) );
na03f02 TIMEBOOST_cell_63444 ( .a(TIMEBOOST_net_13485), .b(FE_OCPN1888_FE_OFN473_n_16992), .c(n_15528), .o(TIMEBOOST_net_20669) );
in01s02 g57994_u0 ( .a(FE_OFN1789_n_9823), .o(g57994_sb) );
na02f02 TIMEBOOST_cell_63343 ( .a(TIMEBOOST_net_20618), .b(n_15695), .o(n_15698) );
na03f10 TIMEBOOST_cell_32076 ( .a(FE_RN_72_0), .b(FE_OCPN1854_n_2071), .c(FE_RN_73_0), .o(TIMEBOOST_net_694) );
in01s01 g57995_u0 ( .a(FE_OFN533_n_9823), .o(g57995_sb) );
na02s01 TIMEBOOST_cell_42962 ( .a(TIMEBOOST_net_12375), .b(FE_OFN951_n_2055), .o(TIMEBOOST_net_10535) );
na02s01 TIMEBOOST_cell_63755 ( .a(TIMEBOOST_net_20863), .b(FE_OFN235_n_9834), .o(TIMEBOOST_net_14678) );
na02s01 TIMEBOOST_cell_54169 ( .a(FE_OFN258_n_9862), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q), .o(TIMEBOOST_net_17302) );
in01s01 g57996_u0 ( .a(FE_OFN535_n_9823), .o(g57996_sb) );
in01s01 TIMEBOOST_cell_35508 ( .a(TIMEBOOST_net_10099), .o(TIMEBOOST_net_10084) );
na02s01 g57996_u2 ( .a(FE_OFN535_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q), .o(g57996_db) );
in01s01 TIMEBOOST_cell_35509 ( .a(TIMEBOOST_net_10100), .o(TIMEBOOST_net_10099) );
in01s01 g57997_u0 ( .a(FE_OFN535_n_9823), .o(g57997_sb) );
na02s01 g57997_u2 ( .a(FE_OFN535_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q), .o(g57997_db) );
na03s02 TIMEBOOST_cell_46429 ( .a(TIMEBOOST_net_12428), .b(FE_OFN563_n_9895), .c(g57921_sb), .o(n_9890) );
na02m02 TIMEBOOST_cell_71396 ( .a(n_2017), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_22906) );
na02s01 g57998_u2 ( .a(FE_OFN1789_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q), .o(g57998_db) );
na03f08 TIMEBOOST_cell_32077 ( .a(n_16451), .b(FE_OCPN1875_n_14526), .c(n_16452), .o(n_16455) );
in01s01 g57999_u0 ( .a(FE_OFN531_n_9823), .o(g57999_sb) );
na04f04 TIMEBOOST_cell_73292 ( .a(TIMEBOOST_net_16968), .b(g52630_sb), .c(TIMEBOOST_net_11642), .d(n_14839), .o(TIMEBOOST_net_22794) );
na03f02 TIMEBOOST_cell_73539 ( .a(TIMEBOOST_net_17508), .b(FE_OFN1232_n_6391), .c(g62570_sb), .o(n_6415) );
no02f02 g57_u0 ( .a(n_15585), .b(n_15562), .o(n_15586) );
in01s01 g58000_u0 ( .a(FE_OFN534_n_9823), .o(g58000_sb) );
na02s01 g58000_u2 ( .a(FE_OFN534_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q), .o(g58000_db) );
na02m02 TIMEBOOST_cell_71238 ( .a(TIMEBOOST_net_7619), .b(g53945_da), .o(TIMEBOOST_net_22827) );
in01s02 g58001_u0 ( .a(FE_OFN533_n_9823), .o(g58001_sb) );
in01s01 TIMEBOOST_cell_35510 ( .a(TIMEBOOST_net_10101), .o(TIMEBOOST_net_10086) );
in01s01 TIMEBOOST_cell_35511 ( .a(TIMEBOOST_net_10102), .o(TIMEBOOST_net_10101) );
in01s01 g58002_u0 ( .a(FE_OFN531_n_9823), .o(g58002_sb) );
na02s01 TIMEBOOST_cell_42803 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q), .o(TIMEBOOST_net_12296) );
na02s01 TIMEBOOST_cell_30997 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_9603) );
in01s01 g58003_u0 ( .a(FE_OFN534_n_9823), .o(g58003_sb) );
na02f04 TIMEBOOST_cell_72211 ( .a(TIMEBOOST_net_23313), .b(g54239_db), .o(TIMEBOOST_net_13509) );
na02s01 g58003_u2 ( .a(FE_OFN534_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q), .o(g58003_db) );
in01s01 TIMEBOOST_cell_45995 ( .a(TIMEBOOST_net_13956), .o(TIMEBOOST_net_13897) );
in01s01 g58004_u0 ( .a(FE_OFN1789_n_9823), .o(g58004_sb) );
na02f02 TIMEBOOST_cell_70653 ( .a(TIMEBOOST_net_22534), .b(g63143_sb), .o(n_4961) );
na03s06 TIMEBOOST_cell_73071 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q), .b(FE_OFN702_n_7845), .c(TIMEBOOST_net_22259), .o(TIMEBOOST_net_14763) );
in01s01 g58005_u0 ( .a(FE_OFN1789_n_9823), .o(g58005_sb) );
na03f02 TIMEBOOST_cell_65839 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(g64078_sb), .c(g64078_db), .o(n_4077) );
na03f02 TIMEBOOST_cell_66445 ( .a(TIMEBOOST_net_17126), .b(FE_OFN1315_n_6624), .c(g62947_sb), .o(n_5987) );
in01s01 g58006_u0 ( .a(FE_OFN533_n_9823), .o(g58006_sb) );
na02s01 g58006_u2 ( .a(FE_OFN533_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q), .o(g58006_db) );
na02m10 TIMEBOOST_cell_54281 ( .a(configuration_pci_err_data_511), .b(wbm_dat_o_10_), .o(TIMEBOOST_net_17358) );
na03f02 TIMEBOOST_cell_73540 ( .a(TIMEBOOST_net_17069), .b(FE_OFN1231_n_6391), .c(g62378_sb), .o(n_6847) );
in01s01 g58008_u0 ( .a(FE_OFN529_n_9899), .o(g58008_sb) );
na04m02 TIMEBOOST_cell_64994 ( .a(n_4452), .b(g65003_sb), .c(g65003_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q), .o(TIMEBOOST_net_17429) );
in01m04 g58009_u0 ( .a(FE_OFN527_n_9899), .o(g58009_sb) );
in01s01 TIMEBOOST_cell_35512 ( .a(TIMEBOOST_net_10103), .o(TIMEBOOST_net_10088) );
na02m08 g58009_u2 ( .a(FE_OFN527_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q), .o(g58009_db) );
in01s01 TIMEBOOST_cell_35513 ( .a(TIMEBOOST_net_10104), .o(TIMEBOOST_net_10103) );
in01s01 g58010_u0 ( .a(FE_OFN527_n_9899), .o(g58010_sb) );
na02s01 g58010_u2 ( .a(FE_OFN527_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q), .o(g58010_db) );
in01s01 g58011_u0 ( .a(FE_OFN525_n_9899), .o(g58011_sb) );
na02s02 TIMEBOOST_cell_63064 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q), .o(TIMEBOOST_net_20479) );
na02f02 TIMEBOOST_cell_49640 ( .a(TIMEBOOST_net_15037), .b(g61778_sb), .o(n_8251) );
in01s01 g58012_u0 ( .a(FE_OFN527_n_9899), .o(g58012_sb) );
na02f02 TIMEBOOST_cell_62447 ( .a(TIMEBOOST_net_20170), .b(TIMEBOOST_net_10284), .o(n_2568) );
na02s02 TIMEBOOST_cell_48724 ( .a(TIMEBOOST_net_14579), .b(TIMEBOOST_net_10464), .o(TIMEBOOST_net_9548) );
na02s02 TIMEBOOST_cell_38271 ( .a(g57909_db), .b(TIMEBOOST_net_10747), .o(n_9906) );
in01s01 g58013_u0 ( .a(FE_OFN528_n_9899), .o(g58013_sb) );
na02s01 g58013_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN528_n_9899), .o(g58013_db) );
in01s01 g58014_u0 ( .a(FE_OFN528_n_9899), .o(g58014_sb) );
na02s01 g58014_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q), .b(FE_OFN528_n_9899), .o(g58014_db) );
na03s02 TIMEBOOST_cell_46381 ( .a(TIMEBOOST_net_12460), .b(g58257_sb), .c(TIMEBOOST_net_12702), .o(TIMEBOOST_net_9562) );
in01s01 g58015_u0 ( .a(FE_OFN529_n_9899), .o(g58015_sb) );
na04f04 TIMEBOOST_cell_36831 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q), .b(FE_OFN1389_n_8567), .c(n_9647), .d(g57285_sb), .o(n_11468) );
na02s01 g58015_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q), .b(FE_OFN529_n_9899), .o(g58015_db) );
in01s01 g58016_u0 ( .a(FE_OFN526_n_9899), .o(g58016_sb) );
na02s02 TIMEBOOST_cell_52906 ( .a(TIMEBOOST_net_16670), .b(g58214_db), .o(TIMEBOOST_net_9404) );
na02f01 TIMEBOOST_cell_70652 ( .a(TIMEBOOST_net_15057), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_22534) );
na03f08 TIMEBOOST_cell_31959 ( .a(n_1325), .b(n_15371), .c(n_7568), .o(TIMEBOOST_net_422) );
in01m10 g58017_u0 ( .a(FE_OFN527_n_9899), .o(g58017_sb) );
na02f02 TIMEBOOST_cell_70202 ( .a(TIMEBOOST_net_14751), .b(FE_OFN2128_n_16497), .o(TIMEBOOST_net_22309) );
na02m02 TIMEBOOST_cell_53580 ( .a(TIMEBOOST_net_17007), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_15320) );
in01s01 g58018_u0 ( .a(FE_OFN526_n_9899), .o(g58018_sb) );
na02m02 TIMEBOOST_cell_28335 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(g65797_sb), .o(TIMEBOOST_net_8272) );
na02s01 g58018_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q), .b(FE_OFN526_n_9899), .o(g58018_db) );
na02m02 TIMEBOOST_cell_69098 ( .a(FE_OFN1642_n_4671), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q), .o(TIMEBOOST_net_21757) );
in01s01 g58019_u0 ( .a(FE_OFN529_n_9899), .o(g58019_sb) );
na04f04 TIMEBOOST_cell_65466 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_513), .c(n_16429), .d(n_15731), .o(n_15732) );
na02s01 g58019_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q), .b(FE_OFN529_n_9899), .o(g58019_db) );
na03f02 TIMEBOOST_cell_34919 ( .a(TIMEBOOST_net_9453), .b(FE_OFN1382_n_8567), .c(g57240_sb), .o(n_10426) );
in01s01 g58020_u0 ( .a(FE_OFN527_n_9899), .o(g58020_sb) );
na03f02 TIMEBOOST_cell_73541 ( .a(TIMEBOOST_net_17505), .b(FE_OFN1231_n_6391), .c(g62688_sb), .o(n_6166) );
na02s01 g58020_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q), .b(FE_OFN527_n_9899), .o(g58020_db) );
na03f02 TIMEBOOST_cell_73542 ( .a(TIMEBOOST_net_17557), .b(FE_OFN1231_n_6391), .c(g62337_sb), .o(n_6924) );
in01s01 g58021_u0 ( .a(FE_OFN525_n_9899), .o(g58021_sb) );
na03f02 TIMEBOOST_cell_73794 ( .a(TIMEBOOST_net_13751), .b(FE_OFN1599_n_13995), .c(FE_OFN1605_n_13997), .o(n_14444) );
na02s01 TIMEBOOST_cell_45239 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q), .o(TIMEBOOST_net_13514) );
in01m08 g58022_u0 ( .a(FE_OFN527_n_9899), .o(g58022_sb) );
na02m02 TIMEBOOST_cell_68787 ( .a(TIMEBOOST_net_21601), .b(g64334_sb), .o(n_3843) );
na02f01 TIMEBOOST_cell_48726 ( .a(TIMEBOOST_net_14580), .b(FE_OFN1051_n_16657), .o(TIMEBOOST_net_10976) );
in01s01 g58023_u0 ( .a(FE_OFN527_n_9899), .o(g58023_sb) );
na03m06 TIMEBOOST_cell_72844 ( .a(g64166_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q), .c(TIMEBOOST_net_12541), .o(TIMEBOOST_net_8322) );
na02s01 g58023_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q), .b(FE_OFN527_n_9899), .o(g58023_db) );
in01s01 g58024_u0 ( .a(FE_OFN525_n_9899), .o(g58024_sb) );
na03f02 TIMEBOOST_cell_64585 ( .a(n_2206), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q), .c(FE_OFN1812_n_7845), .o(TIMEBOOST_net_15101) );
na02f01 TIMEBOOST_cell_49348 ( .a(TIMEBOOST_net_14891), .b(FE_OFN1095_g64577_p), .o(TIMEBOOST_net_12955) );
in01s01 g58025_u0 ( .a(FE_OFN527_n_9899), .o(g58025_sb) );
no03f04 TIMEBOOST_cell_73682 ( .a(n_4652), .b(n_12595), .c(n_4879), .o(g59345_p) );
na02s01 TIMEBOOST_cell_42961 ( .a(pci_target_unit_fifos_pcir_data_in), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q), .o(TIMEBOOST_net_12375) );
na02s02 TIMEBOOST_cell_37845 ( .a(TIMEBOOST_net_10534), .b(g65726_sb), .o(n_1938) );
in01s01 g58026_u0 ( .a(FE_OFN527_n_9899), .o(g58026_sb) );
na02s02 TIMEBOOST_cell_37847 ( .a(TIMEBOOST_net_10535), .b(g65696_sb), .o(n_1950) );
in01s01 g58027_u0 ( .a(FE_OFN528_n_9899), .o(g58027_sb) );
na03f02 TIMEBOOST_cell_34915 ( .a(TIMEBOOST_net_9560), .b(FE_OFN1411_n_8567), .c(g57507_sb), .o(n_10325) );
na02s01 g58027_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q), .b(FE_OFN528_n_9899), .o(g58027_db) );
in01m06 g58028_u0 ( .a(FE_OFN527_n_9899), .o(g58028_sb) );
na02m02 TIMEBOOST_cell_68850 ( .a(n_4476), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q), .o(TIMEBOOST_net_21633) );
na02m10 g58028_u2 ( .a(FE_OFN527_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q), .o(g58028_db) );
in01s01 g58029_u0 ( .a(FE_OFN525_n_9899), .o(g58029_sb) );
na02s01 TIMEBOOST_cell_63016 ( .a(g62007_sb), .b(g62007_db), .o(TIMEBOOST_net_20455) );
na02s01 TIMEBOOST_cell_42959 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q), .o(TIMEBOOST_net_12374) );
na03f02 TIMEBOOST_cell_73436 ( .a(TIMEBOOST_net_20539), .b(FE_OFN1288_n_4098), .c(g62884_sb), .o(n_6109) );
in01s01 g58030_u0 ( .a(FE_OFN526_n_9899), .o(g58030_sb) );
na03f02 TIMEBOOST_cell_73543 ( .a(TIMEBOOST_net_20582), .b(FE_OFN1236_n_6391), .c(g62977_sb), .o(n_5928) );
na02m02 TIMEBOOST_cell_48638 ( .a(TIMEBOOST_net_14536), .b(g65238_sb), .o(n_2645) );
in01s01 g58031_u0 ( .a(FE_OFN528_n_9899), .o(g58031_sb) );
na02m01 g64944_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q), .b(FE_OFN649_n_4497), .o(g64944_db) );
na03f02 TIMEBOOST_cell_73501 ( .a(TIMEBOOST_net_8846), .b(FE_OFN1166_n_5615), .c(g61676_sb), .o(n_4891) );
na02s01 TIMEBOOST_cell_38451 ( .a(TIMEBOOST_net_10837), .b(g58099_db), .o(n_9701) );
in01s01 g58032_u0 ( .a(FE_OFN526_n_9899), .o(g58032_sb) );
na02s01 TIMEBOOST_cell_28341 ( .a(configuration_wb_err_data_594), .b(parchk_pci_ad_out_in_1191), .o(TIMEBOOST_net_8275) );
na02s02 g58032_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q), .b(FE_OFN526_n_9899), .o(g58032_db) );
na03m02 TIMEBOOST_cell_72596 ( .a(n_3783), .b(FE_OFN652_n_4508), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q), .o(TIMEBOOST_net_22027) );
in01s01 g58033_u0 ( .a(FE_OFN526_n_9899), .o(g58033_sb) );
na03m02 TIMEBOOST_cell_65403 ( .a(wbs_sel_i_2_), .b(g63586_sb), .c(g63586_db), .o(n_4102) );
na02s01 g58033_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q), .b(FE_OFN526_n_9899), .o(g58033_db) );
na02f01 TIMEBOOST_cell_52395 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_16415) );
in01s01 g58034_u0 ( .a(FE_OFN528_n_9899), .o(g58034_sb) );
na02s01 g58034_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q), .b(FE_OFN528_n_9899), .o(g58034_db) );
na02s01 TIMEBOOST_cell_30971 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_24__Q), .b(FE_OFN227_n_9841), .o(TIMEBOOST_net_9590) );
in01s01 g58035_u0 ( .a(FE_OFN525_n_9899), .o(g58035_sb) );
na02s01 TIMEBOOST_cell_49454 ( .a(TIMEBOOST_net_14944), .b(FE_OFN596_n_9694), .o(TIMEBOOST_net_12991) );
na02m06 TIMEBOOST_cell_72222 ( .a(TIMEBOOST_net_10052), .b(configuration_wb_err_addr_544), .o(TIMEBOOST_net_23319) );
in01s01 g58036_u0 ( .a(FE_OFN525_n_9899), .o(g58036_sb) );
na02m02 TIMEBOOST_cell_69135 ( .a(TIMEBOOST_net_21775), .b(TIMEBOOST_net_12735), .o(TIMEBOOST_net_17564) );
na02f02 TIMEBOOST_cell_50676 ( .a(TIMEBOOST_net_15555), .b(TIMEBOOST_net_11526), .o(TIMEBOOST_net_9457) );
in01s01 g58037_u0 ( .a(FE_OFN528_n_9899), .o(g58037_sb) );
na02m01 TIMEBOOST_cell_53912 ( .a(TIMEBOOST_net_17173), .b(TIMEBOOST_net_12991), .o(TIMEBOOST_net_9400) );
na02s01 g58037_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN528_n_9899), .o(g58037_db) );
na02s01 TIMEBOOST_cell_38401 ( .a(TIMEBOOST_net_10812), .b(g58233_db), .o(n_9046) );
na02s01 g58038_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN527_n_9899), .o(g58038_db) );
na02m02 TIMEBOOST_cell_72006 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q), .o(TIMEBOOST_net_23211) );
in01s01 g58039_u0 ( .a(FE_OFN606_n_9904), .o(g58039_sb) );
na03f02 TIMEBOOST_cell_73368 ( .a(TIMEBOOST_net_16718), .b(FE_OFN1299_n_5763), .c(g62046_sb), .o(n_7766) );
na02s01 g58039_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q), .b(FE_OFN606_n_9904), .o(g58039_db) );
na02s01 TIMEBOOST_cell_52615 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_16525) );
in01s01 g58040_u0 ( .a(FE_OFN606_n_9904), .o(g58040_sb) );
na02s01 TIMEBOOST_cell_28343 ( .a(configuration_wb_err_data_572), .b(parchk_pci_ad_out_in_1169), .o(TIMEBOOST_net_8276) );
na02s01 g58040_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q), .b(FE_OFN606_n_9904), .o(g58040_db) );
in01s01 g58041_u0 ( .a(FE_OFN608_n_9904), .o(g58041_sb) );
na02m01 TIMEBOOST_cell_28345 ( .a(configuration_wb_err_data_593), .b(parchk_pci_ad_out_in_1190), .o(TIMEBOOST_net_8277) );
na02s01 g58041_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q), .b(FE_OFN608_n_9904), .o(g58041_db) );
in01s01 g58042_u0 ( .a(n_9904), .o(g58042_sb) );
na02s01 TIMEBOOST_cell_47770 ( .a(TIMEBOOST_net_14102), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_12380) );
in01s02 TIMEBOOST_cell_67798 ( .a(TIMEBOOST_net_21225), .o(TIMEBOOST_net_21224) );
in01m06 g58043_u0 ( .a(FE_OFN1794_n_9904), .o(g58043_sb) );
na04f02 TIMEBOOST_cell_73502 ( .a(n_2178), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q), .c(FE_OFN2212_n_8407), .d(g62018_sb), .o(n_7859) );
na02m08 g58043_u2 ( .a(FE_OFN1794_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q), .o(g58043_db) );
na02f02 TIMEBOOST_cell_70667 ( .a(TIMEBOOST_net_22541), .b(g63188_sb), .o(n_4943) );
in01s01 g58044_u0 ( .a(FE_OFN606_n_9904), .o(g58044_sb) );
na02m01 TIMEBOOST_cell_51859 ( .a(g64810_sb), .b(n_3747), .o(TIMEBOOST_net_16147) );
na02s01 g58044_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q), .b(FE_OFN606_n_9904), .o(g58044_db) );
in01s01 g58045_u0 ( .a(FE_OFN606_n_9904), .o(g58045_sb) );
na02s01 g58045_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q), .b(FE_OFN606_n_9904), .o(g58045_db) );
na03f02 TIMEBOOST_cell_66292 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q), .b(g63198_sb), .c(g63198_db), .o(n_5768) );
in01s01 g58046_u0 ( .a(FE_OFN608_n_9904), .o(g58046_sb) );
na02s01 g58046_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q), .b(FE_OFN608_n_9904), .o(g58046_db) );
in01s01 TIMEBOOST_cell_67757 ( .a(pci_target_unit_fifos_pcir_data_in_164), .o(TIMEBOOST_net_21184) );
in01s01 g58047_u0 ( .a(FE_OFN1793_n_9904), .o(g58047_sb) );
na02s01 TIMEBOOST_cell_28347 ( .a(configuration_wb_err_cs_bit_564), .b(conf_wb_err_bc_in_846), .o(TIMEBOOST_net_8278) );
na03f02 TIMEBOOST_cell_34942 ( .a(TIMEBOOST_net_9536), .b(FE_OFN1399_n_8567), .c(g57252_sb), .o(n_11503) );
na02s01 TIMEBOOST_cell_53959 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q), .o(TIMEBOOST_net_17197) );
in01s01 g58048_u0 ( .a(FE_OFN1795_n_9904), .o(g58048_sb) );
na02s02 g58048_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q), .b(FE_OFN1795_n_9904), .o(g58048_db) );
na02m01 TIMEBOOST_cell_53365 ( .a(TIMEBOOST_net_12408), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_16900) );
in01s01 g58049_u0 ( .a(FE_OFN606_n_9904), .o(g58049_sb) );
na03f01 TIMEBOOST_cell_68226 ( .a(n_2651), .b(n_1847), .c(FE_OFN989_n_574), .o(TIMEBOOST_net_21321) );
na02s01 g58049_u2 ( .a(FE_OFN606_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q), .o(g58049_db) );
na02s01 TIMEBOOST_cell_43687 ( .a(FE_OFN1789_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q), .o(TIMEBOOST_net_12738) );
in01s01 g58050_u0 ( .a(FE_OFN606_n_9904), .o(g58050_sb) );
na02s01 g58050_u2 ( .a(FE_OFN606_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q), .o(g58050_db) );
in01s01 g58051_u0 ( .a(FE_OFN607_n_9904), .o(g58051_sb) );
na02m01 TIMEBOOST_cell_68558 ( .a(FE_OFN624_n_4409), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q), .o(TIMEBOOST_net_21487) );
na02s01 g58051_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q), .b(FE_OFN607_n_9904), .o(g58051_db) );
na02s01 TIMEBOOST_cell_31085 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_9647) );
in01s01 g58052_u0 ( .a(FE_OFN1794_n_9904), .o(g58052_sb) );
na02f02 TIMEBOOST_cell_54372 ( .a(TIMEBOOST_net_17403), .b(FE_OFN1214_n_4151), .o(TIMEBOOST_net_15341) );
na02m02 TIMEBOOST_cell_70171 ( .a(TIMEBOOST_net_22293), .b(g64081_sb), .o(n_4074) );
in01s01 g58053_u0 ( .a(FE_OFN1793_n_9904), .o(g58053_sb) );
na02s01 g58054_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q), .b(n_9904), .o(g58054_db) );
na03f02 TIMEBOOST_cell_73452 ( .a(TIMEBOOST_net_17378), .b(FE_OFN1248_n_4093), .c(g62907_sb), .o(n_6063) );
in01s01 g58055_u0 ( .a(FE_OFN1793_n_9904), .o(g58055_sb) );
na03m02 TIMEBOOST_cell_65044 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q), .b(TIMEBOOST_net_9793), .c(g64351_sb), .o(n_3827) );
in01s01 g58056_u0 ( .a(FE_OFN606_n_9904), .o(g58056_sb) );
na02s01 TIMEBOOST_cell_49279 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q), .b(FE_OFN602_n_9687), .o(TIMEBOOST_net_14857) );
na02s01 g58056_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q), .b(FE_OFN606_n_9904), .o(g58056_db) );
in01s01 g58057_u0 ( .a(FE_OFN1794_n_9904), .o(g58057_sb) );
na02f01 TIMEBOOST_cell_68051 ( .a(TIMEBOOST_net_21233), .b(wbu_addr_in_255), .o(TIMEBOOST_net_12309) );
na02s01 g58057_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q), .b(FE_OFN1794_n_9904), .o(g58057_db) );
na03s02 TIMEBOOST_cell_67873 ( .a(TIMEBOOST_net_21199), .b(g65754_sb), .c(g65754_db), .o(n_1921) );
in01s01 g58058_u0 ( .a(FE_OFN607_n_9904), .o(g58058_sb) );
na03f02 TIMEBOOST_cell_47039 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_12__Q), .b(n_13221), .c(FE_OFN2070_n_15978), .o(TIMEBOOST_net_11764) );
na02s01 g58058_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q), .b(FE_OFN607_n_9904), .o(g58058_db) );
na02m01 TIMEBOOST_cell_62634 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_146), .o(TIMEBOOST_net_20264) );
in01s01 g58059_u0 ( .a(FE_OFN1795_n_9904), .o(g58059_sb) );
na03f01 TIMEBOOST_cell_47372 ( .a(FE_OFN1583_n_12306), .b(TIMEBOOST_net_13689), .c(FE_OFN1760_n_10780), .o(n_12741) );
na03f02 TIMEBOOST_cell_34944 ( .a(TIMEBOOST_net_9454), .b(FE_OFN1391_n_8567), .c(g57236_sb), .o(n_10432) );
in01s01 g58060_u0 ( .a(FE_OFN606_n_9904), .o(g58060_sb) );
na02f02 TIMEBOOST_cell_47592 ( .a(TIMEBOOST_net_14013), .b(n_2214), .o(TIMEBOOST_net_85) );
na03f02 TIMEBOOST_cell_47373 ( .a(FE_OFN1584_n_12306), .b(TIMEBOOST_net_13690), .c(FE_OFN1761_n_10780), .o(n_12514) );
na02s01 g58061_u2 ( .a(FE_OFN608_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q), .o(g58061_db) );
na02m06 TIMEBOOST_cell_69239 ( .a(TIMEBOOST_net_21827), .b(n_4465), .o(TIMEBOOST_net_20367) );
in01s02 g58062_u0 ( .a(FE_OFN1795_n_9904), .o(g58062_sb) );
na02s01 g58062_u2 ( .a(FE_OFN1795_n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q), .o(g58062_db) );
in01s01 g58063_u0 ( .a(FE_OFN606_n_9904), .o(g58063_sb) );
na03f02 TIMEBOOST_cell_73180 ( .a(TIMEBOOST_net_16950), .b(FE_OFN1150_n_13249), .c(g54132_sb), .o(n_13467) );
na02s01 g58063_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q), .b(FE_OFN606_n_9904), .o(g58063_db) );
na02f01 TIMEBOOST_cell_39480 ( .a(TIMEBOOST_net_8325), .b(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_11352) );
na02f02 TIMEBOOST_cell_50486 ( .a(TIMEBOOST_net_15460), .b(g62984_sb), .o(n_5914) );
na02s01 g58064_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q), .b(FE_OFN607_n_9904), .o(g58064_db) );
na02s04 TIMEBOOST_cell_43471 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q), .b(g65919_sb), .o(TIMEBOOST_net_12630) );
na02f01 TIMEBOOST_cell_53044 ( .a(TIMEBOOST_net_16739), .b(FE_OFN1180_n_3476), .o(TIMEBOOST_net_15301) );
na02f02 TIMEBOOST_cell_49810 ( .a(TIMEBOOST_net_15122), .b(g62810_sb), .o(n_5358) );
in01s01 g58066_u0 ( .a(FE_OFN606_n_9904), .o(g58066_sb) );
na02s01 g58066_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q), .b(FE_OFN606_n_9904), .o(g58066_db) );
in01s01 TIMEBOOST_cell_63539 ( .a(TIMEBOOST_net_20719), .o(TIMEBOOST_net_20718) );
na02m01 g67069_u2 ( .a(pci_ad_i_12_), .b(n_574), .o(g67069_db) );
na02s01 g58067_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q), .b(FE_OFN608_n_9904), .o(g58067_db) );
na03f02 TIMEBOOST_cell_70646 ( .a(n_4037), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q), .c(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_22531) );
in01s01 g58068_u0 ( .a(FE_OFN1793_n_9904), .o(g58068_sb) );
na02s01 TIMEBOOST_cell_63132 ( .a(FE_OFN551_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q), .o(TIMEBOOST_net_20513) );
na04s02 TIMEBOOST_cell_73091 ( .a(TIMEBOOST_net_10784), .b(g65832_sb), .c(g61897_sb), .d(g61897_db), .o(n_8032) );
na02f01 TIMEBOOST_cell_42982 ( .a(FE_OFN918_n_4725), .b(TIMEBOOST_net_12385), .o(TIMEBOOST_net_10448) );
in01m02 g58069_u0 ( .a(FE_OFN576_n_9902), .o(g58069_sb) );
na02m02 TIMEBOOST_cell_49428 ( .a(TIMEBOOST_net_14931), .b(g57910_sb), .o(TIMEBOOST_net_12977) );
na03f02 TIMEBOOST_cell_66339 ( .a(TIMEBOOST_net_21009), .b(FE_OFN1232_n_6391), .c(g62355_sb), .o(n_6889) );
in01s01 g58070_u0 ( .a(FE_OFN577_n_9902), .o(g58070_sb) );
na02s01 TIMEBOOST_cell_45383 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q), .o(TIMEBOOST_net_13586) );
in01s01 TIMEBOOST_cell_73993 ( .a(TIMEBOOST_net_23557), .o(TIMEBOOST_net_23558) );
in01m02 g58071_u0 ( .a(FE_OFN575_n_9902), .o(g58071_sb) );
na03m02 TIMEBOOST_cell_72591 ( .a(TIMEBOOST_net_21437), .b(g65020_sb), .c(TIMEBOOST_net_21667), .o(TIMEBOOST_net_17421) );
na02s01 g58071_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q), .b(FE_OFN575_n_9902), .o(g58071_db) );
in01s01 g58072_u0 ( .a(FE_OFN574_n_9902), .o(g58072_sb) );
na02s04 TIMEBOOST_cell_68124 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_87), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_21270) );
na03m08 TIMEBOOST_cell_65116 ( .a(n_3777), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q), .c(FE_OFN666_n_4495), .o(TIMEBOOST_net_14397) );
in01s01 g58073_u0 ( .a(FE_OFN577_n_9902), .o(g58073_sb) );
na02m10 TIMEBOOST_cell_52973 ( .a(wishbone_slave_unit_pcim_sm_data_in_643), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q), .o(TIMEBOOST_net_16704) );
na03m04 TIMEBOOST_cell_72820 ( .a(g64753_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q), .c(TIMEBOOST_net_10615), .o(TIMEBOOST_net_17362) );
in01s01 g58074_u0 ( .a(FE_OFN576_n_9902), .o(g58074_sb) );
na02s01 TIMEBOOST_cell_68052 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_71), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_21234) );
na02s01 g58074_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q), .b(FE_OFN576_n_9902), .o(g58074_db) );
in01m01 g58075_u0 ( .a(FE_OFN576_n_9902), .o(g58075_sb) );
na02s01 TIMEBOOST_cell_49429 ( .a(FE_OFN1648_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q), .o(TIMEBOOST_net_14932) );
na02m10 TIMEBOOST_cell_45385 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q), .o(TIMEBOOST_net_13587) );
na03m02 TIMEBOOST_cell_65257 ( .a(TIMEBOOST_net_14479), .b(g64274_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q), .o(TIMEBOOST_net_15063) );
in01s01 g58076_u0 ( .a(FE_OFN577_n_9902), .o(g58076_sb) );
na02f02 TIMEBOOST_cell_62967 ( .a(TIMEBOOST_net_20430), .b(g54157_sb), .o(FE_RN_213_0) );
na02s01 g58076_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q), .b(FE_OFN577_n_9902), .o(g58076_db) );
in01s01 g58077_u0 ( .a(FE_OFN575_n_9902), .o(g58077_sb) );
na02m02 TIMEBOOST_cell_53378 ( .a(TIMEBOOST_net_16906), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_14521) );
na02s01 g58077_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q), .b(FE_OFN575_n_9902), .o(g58077_db) );
na02s02 TIMEBOOST_cell_70471 ( .a(TIMEBOOST_net_22443), .b(g58205_sb), .o(n_9582) );
in01m01 g58078_u0 ( .a(FE_OFN577_n_9902), .o(g58078_sb) );
na03f02 TIMEBOOST_cell_72527 ( .a(TIMEBOOST_net_21393), .b(g64141_sb), .c(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_22489) );
na02s01 g58078_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q), .b(FE_OFN577_n_9902), .o(g58078_db) );
na02m02 TIMEBOOST_cell_68852 ( .a(FE_OFN647_n_4497), .b(n_4343), .o(TIMEBOOST_net_21634) );
in01m02 g58079_u0 ( .a(FE_OFN577_n_9902), .o(g58079_sb) );
na02m02 TIMEBOOST_cell_28367 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q), .b(g65356_sb), .o(TIMEBOOST_net_8288) );
in01s01 TIMEBOOST_cell_67800 ( .a(TIMEBOOST_net_21227), .o(TIMEBOOST_net_21226) );
na03f02 TIMEBOOST_cell_66289 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q), .b(g62516_sb), .c(g62516_db), .o(n_6546) );
in01s01 g58080_u0 ( .a(FE_OFN577_n_9902), .o(g58080_sb) );
na02s01 g58080_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q), .b(FE_OFN577_n_9902), .o(g58080_db) );
in01s01 TIMEBOOST_cell_72357 ( .a(TIMEBOOST_net_23389), .o(TIMEBOOST_net_23390) );
in01f02 g58081_u0 ( .a(FE_OFN574_n_9902), .o(g58081_sb) );
na02m02 g58081_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q), .b(FE_OFN574_n_9902), .o(g58081_db) );
na02m02 TIMEBOOST_cell_49326 ( .a(TIMEBOOST_net_14880), .b(g64149_sb), .o(TIMEBOOST_net_8783) );
in01m01 g58082_u0 ( .a(FE_OFN577_n_9902), .o(g58082_sb) );
na04m02 TIMEBOOST_cell_67303 ( .a(TIMEBOOST_net_10489), .b(n_4488), .c(g64842_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q), .o(TIMEBOOST_net_17536) );
na02s01 g58082_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q), .b(FE_OFN577_n_9902), .o(g58082_db) );
na02f01 TIMEBOOST_cell_70348 ( .a(TIMEBOOST_net_17292), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_22382) );
in01s01 g58083_u0 ( .a(FE_OFN575_n_9902), .o(g58083_sb) );
na02s01 TIMEBOOST_cell_28369 ( .a(g61705_sb), .b(g61776_db), .o(TIMEBOOST_net_8289) );
na02s01 g58083_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q), .b(FE_OFN575_n_9902), .o(g58083_db) );
na02s01 TIMEBOOST_cell_49475 ( .a(g57929_sb), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_14955) );
in01s01 g58084_u0 ( .a(FE_OFN575_n_9902), .o(g58084_sb) );
na02s01 g58084_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q), .b(FE_OFN575_n_9902), .o(g58084_db) );
na02s01 TIMEBOOST_cell_47535 ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .b(wishbone_slave_unit_delayed_write_data_comp_wdata_out_76), .o(TIMEBOOST_net_13985) );
na02s01 g58085_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q), .b(FE_OFN574_n_9902), .o(g58085_db) );
na02m10 TIMEBOOST_cell_43945 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61), .b(pci_target_unit_pcit_if_strd_addr_in_697), .o(TIMEBOOST_net_12867) );
in01m01 g58086_u0 ( .a(FE_OFN575_n_9902), .o(g58086_sb) );
na02s01 TIMEBOOST_cell_49446 ( .a(TIMEBOOST_net_14940), .b(FE_OFN600_n_9687), .o(TIMEBOOST_net_12987) );
na04f04 TIMEBOOST_cell_42465 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q), .b(n_13168), .c(FE_OFN1327_n_13547), .d(g53923_sb), .o(n_13521) );
na02s02 TIMEBOOST_cell_28333 ( .a(TIMEBOOST_net_21159), .b(g65788_sb), .o(TIMEBOOST_net_8271) );
in01m01 g58087_u0 ( .a(FE_OFN577_n_9902), .o(g58087_sb) );
na02f02 TIMEBOOST_cell_38670 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q), .b(g64237_sb), .o(TIMEBOOST_net_10947) );
na02s01 g58087_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q), .b(FE_OFN577_n_9902), .o(g58087_db) );
na02f02 TIMEBOOST_cell_70647 ( .a(TIMEBOOST_net_22531), .b(g62723_sb), .o(n_5537) );
in01s01 g58088_u0 ( .a(FE_OFN576_n_9902), .o(g58088_sb) );
na02s01 g58088_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q), .b(FE_OFN576_n_9902), .o(g58088_db) );
na02m02 TIMEBOOST_cell_70936 ( .a(TIMEBOOST_net_20540), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_22676) );
in01s01 g58089_u0 ( .a(FE_OFN577_n_9902), .o(g58089_sb) );
na02s01 g58089_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q), .b(FE_OFN577_n_9902), .o(g58089_db) );
in01m01 g58090_u0 ( .a(FE_OFN574_n_9902), .o(g58090_sb) );
in01s01 TIMEBOOST_cell_73878 ( .a(n_8012), .o(TIMEBOOST_net_23443) );
na02m01 g58090_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q), .b(FE_OFN574_n_9902), .o(g58090_db) );
in01m01 g58091_u0 ( .a(FE_OFN577_n_9902), .o(g58091_sb) );
na04f02 TIMEBOOST_cell_73293 ( .a(n_1750), .b(g62716_sb), .c(g60682_da), .d(TIMEBOOST_net_22446), .o(n_5644) );
na02s01 TIMEBOOST_cell_38815 ( .a(TIMEBOOST_net_11019), .b(g65858_sb), .o(n_2581) );
in01s01 g58092_u0 ( .a(FE_OFN576_n_9902), .o(g58092_sb) );
na02s01 g58092_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q), .b(FE_OFN576_n_9902), .o(g58092_db) );
in01f02 g58093_u0 ( .a(FE_OFN575_n_9902), .o(g58093_sb) );
na03m02 TIMEBOOST_cell_73033 ( .a(TIMEBOOST_net_21741), .b(FE_OFN639_n_4669), .c(TIMEBOOST_net_23373), .o(TIMEBOOST_net_17029) );
na04f04 TIMEBOOST_cell_67686 ( .a(FE_OCPN1901_n_16810), .b(n_14911), .c(FE_OCPN1903_FE_OFN1061_n_16720), .d(TIMEBOOST_net_11894), .o(FE_RN_415_0) );
in01m02 g58094_u0 ( .a(FE_OFN577_n_9902), .o(g58094_sb) );
na02m02 g58094_u2 ( .a(FE_OFN577_n_9902), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q), .o(g58094_db) );
in01s01 g58095_u0 ( .a(FE_OFN576_n_9902), .o(g58095_sb) );
na03m06 TIMEBOOST_cell_73028 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(FE_OFN1031_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q), .o(TIMEBOOST_net_23311) );
na02s01 g58095_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q), .b(FE_OFN576_n_9902), .o(g58095_db) );
in01m01 g58096_u0 ( .a(FE_OFN574_n_9902), .o(g58096_sb) );
na03f06 TIMEBOOST_cell_73219 ( .a(TIMEBOOST_net_16956), .b(FE_OFN1148_n_13249), .c(g54137_sb), .o(n_13273) );
na03s01 TIMEBOOST_cell_72456 ( .a(pci_target_unit_del_sync_bc_in_202), .b(g66411_db), .c(g66399_sb), .o(n_2524) );
in01m02 g58097_u0 ( .a(FE_OFN574_n_9902), .o(g58097_sb) );
na02f01 TIMEBOOST_cell_54192 ( .a(TIMEBOOST_net_17313), .b(FE_OFN877_g64577_p), .o(TIMEBOOST_net_15152) );
na02s01 g58097_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q), .b(FE_OFN574_n_9902), .o(g58097_db) );
na03m02 TIMEBOOST_cell_65216 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q), .b(FE_OFN1676_n_4655), .c(n_4479), .o(TIMEBOOST_net_20366) );
na02s01 g58098_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q), .b(FE_OFN575_n_9902), .o(g58098_db) );
na02s01 TIMEBOOST_cell_48816 ( .a(TIMEBOOST_net_14625), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_11117) );
in01s01 g58099_u0 ( .a(FE_OFN534_n_9823), .o(g58099_sb) );
na02s01 g58099_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q), .b(FE_OFN534_n_9823), .o(g58099_db) );
na03f01 TIMEBOOST_cell_73294 ( .a(TIMEBOOST_net_328), .b(n_4098), .c(TIMEBOOST_net_17353), .o(n_6338) );
in01s01 g58100_u0 ( .a(FE_OFN535_n_9823), .o(g58100_sb) );
na02m02 TIMEBOOST_cell_50675 ( .a(g58306_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q), .o(TIMEBOOST_net_15555) );
na02m02 TIMEBOOST_cell_68965 ( .a(TIMEBOOST_net_21690), .b(TIMEBOOST_net_10576), .o(TIMEBOOST_net_17382) );
in01s01 g58101_u0 ( .a(FE_OFN519_n_9697), .o(g58101_sb) );
in01s02 g58102_u0 ( .a(FE_OFN595_n_9694), .o(g58102_sb) );
na02s01 g58102_u2 ( .a(FE_OFN595_n_9694), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q), .o(g58102_db) );
na02s01 TIMEBOOST_cell_43345 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_12567) );
in01s01 g58103_u0 ( .a(FE_OFN588_n_9692), .o(g58103_sb) );
na02m01 TIMEBOOST_cell_71912 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q), .b(FE_OFN1624_n_4438), .o(TIMEBOOST_net_23164) );
in01s01 g58104_u0 ( .a(FE_OFN587_n_9692), .o(g58104_sb) );
na03m06 TIMEBOOST_cell_68372 ( .a(FE_OFN906_n_4736), .b(TIMEBOOST_net_12319), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q), .o(TIMEBOOST_net_21394) );
na03m02 TIMEBOOST_cell_72718 ( .a(g64996_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q), .c(TIMEBOOST_net_16213), .o(TIMEBOOST_net_17540) );
na03s01 TIMEBOOST_cell_68086 ( .a(n_16871), .b(n_16864), .c(wishbone_slave_unit_pci_initiator_sm_rdata_selector), .o(TIMEBOOST_net_21251) );
in01m06 g58105_u0 ( .a(FE_OFN1803_n_9690), .o(g58105_sb) );
na02m02 TIMEBOOST_cell_71916 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q), .b(FE_OFN1625_n_4438), .o(TIMEBOOST_net_23166) );
na02m10 g58105_u2 ( .a(FE_OFN1803_n_9690), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q), .o(g58105_db) );
na02s01 TIMEBOOST_cell_53235 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_788), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q), .o(TIMEBOOST_net_16835) );
in01s01 g58106_u0 ( .a(FE_OFN602_n_9687), .o(g58106_sb) );
na03f02 TIMEBOOST_cell_73694 ( .a(n_9976), .b(n_10560), .c(FE_RN_233_0), .o(n_12133) );
in01s01 g58107_u0 ( .a(FE_OFN601_n_9687), .o(g58107_sb) );
na02s01 g58107_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q), .b(FE_OFN601_n_9687), .o(g58107_db) );
in01s02 g58108_u0 ( .a(FE_OFN600_n_9687), .o(g58108_sb) );
na03f04 TIMEBOOST_cell_64580 ( .a(TIMEBOOST_net_553), .b(n_4086), .c(n_15762), .o(n_4792) );
na02m02 TIMEBOOST_cell_68475 ( .a(TIMEBOOST_net_21445), .b(TIMEBOOST_net_10335), .o(TIMEBOOST_net_17480) );
in01s02 g58110_u0 ( .a(FE_OFN601_n_9687), .o(g58110_sb) );
na02m01 TIMEBOOST_cell_42802 ( .a(TIMEBOOST_net_12295), .b(FE_OFN935_n_2292), .o(TIMEBOOST_net_10234) );
na03f08 TIMEBOOST_cell_72433 ( .a(n_1986), .b(n_2929), .c(n_2931), .o(n_2930) );
in01s01 g58111_u0 ( .a(FE_OFN602_n_9687), .o(g58111_sb) );
in01s01 TIMEBOOST_cell_73967 ( .a(TIMEBOOST_net_23531), .o(TIMEBOOST_net_23532) );
na02s01 g58111_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q), .b(FE_OFN602_n_9687), .o(g58111_db) );
na02s02 TIMEBOOST_cell_38813 ( .a(TIMEBOOST_net_11018), .b(g65892_sb), .o(n_2572) );
in01s01 g58112_u0 ( .a(FE_OFN602_n_9687), .o(g58112_sb) );
na02m02 TIMEBOOST_cell_49351 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(FE_OFN1059_n_4727), .o(TIMEBOOST_net_14893) );
na02s01 g58112_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q), .b(FE_OFN602_n_9687), .o(g58112_db) );
na02f08 TIMEBOOST_cell_47530 ( .a(TIMEBOOST_net_13982), .b(n_279), .o(n_15370) );
in01s01 g58113_u0 ( .a(FE_OFN601_n_9687), .o(g58113_sb) );
na02m02 TIMEBOOST_cell_69572 ( .a(n_4442), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q), .o(TIMEBOOST_net_21994) );
na02s01 g58113_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q), .b(FE_OFN601_n_9687), .o(g58113_db) );
na02m02 TIMEBOOST_cell_49180 ( .a(TIMEBOOST_net_14807), .b(g61861_sb), .o(n_8116) );
in01s02 g58114_u0 ( .a(FE_OFN600_n_9687), .o(g58114_sb) );
na02f02 TIMEBOOST_cell_71038 ( .a(TIMEBOOST_net_20531), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_22727) );
na02m02 TIMEBOOST_cell_69003 ( .a(TIMEBOOST_net_21709), .b(TIMEBOOST_net_17221), .o(TIMEBOOST_net_13229) );
in01s02 g58115_u0 ( .a(FE_OFN600_n_9687), .o(g58115_sb) );
na02m02 TIMEBOOST_cell_48380 ( .a(TIMEBOOST_net_14407), .b(TIMEBOOST_net_10773), .o(TIMEBOOST_net_9458) );
in01s01 g58116_u0 ( .a(FE_OFN601_n_9687), .o(g58116_sb) );
na03s02 TIMEBOOST_cell_41726 ( .a(g58314_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q), .c(g58314_db), .o(n_9498) );
na02s01 g58116_u2 ( .a(FE_OFN601_n_9687), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q), .o(g58116_db) );
in01s01 g58117_u0 ( .a(FE_OFN602_n_9687), .o(g58117_sb) );
na03m02 TIMEBOOST_cell_72886 ( .a(g61864_sb), .b(g61896_db), .c(n_1886), .o(n_8034) );
in01s01 g58118_u0 ( .a(FE_OFN601_n_9687), .o(g58118_sb) );
na03m02 TIMEBOOST_cell_65074 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q), .c(FE_OFN1625_n_4438), .o(TIMEBOOST_net_16261) );
na02m10 TIMEBOOST_cell_52975 ( .a(wishbone_slave_unit_pcim_sm_data_in_661), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q), .o(TIMEBOOST_net_16705) );
na03f02 TIMEBOOST_cell_73774 ( .a(TIMEBOOST_net_13729), .b(FE_OFN1586_n_13736), .c(FE_OCP_RBN1996_n_13971), .o(n_14254) );
in01s01 g58119_u0 ( .a(FE_OFN601_n_9687), .o(g58119_sb) );
na03f02 TIMEBOOST_cell_73813 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_13777), .c(FE_OFN1769_n_14054), .o(g53223_p) );
na04m20 TIMEBOOST_cell_72435 ( .a(n_4725), .b(TIMEBOOST_net_16563), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q), .d(g60689_sb), .o(TIMEBOOST_net_20929) );
na02s01 TIMEBOOST_cell_51645 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q), .o(TIMEBOOST_net_16040) );
in01s01 g58120_u0 ( .a(FE_OFN2254_n_9687), .o(g58120_sb) );
na03m02 TIMEBOOST_cell_72792 ( .a(TIMEBOOST_net_23164), .b(g64982_sb), .c(TIMEBOOST_net_21850), .o(TIMEBOOST_net_17112) );
na04s02 TIMEBOOST_cell_67439 ( .a(wbs_dat_i_21_), .b(TIMEBOOST_net_577), .c(g63602_sb), .d(g63602_db), .o(n_7185) );
na03s02 TIMEBOOST_cell_72447 ( .a(pciu_pciif_idsel_reg_in), .b(g67051_sb), .c(TIMEBOOST_net_14099), .o(n_1452) );
no03s02 TIMEBOOST_cell_68088 ( .a(TIMEBOOST_net_9), .b(n_748), .c(TIMEBOOST_net_47), .o(TIMEBOOST_net_21252) );
na02s01 g58121_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q), .b(FE_OFN600_n_9687), .o(g58121_db) );
na02m10 TIMEBOOST_cell_45303 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q), .o(TIMEBOOST_net_13546) );
na03f02 TIMEBOOST_cell_34809 ( .a(TIMEBOOST_net_9481), .b(FE_OFN1392_n_8567), .c(g57118_sb), .o(n_11628) );
na02s01 g58122_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q), .b(FE_OFN600_n_9687), .o(g58122_db) );
na02m01 TIMEBOOST_cell_72022 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q), .b(FE_OFN648_n_4497), .o(TIMEBOOST_net_23219) );
in01s04 g58123_u0 ( .a(FE_OFN603_n_9687), .o(g58123_sb) );
na02m01 TIMEBOOST_cell_48669 ( .a(pci_target_unit_fifos_pciw_addr_data_in_145), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q), .o(TIMEBOOST_net_14552) );
na02f02 TIMEBOOST_cell_54356 ( .a(TIMEBOOST_net_17395), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_15520) );
na02m01 TIMEBOOST_cell_48671 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q), .o(TIMEBOOST_net_14553) );
in01s01 g58124_u0 ( .a(FE_OFN601_n_9687), .o(g58124_sb) );
na02s01 TIMEBOOST_cell_38558 ( .a(g57948_sb), .b(FE_OFN254_n_9825), .o(TIMEBOOST_net_10891) );
na02s01 TIMEBOOST_cell_45387 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q), .o(TIMEBOOST_net_13588) );
na02s01 TIMEBOOST_cell_38559 ( .a(TIMEBOOST_net_10891), .b(g57976_db), .o(n_9826) );
in01s01 g58125_u0 ( .a(FE_OFN601_n_9687), .o(g58125_sb) );
na02s02 TIMEBOOST_cell_38560 ( .a(g57938_sb), .b(FE_OFN241_n_9830), .o(TIMEBOOST_net_10892) );
na02m10 TIMEBOOST_cell_52977 ( .a(wishbone_slave_unit_pcim_sm_data_in_652), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q), .o(TIMEBOOST_net_16706) );
na02s02 TIMEBOOST_cell_38561 ( .a(TIMEBOOST_net_10892), .b(g57938_db), .o(n_9872) );
in01s01 g58126_u0 ( .a(FE_OFN602_n_9687), .o(g58126_sb) );
na02s02 TIMEBOOST_cell_52366 ( .a(TIMEBOOST_net_16400), .b(g58170_db), .o(TIMEBOOST_net_9378) );
na02s01 g58126_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q), .b(FE_OFN602_n_9687), .o(g58126_db) );
na02s01 TIMEBOOST_cell_47614 ( .a(TIMEBOOST_net_14024), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_401), .o(n_13228) );
in01m02 g58127_u0 ( .a(FE_OFN2253_n_9687), .o(g58127_sb) );
na02m02 TIMEBOOST_cell_68528 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q), .b(n_3741), .o(TIMEBOOST_net_21472) );
na02s01 TIMEBOOST_cell_38677 ( .a(TIMEBOOST_net_10950), .b(g63564_sb), .o(n_4598) );
in01s02 g58128_u0 ( .a(FE_OFN601_n_9687), .o(g58128_sb) );
na02s01 g58128_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q), .b(FE_OFN601_n_9687), .o(g58128_db) );
na02s01 TIMEBOOST_cell_49482 ( .a(TIMEBOOST_net_14958), .b(TIMEBOOST_net_12449), .o(TIMEBOOST_net_9420) );
in01s01 g58129_u0 ( .a(FE_OFN601_n_9687), .o(g58129_sb) );
na02f02 TIMEBOOST_cell_69955 ( .a(TIMEBOOST_net_22185), .b(g52638_db), .o(n_14753) );
na02f02 TIMEBOOST_cell_70133 ( .a(TIMEBOOST_net_22274), .b(g62010_sb), .o(n_7875) );
na02m02 g64783_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q), .b(FE_OFN669_n_4505), .o(g64783_db) );
in01s01 g58130_u0 ( .a(FE_OFN602_n_9687), .o(g58130_sb) );
na02s01 g58130_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q), .b(FE_OFN602_n_9687), .o(g58130_db) );
na02f02 TIMEBOOST_cell_70323 ( .a(TIMEBOOST_net_22369), .b(g62859_sb), .o(n_5248) );
na02f02 TIMEBOOST_cell_48626 ( .a(TIMEBOOST_net_14530), .b(g65229_sb), .o(n_2658) );
in01s02 g58132_u0 ( .a(FE_OFN601_n_9687), .o(g58132_sb) );
na02f10 TIMEBOOST_cell_52839 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_778), .o(TIMEBOOST_net_16637) );
na02s01 g58132_u2 ( .a(FE_OFN601_n_9687), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q), .o(g58132_db) );
na02f02 TIMEBOOST_cell_70927 ( .a(TIMEBOOST_net_22671), .b(g62454_sb), .o(n_6689) );
in01s01 g58133_u0 ( .a(FE_OFN602_n_9687), .o(g58133_sb) );
na03f02 TIMEBOOST_cell_35051 ( .a(TIMEBOOST_net_9603), .b(FE_OFN1436_n_9372), .c(g58456_sb), .o(n_9400) );
na02s01 g58133_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q), .b(FE_OFN602_n_9687), .o(g58133_db) );
na02m02 TIMEBOOST_cell_69421 ( .a(TIMEBOOST_net_21918), .b(g65002_sb), .o(TIMEBOOST_net_17577) );
na03f02 TIMEBOOST_cell_67875 ( .a(n_4672), .b(g64912_sb), .c(g64912_db), .o(TIMEBOOST_net_328) );
na02s02 TIMEBOOST_cell_43660 ( .a(TIMEBOOST_net_12724), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_11009) );
na03s02 TIMEBOOST_cell_73029 ( .a(TIMEBOOST_net_12720), .b(FE_OFN775_n_15366), .c(g65893_sb), .o(n_2583) );
na03f02 TIMEBOOST_cell_34755 ( .a(TIMEBOOST_net_9407), .b(FE_OFN1421_n_8567), .c(g57255_sb), .o(n_11499) );
in01s02 TIMEBOOST_cell_67102 ( .a(TIMEBOOST_net_21136), .o(n_2079) );
in01s01 g58136_u0 ( .a(FE_OFN602_n_9687), .o(g58136_sb) );
na02s01 TIMEBOOST_cell_38916 ( .a(FE_OFN1021_n_11877), .b(wbu_addr_in_279), .o(TIMEBOOST_net_11070) );
na02s01 g58137_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q), .b(FE_OFN600_n_9687), .o(g58137_db) );
in01s01 g58138_u0 ( .a(FE_OFN519_n_9697), .o(g58138_sb) );
na03f03 TIMEBOOST_cell_73711 ( .a(TIMEBOOST_net_13547), .b(n_12010), .c(FE_OFN1746_n_12004), .o(n_12649) );
na02s01 g58138_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q), .b(FE_OFN519_n_9697), .o(g58138_db) );
in01s01 TIMEBOOST_cell_63538 ( .a(TIMEBOOST_net_20718), .o(wbs_adr_i_10_) );
in01s02 g58139_u0 ( .a(FE_OFN517_n_9697), .o(g58139_sb) );
na03f10 TIMEBOOST_cell_64276 ( .a(conf_wb_err_addr_in_970), .b(conf_wb_err_addr_in_969), .c(n_531), .o(TIMEBOOST_net_12257) );
na02s02 g58139_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q), .b(FE_OFN517_n_9697), .o(g58139_db) );
na04f02 TIMEBOOST_cell_73220 ( .a(FE_OFN2022_n_4778), .b(TIMEBOOST_net_16658), .c(TIMEBOOST_net_629), .d(g63615_sb), .o(n_7145) );
in01s01 g58140_u0 ( .a(FE_OFN516_n_9697), .o(g58140_sb) );
na03s02 TIMEBOOST_cell_41734 ( .a(g58408_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q), .c(g58408_db), .o(n_9432) );
na02s01 g58140_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q), .b(FE_OFN516_n_9697), .o(g58140_db) );
in01s01 g58141_u0 ( .a(FE_OFN515_n_9697), .o(g58141_sb) );
na03f02 TIMEBOOST_cell_73568 ( .a(TIMEBOOST_net_17076), .b(FE_OFN1231_n_6391), .c(g62980_sb), .o(n_5922) );
na02s01 g58141_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q), .b(FE_OFN515_n_9697), .o(g58141_db) );
na02f02 TIMEBOOST_cell_54308 ( .a(TIMEBOOST_net_17371), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_15435) );
in01s01 g58142_u0 ( .a(FE_OFN517_n_9697), .o(g58142_sb) );
na02s01 g58142_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q), .b(FE_OFN517_n_9697), .o(g58142_db) );
na02f02 TIMEBOOST_cell_38971 ( .a(TIMEBOOST_net_11097), .b(g58311_db), .o(n_9500) );
in01s01 g58143_u0 ( .a(FE_OFN518_n_9697), .o(g58143_sb) );
na02s01 g58143_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q), .b(FE_OFN518_n_9697), .o(g58143_db) );
in01s01 g58144_u0 ( .a(FE_OFN518_n_9697), .o(g58144_sb) );
na02s01 g58144_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q), .b(FE_OFN518_n_9697), .o(g58144_db) );
in01s01 g58145_u0 ( .a(FE_OFN517_n_9697), .o(g58145_sb) );
na02s01 g58145_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q), .b(FE_OFN517_n_9697), .o(g58145_db) );
in01s01 g58146_u0 ( .a(FE_OFN517_n_9697), .o(g58146_sb) );
na03f02 TIMEBOOST_cell_34863 ( .a(TIMEBOOST_net_9414), .b(FE_OFN1397_n_8567), .c(g57261_sb), .o(n_10419) );
na02s01 g58146_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q), .b(FE_OFN517_n_9697), .o(g58146_db) );
na02s01 TIMEBOOST_cell_53961 ( .a(pci_target_unit_fifos_pcir_data_in), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q), .o(TIMEBOOST_net_17198) );
in01s01 g58147_u0 ( .a(FE_OFN517_n_9697), .o(g58147_sb) );
na02s01 g58147_u2 ( .a(FE_OFN517_n_9697), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q), .o(g58147_db) );
in01s01 g58148_u0 ( .a(FE_OFN517_n_9697), .o(g58148_sb) );
na02s01 g58148_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q), .b(FE_OFN517_n_9697), .o(g58148_db) );
in01s01 g58149_u0 ( .a(FE_OFN519_n_9697), .o(g58149_sb) );
na03s02 TIMEBOOST_cell_64411 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q), .b(FE_OFN603_n_9687), .c(g58123_sb), .o(TIMEBOOST_net_14651) );
na02s01 g58149_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q), .b(FE_OFN519_n_9697), .o(g58149_db) );
na02s01 TIMEBOOST_cell_53039 ( .a(configuration_pci_err_data_505), .b(wbm_dat_o_4_), .o(TIMEBOOST_net_16737) );
in01s01 g58150_u0 ( .a(FE_OFN518_n_9697), .o(g58150_sb) );
na03f02 TIMEBOOST_cell_65319 ( .a(TIMEBOOST_net_16309), .b(n_5633), .c(g62077_sb), .o(n_5634) );
na02s01 TIMEBOOST_cell_43021 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_140), .o(TIMEBOOST_net_12405) );
na03m02 TIMEBOOST_cell_72763 ( .a(TIMEBOOST_net_21542), .b(g64882_sb), .c(TIMEBOOST_net_21856), .o(TIMEBOOST_net_17368) );
na02s01 g58151_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q), .b(FE_OFN515_n_9697), .o(g58151_db) );
na02m06 TIMEBOOST_cell_71894 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q), .b(pci_target_unit_fifos_pciw_cbe_in), .o(TIMEBOOST_net_23155) );
in01s01 g58152_u0 ( .a(FE_OFN517_n_9697), .o(g58152_sb) );
no04f04 TIMEBOOST_cell_73801 ( .a(FE_RN_831_0), .b(FE_RN_832_0), .c(FE_RN_833_0), .d(n_16233), .o(n_16234) );
na02s02 TIMEBOOST_cell_48738 ( .a(TIMEBOOST_net_14586), .b(g57928_sb), .o(TIMEBOOST_net_9419) );
in01s01 g58153_u0 ( .a(FE_OFN516_n_9697), .o(g58153_sb) );
na02s01 g58153_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q), .b(FE_OFN516_n_9697), .o(g58153_db) );
na03s02 TIMEBOOST_cell_73092 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(FE_OFN2113_n_2053), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q), .o(TIMEBOOST_net_22250) );
in01s01 g58154_u0 ( .a(FE_OFN516_n_9697), .o(g58154_sb) );
na02s01 g58154_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q), .b(FE_OFN516_n_9697), .o(g58154_db) );
na02m02 TIMEBOOST_cell_63131 ( .a(TIMEBOOST_net_20512), .b(FE_OFN568_n_9528), .o(TIMEBOOST_net_16430) );
na02m02 TIMEBOOST_cell_53401 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(g65728_sb), .o(TIMEBOOST_net_16918) );
na02s01 g58155_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q), .b(FE_OFN517_n_9697), .o(g58155_db) );
na02m01 TIMEBOOST_cell_71868 ( .a(TIMEBOOST_net_17205), .b(FE_OFN1784_n_1699), .o(TIMEBOOST_net_23142) );
in01s01 g58156_u0 ( .a(FE_OFN516_n_9697), .o(g58156_sb) );
na03s01 TIMEBOOST_cell_72444 ( .a(g58054_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q), .c(g58042_sb), .o(TIMEBOOST_net_12402) );
na02m02 TIMEBOOST_cell_69579 ( .a(TIMEBOOST_net_21997), .b(TIMEBOOST_net_20286), .o(TIMEBOOST_net_14594) );
in01s01 TIMEBOOST_cell_35514 ( .a(TIMEBOOST_net_10105), .o(TIMEBOOST_net_10090) );
na02m02 TIMEBOOST_cell_48608 ( .a(TIMEBOOST_net_14521), .b(g65232_sb), .o(n_2655) );
na04f04 TIMEBOOST_cell_24555 ( .a(n_9227), .b(g57129_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q), .d(FE_OFN1402_n_8567), .o(n_10841) );
in01s01 g58158_u0 ( .a(FE_OFN518_n_9697), .o(g58158_sb) );
na02m10 TIMEBOOST_cell_45305 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q), .o(TIMEBOOST_net_13547) );
na02s01 g58158_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q), .b(FE_OFN518_n_9697), .o(g58158_db) );
na02m01 TIMEBOOST_cell_47577 ( .a(g58770_sb), .b(n_8831), .o(TIMEBOOST_net_14006) );
in01s01 g58159_u0 ( .a(FE_OFN517_n_9697), .o(g58159_sb) );
na02s01 g58159_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q), .b(FE_OFN517_n_9697), .o(g58159_db) );
na03f02 TIMEBOOST_cell_71160 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_385), .b(FE_OFN1001_n_15978), .c(g53940_sb), .o(TIMEBOOST_net_22788) );
in01m01 g58160_u0 ( .a(FE_OFN515_n_9697), .o(g58160_sb) );
na02s01 g58160_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q), .b(FE_OFN515_n_9697), .o(g58160_db) );
in01f10 g58161_u0 ( .a(FE_OFN515_n_9697), .o(g58161_sb) );
na02m06 TIMEBOOST_cell_38678 ( .a(g64242_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q), .o(TIMEBOOST_net_10951) );
na02m04 TIMEBOOST_cell_38679 ( .a(TIMEBOOST_net_10951), .b(g64242_db), .o(n_3930) );
in01s01 g58162_u0 ( .a(FE_OFN518_n_9697), .o(g58162_sb) );
na02f01 TIMEBOOST_cell_43412 ( .a(TIMEBOOST_net_12600), .b(g64786_db), .o(n_3765) );
na02s01 g58162_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q), .b(FE_OFN518_n_9697), .o(g58162_db) );
in01s01 g58163_u0 ( .a(FE_OFN517_n_9697), .o(g58163_sb) );
na02s02 TIMEBOOST_cell_47671 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q), .b(g65957_sb), .o(TIMEBOOST_net_14053) );
in01s01 g58164_u0 ( .a(FE_OFN515_n_9697), .o(g58164_sb) );
na03f02 TIMEBOOST_cell_73369 ( .a(TIMEBOOST_net_16717), .b(FE_OFN1301_n_5763), .c(g62035_sb), .o(n_7781) );
na02m01 TIMEBOOST_cell_63654 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q), .o(TIMEBOOST_net_20813) );
in01s01 g58165_u0 ( .a(FE_OFN518_n_9697), .o(g58165_sb) );
na02f01 TIMEBOOST_cell_72101 ( .a(TIMEBOOST_net_23258), .b(g64090_db), .o(n_4065) );
na02s01 g58165_u2 ( .a(FE_OFN518_n_9697), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q), .o(g58165_db) );
na02s02 TIMEBOOST_cell_63130 ( .a(FE_OFN245_n_9114), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q), .o(TIMEBOOST_net_20512) );
na02s01 g58166_u2 ( .a(FE_OFN517_n_9697), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q), .o(g58166_db) );
na03f02 TIMEBOOST_cell_67030 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_16531), .c(FE_OFN1600_n_13995), .o(n_14472) );
in01s01 g58167_u0 ( .a(FE_OFN517_n_9697), .o(g58167_sb) );
na02s01 TIMEBOOST_cell_69606 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_22011) );
na04m08 TIMEBOOST_cell_64827 ( .a(n_4465), .b(FE_OFN622_n_4409), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q), .d(g65013_sb), .o(n_4345) );
na02s01 g58168_u2 ( .a(FE_OFN516_n_9697), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q), .o(g58168_db) );
no02f02 TIMEBOOST_cell_51374 ( .a(TIMEBOOST_net_15904), .b(FE_RN_703_0), .o(FE_RN_704_0) );
in01s02 g58169_u0 ( .a(FE_OFN587_n_9692), .o(g58169_sb) );
na02m01 TIMEBOOST_cell_49261 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q), .b(FE_OFN574_n_9902), .o(TIMEBOOST_net_14848) );
na02f04 TIMEBOOST_cell_62905 ( .a(TIMEBOOST_net_20399), .b(FE_OFN1147_n_13249), .o(TIMEBOOST_net_15215) );
no02f02 TIMEBOOST_cell_71815 ( .a(TIMEBOOST_net_23115), .b(n_14434), .o(FE_RN_847_0) );
in01s01 g58170_u0 ( .a(FE_OFN588_n_9692), .o(g58170_sb) );
na02s02 TIMEBOOST_cell_49468 ( .a(TIMEBOOST_net_14951), .b(TIMEBOOST_net_13122), .o(TIMEBOOST_net_9356) );
na02s01 g58170_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q), .b(FE_OFN588_n_9692), .o(g58170_db) );
na02s02 TIMEBOOST_cell_71914 ( .a(g58192_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q), .o(TIMEBOOST_net_23165) );
in01s01 g58171_u0 ( .a(FE_OFN584_n_9692), .o(g58171_sb) );
na02m02 TIMEBOOST_cell_28409 ( .a(FE_OFN223_n_9844), .b(FE_OFN1692_n_9528), .o(TIMEBOOST_net_8309) );
na02s02 g58171_u2 ( .a(FE_OFN584_n_9692), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q), .o(g58171_db) );
na02f02 TIMEBOOST_cell_28410 ( .a(TIMEBOOST_net_8309), .b(g58284_da), .o(n_9518) );
in01s01 g58172_u0 ( .a(FE_OFN585_n_9692), .o(g58172_sb) );
na03s01 TIMEBOOST_cell_72457 ( .a(pci_target_unit_del_sync_bc_in_201), .b(FE_OFN2094_n_2520), .c(g66425_db), .o(n_2501) );
na02s02 TIMEBOOST_cell_49296 ( .a(TIMEBOOST_net_14865), .b(TIMEBOOST_net_10843), .o(TIMEBOOST_net_9479) );
in01s01 g58173_u0 ( .a(FE_OFN588_n_9692), .o(g58173_sb) );
na02f02 TIMEBOOST_cell_70654 ( .a(TIMEBOOST_net_20468), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_22535) );
na02s02 g58173_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q), .b(FE_OFN588_n_9692), .o(g58173_db) );
in01s01 g58174_u0 ( .a(FE_OFN589_n_9692), .o(g58174_sb) );
na02f02 TIMEBOOST_cell_70475 ( .a(TIMEBOOST_net_22445), .b(n_3373), .o(TIMEBOOST_net_415) );
na02s01 g58174_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q), .b(FE_OFN589_n_9692), .o(g58174_db) );
na02s01 TIMEBOOST_cell_38801 ( .a(TIMEBOOST_net_11012), .b(g65813_sb), .o(n_2574) );
in01s01 g58175_u0 ( .a(FE_OFN589_n_9692), .o(g58175_sb) );
na03f06 TIMEBOOST_cell_73174 ( .a(TIMEBOOST_net_16636), .b(g52634_sb), .c(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_5668) );
na02s01 g58175_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q), .b(FE_OFN589_n_9692), .o(g58175_db) );
na03f02 TIMEBOOST_cell_73453 ( .a(TIMEBOOST_net_17004), .b(FE_OFN1257_n_4143), .c(g62970_sb), .o(n_5942) );
in01s01 g58176_u0 ( .a(FE_OFN587_n_9692), .o(g58176_sb) );
na04f04 TIMEBOOST_cell_35023 ( .a(n_9053), .b(g57354_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q), .d(FE_OFN1407_n_8567), .o(n_10388) );
na02s01 g58176_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q), .b(FE_OFN587_n_9692), .o(g58176_db) );
na02m10 TIMEBOOST_cell_45623 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q), .o(TIMEBOOST_net_13706) );
in01s01 g58177_u0 ( .a(FE_OFN588_n_9692), .o(g58177_sb) );
na02m02 TIMEBOOST_cell_70223 ( .a(TIMEBOOST_net_22319), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_16413) );
na02s01 g58177_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q), .b(FE_OFN584_n_9692), .o(g58177_db) );
na04f04 TIMEBOOST_cell_73295 ( .a(TIMEBOOST_net_20415), .b(TIMEBOOST_net_7214), .c(FE_OFN877_g64577_p), .d(g63106_sb), .o(n_5042) );
in01s01 g58178_u0 ( .a(FE_OFN587_n_9692), .o(g58178_sb) );
na02s02 TIMEBOOST_cell_28413 ( .a(FE_OFN569_n_9528), .b(n_8892), .o(TIMEBOOST_net_8311) );
na04m04 TIMEBOOST_cell_36023 ( .a(g62005_sb), .b(n_2158), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q), .d(FE_OFN712_n_8140), .o(n_7885) );
in01s02 g58179_u0 ( .a(FE_OFN587_n_9692), .o(g58179_sb) );
no04f06 TIMEBOOST_cell_64368 ( .a(n_2869), .b(n_287), .c(FE_RN_627_0), .d(FE_RN_628_0), .o(TIMEBOOST_net_155) );
na02s01 g58179_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q), .b(FE_OFN587_n_9692), .o(g58179_db) );
na03f02 TIMEBOOST_cell_72981 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(FE_OFN1055_n_4727), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q), .o(TIMEBOOST_net_22144) );
in01s01 g58180_u0 ( .a(FE_OFN588_n_9692), .o(g58180_sb) );
na02f02 TIMEBOOST_cell_71163 ( .a(TIMEBOOST_net_22789), .b(g54199_sb), .o(n_13419) );
na03f02 TIMEBOOST_cell_66879 ( .a(FE_OFN1562_n_12502), .b(FE_OCPN1825_n_12030), .c(TIMEBOOST_net_13537), .o(n_12510) );
na02m02 TIMEBOOST_cell_68869 ( .a(TIMEBOOST_net_21642), .b(TIMEBOOST_net_10431), .o(TIMEBOOST_net_21034) );
in01s01 g58181_u0 ( .a(FE_OFN585_n_9692), .o(g58181_sb) );
na04f04 TIMEBOOST_cell_35024 ( .a(n_8993), .b(g57591_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q), .d(FE_OFN1384_n_8567), .o(n_10288) );
in01s01 TIMEBOOST_cell_63547 ( .a(TIMEBOOST_net_20726), .o(TIMEBOOST_net_20727) );
na04f04 TIMEBOOST_cell_35025 ( .a(n_9413), .b(g57582_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q), .d(FE_OFN1385_n_8567), .o(n_11167) );
in01s01 g58182_u0 ( .a(FE_OFN588_n_9692), .o(g58182_sb) );
na03m06 TIMEBOOST_cell_69914 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q), .b(FE_OFN1051_n_16657), .c(pci_target_unit_fifos_pciw_addr_data_in_137), .o(TIMEBOOST_net_22165) );
na02f02 TIMEBOOST_cell_70071 ( .a(TIMEBOOST_net_22243), .b(g61704_sb), .o(n_8419) );
na02f02 TIMEBOOST_cell_71491 ( .a(TIMEBOOST_net_22953), .b(TIMEBOOST_net_8849), .o(n_14821) );
in01s01 g58183_u0 ( .a(FE_OFN584_n_9692), .o(g58183_sb) );
in01s01 TIMEBOOST_cell_73839 ( .a(TIMEBOOST_net_23403), .o(TIMEBOOST_net_23404) );
na02s02 g58183_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q), .b(FE_OFN584_n_9692), .o(g58183_db) );
in01s01 g58184_u0 ( .a(FE_OFN585_n_9692), .o(g58184_sb) );
na02s01 TIMEBOOST_cell_50035 ( .a(configuration_pci_err_data_532), .b(wbm_dat_o_31_), .o(TIMEBOOST_net_15235) );
na02s01 TIMEBOOST_cell_52397 ( .a(g58488_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q), .o(TIMEBOOST_net_16416) );
in01s02 g58185_u0 ( .a(FE_OFN584_n_9692), .o(g58185_sb) );
na03f02 TIMEBOOST_cell_73606 ( .a(TIMEBOOST_net_17551), .b(FE_OFN1213_n_4151), .c(g62388_sb), .o(n_6824) );
na02s02 TIMEBOOST_cell_70868 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q), .o(TIMEBOOST_net_22642) );
na02m02 TIMEBOOST_cell_69560 ( .a(g64851_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q), .o(TIMEBOOST_net_21988) );
in01s01 g58186_u0 ( .a(FE_OFN584_n_9692), .o(g58186_sb) );
na02m02 TIMEBOOST_cell_53014 ( .a(TIMEBOOST_net_16724), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_15312) );
na02m06 TIMEBOOST_cell_45475 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q), .o(TIMEBOOST_net_13632) );
na04m08 TIMEBOOST_cell_72950 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q), .b(FE_OFN1810_n_4454), .c(n_3747), .d(g64919_sb), .o(n_3684) );
in01s01 g58187_u0 ( .a(FE_OFN589_n_9692), .o(g58187_sb) );
na03f02 TIMEBOOST_cell_72951 ( .a(pci_target_unit_del_sync_addr_in_214), .b(g65247_sb), .c(TIMEBOOST_net_7157), .o(n_2635) );
na02s01 g58187_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q), .b(FE_OFN589_n_9692), .o(g58187_db) );
in01s01 g58188_u0 ( .a(FE_OFN588_n_9692), .o(g58188_sb) );
na03m02 TIMEBOOST_cell_72822 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q), .b(g65332_sb), .c(TIMEBOOST_net_22261), .o(TIMEBOOST_net_17432) );
in01s02 g58189_u0 ( .a(FE_OFN587_n_9692), .o(g58189_sb) );
na02s01 TIMEBOOST_cell_53963 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q), .o(TIMEBOOST_net_17199) );
na02s02 TIMEBOOST_cell_52398 ( .a(TIMEBOOST_net_16416), .b(TIMEBOOST_net_11195), .o(TIMEBOOST_net_9449) );
in01m06 g58190_u0 ( .a(FE_OFN585_n_9692), .o(g58190_sb) );
na02m02 TIMEBOOST_cell_69561 ( .a(TIMEBOOST_net_21988), .b(TIMEBOOST_net_14398), .o(TIMEBOOST_net_17124) );
na02m08 g58190_u2 ( .a(FE_OFN585_n_9692), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q), .o(g58190_db) );
na02f04 TIMEBOOST_cell_69852 ( .a(pciu_am1_in_534), .b(n_4806), .o(TIMEBOOST_net_22134) );
in01s01 g58191_u0 ( .a(FE_OFN589_n_9692), .o(g58191_sb) );
na02m02 TIMEBOOST_cell_69072 ( .a(n_38), .b(FE_OFN619_n_4490), .o(TIMEBOOST_net_21744) );
na02s01 g58191_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q), .b(FE_OFN589_n_9692), .o(g58191_db) );
na02s02 TIMEBOOST_cell_63007 ( .a(TIMEBOOST_net_20450), .b(g57994_sb), .o(TIMEBOOST_net_14469) );
in01s02 g58192_u0 ( .a(FE_OFN587_n_9692), .o(g58192_sb) );
na02s01 TIMEBOOST_cell_45307 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q), .o(TIMEBOOST_net_13548) );
in01s01 g58193_u0 ( .a(FE_OFN589_n_9692), .o(g58193_sb) );
na02s02 g58193_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q), .b(FE_OFN589_n_9692), .o(g58193_db) );
na03s01 TIMEBOOST_cell_22706 ( .a(FE_OFN270_n_9836), .b(g58158_sb), .c(g58158_db), .o(n_9631) );
in01s01 g58194_u0 ( .a(FE_OFN585_n_9692), .o(g58194_sb) );
in01s01 TIMEBOOST_cell_63546 ( .a(pci_target_unit_fifos_pcir_data_in_187), .o(TIMEBOOST_net_20726) );
in01s01 TIMEBOOST_cell_73879 ( .a(TIMEBOOST_net_23443), .o(TIMEBOOST_net_23444) );
in01s01 g58195_u0 ( .a(FE_OFN585_n_9692), .o(g58195_sb) );
na02m01 TIMEBOOST_cell_4282 ( .a(g52485_da), .b(FE_OFN1025_n_11877), .o(TIMEBOOST_net_701) );
na02s01 TIMEBOOST_cell_62978 ( .a(configuration_wb_err_addr_557), .b(conf_wb_err_addr_in_966), .o(TIMEBOOST_net_20436) );
na02s02 TIMEBOOST_cell_63309 ( .a(TIMEBOOST_net_20601), .b(g58229_sb), .o(TIMEBOOST_net_9354) );
in01s02 g58196_u0 ( .a(FE_OFN587_n_9692), .o(g58196_sb) );
na03f02 TIMEBOOST_cell_73544 ( .a(TIMEBOOST_net_17079), .b(FE_OFN1230_n_6391), .c(g62987_sb), .o(n_5908) );
na03s01 TIMEBOOST_cell_68132 ( .a(g54216_sb), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_406), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q), .o(TIMEBOOST_net_21274) );
na03m02 TIMEBOOST_cell_73545 ( .a(TIMEBOOST_net_7598), .b(g54194_sb), .c(g54194_db), .o(n_13357) );
in01s01 g58197_u0 ( .a(FE_OFN584_n_9692), .o(g58197_sb) );
na02s03 TIMEBOOST_cell_4278 ( .a(g52483_da), .b(FE_OFN8_n_11877), .o(TIMEBOOST_net_699) );
na02s01 g58197_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q), .b(FE_OFN584_n_9692), .o(g58197_db) );
in01s01 g58198_u0 ( .a(FE_OFN595_n_9694), .o(g58198_sb) );
na02m10 TIMEBOOST_cell_69602 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q), .o(TIMEBOOST_net_22009) );
na02s01 g58198_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q), .b(FE_OFN595_n_9694), .o(g58198_db) );
na02m01 TIMEBOOST_cell_69152 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q), .o(TIMEBOOST_net_21784) );
in01s01 g58199_u0 ( .a(FE_OFN596_n_9694), .o(g58199_sb) );
na02s01 g58199_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q), .b(FE_OFN596_n_9694), .o(g58199_db) );
na03m02 TIMEBOOST_cell_73093 ( .a(g65324_da), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q), .c(TIMEBOOST_net_14662), .o(TIMEBOOST_net_17395) );
in01s01 g58200_u0 ( .a(FE_OFN592_n_9694), .o(g58200_sb) );
na03f02 TIMEBOOST_cell_67020 ( .a(FE_OFN1586_n_13736), .b(TIMEBOOST_net_16071), .c(FE_OCP_RBN1999_n_13971), .o(n_16207) );
na02s01 g58200_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q), .b(FE_OFN592_n_9694), .o(g58200_db) );
na03f06 TIMEBOOST_cell_64364 ( .a(n_1414), .b(n_1413), .c(n_2228), .o(TIMEBOOST_net_88) );
in01s01 g58201_u0 ( .a(FE_OFN593_n_9694), .o(g58201_sb) );
na02s01 g58201_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q), .b(FE_OFN593_n_9694), .o(g58201_db) );
na02m02 TIMEBOOST_cell_68568 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q), .b(FE_OFN630_n_4454), .o(TIMEBOOST_net_21492) );
in01s01 g58202_u0 ( .a(FE_OFN596_n_9694), .o(g58202_sb) );
na02s01 g58202_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q), .b(FE_OFN596_n_9694), .o(g58202_db) );
na02m02 TIMEBOOST_cell_4266 ( .a(g52475_da), .b(FE_OFN1023_n_11877), .o(TIMEBOOST_net_693) );
in01s01 g58203_u0 ( .a(FE_OFN597_n_9694), .o(g58203_sb) );
na02s01 g58203_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q), .b(FE_OFN597_n_9694), .o(g58203_db) );
na03f02 TIMEBOOST_cell_73546 ( .a(TIMEBOOST_net_17070), .b(FE_OFN1230_n_6391), .c(g62370_sb), .o(n_6863) );
in01s02 g58204_u0 ( .a(FE_OFN597_n_9694), .o(g58204_sb) );
na02s01 g58204_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN597_n_9694), .o(g58204_db) );
in01s02 g58205_u0 ( .a(FE_OFN592_n_9694), .o(g58205_sb) );
na03f10 TIMEBOOST_cell_70286 ( .a(TIMEBOOST_net_14988), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q), .c(FE_OFN1147_n_13249), .o(TIMEBOOST_net_22351) );
na02f02 TIMEBOOST_cell_30899 ( .a(n_9035), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q), .o(TIMEBOOST_net_9554) );
in01s02 g58206_u0 ( .a(FE_OFN596_n_9694), .o(g58206_sb) );
na02f01 TIMEBOOST_cell_28423 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(FE_OFN1031_n_4732), .o(TIMEBOOST_net_8316) );
na02f01 TIMEBOOST_cell_71774 ( .a(TIMEBOOST_net_13698), .b(FE_OFN1774_n_13800), .o(TIMEBOOST_net_23095) );
in01s01 g58207_u0 ( .a(FE_OFN595_n_9694), .o(g58207_sb) );
na03m06 TIMEBOOST_cell_67823 ( .a(n_3744), .b(n_83), .c(FE_OFN667_n_4495), .o(TIMEBOOST_net_10432) );
na02s01 g58207_u2 ( .a(FE_OFN595_n_9694), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q), .o(g58207_db) );
na02f02 TIMEBOOST_cell_70834 ( .a(TIMEBOOST_net_16694), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_22625) );
in01s01 g58208_u0 ( .a(FE_OFN595_n_9694), .o(g58208_sb) );
na03m02 TIMEBOOST_cell_72556 ( .a(g64770_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q), .c(TIMEBOOST_net_14464), .o(TIMEBOOST_net_13225) );
na02s01 g58208_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q), .b(FE_OFN595_n_9694), .o(g58208_db) );
na03f02 TIMEBOOST_cell_73607 ( .a(TIMEBOOST_net_17469), .b(FE_OFN1206_n_6356), .c(g63174_sb), .o(n_5796) );
in01s02 g58209_u0 ( .a(FE_OFN597_n_9694), .o(g58209_sb) );
na02s01 g58209_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q), .b(FE_OFN597_n_9694), .o(g58209_db) );
in01s02 g58210_u0 ( .a(FE_OFN595_n_9694), .o(g58210_sb) );
na03m02 TIMEBOOST_cell_72697 ( .a(TIMEBOOST_net_21566), .b(FE_OFN649_n_4497), .c(TIMEBOOST_net_21915), .o(TIMEBOOST_net_13247) );
na02s01 g58210_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN595_n_9694), .o(g58210_db) );
na03s01 TIMEBOOST_cell_64307 ( .a(TIMEBOOST_net_8632), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q), .o(TIMEBOOST_net_16811) );
in01s01 g58211_u0 ( .a(FE_OFN596_n_9694), .o(g58211_sb) );
na03s02 TIMEBOOST_cell_46695 ( .a(TIMEBOOST_net_12804), .b(g58325_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q), .o(TIMEBOOST_net_9446) );
in01s01 TIMEBOOST_cell_73880 ( .a(n_7957), .o(TIMEBOOST_net_23445) );
in01s02 g58212_u0 ( .a(FE_OFN592_n_9694), .o(g58212_sb) );
na04f04 TIMEBOOST_cell_67700 ( .a(TIMEBOOST_net_16859), .b(FE_OFN2198_n_10256), .c(g52608_sb), .d(TIMEBOOST_net_698), .o(n_11863) );
na02s01 TIMEBOOST_cell_42881 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q), .o(TIMEBOOST_net_12335) );
in01s01 g58213_u0 ( .a(FE_OFN592_n_9694), .o(g58213_sb) );
na02m04 TIMEBOOST_cell_69068 ( .a(g64863_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_21742) );
na02s01 g58213_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q), .b(FE_OFN592_n_9694), .o(g58213_db) );
na02f02 TIMEBOOST_cell_69753 ( .a(TIMEBOOST_net_22084), .b(g65940_db), .o(n_2579) );
in01s01 g58214_u0 ( .a(FE_OFN593_n_9694), .o(g58214_sb) );
no03f04 TIMEBOOST_cell_71814 ( .a(FE_RN_845_0), .b(FE_RN_844_0), .c(FE_RN_843_0), .o(TIMEBOOST_net_23115) );
na02s01 g58214_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q), .b(FE_OFN593_n_9694), .o(g58214_db) );
na02s02 TIMEBOOST_cell_52231 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q), .b(g65842_sb), .o(TIMEBOOST_net_16333) );
in01s01 g58215_u0 ( .a(FE_OFN596_n_9694), .o(g58215_sb) );
na04f04 TIMEBOOST_cell_67694 ( .a(TIMEBOOST_net_16854), .b(FE_OFN2198_n_10256), .c(g52622_sb), .d(TIMEBOOST_net_701), .o(n_11849) );
na03f02 TIMEBOOST_cell_66691 ( .a(TIMEBOOST_net_16787), .b(FE_OFN1315_n_6624), .c(g62622_sb), .o(n_6313) );
in01s01 g58216_u0 ( .a(FE_OFN596_n_9694), .o(g58216_sb) );
na02f01 TIMEBOOST_cell_54220 ( .a(TIMEBOOST_net_17327), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_15147) );
na02s01 TIMEBOOST_cell_42885 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q), .o(TIMEBOOST_net_12337) );
in01s02 g58217_u0 ( .a(FE_OFN597_n_9694), .o(g58217_sb) );
na02s01 g58217_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q), .b(FE_OFN597_n_9694), .o(g58217_db) );
in01s01 g58218_u0 ( .a(FE_OFN596_n_9694), .o(g58218_sb) );
na02m02 TIMEBOOST_cell_62826 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q), .b(pci_target_unit_fifos_pciw_control_in_156), .o(TIMEBOOST_net_20360) );
na02m01 TIMEBOOST_cell_68740 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q), .b(FE_OFN661_n_4392), .o(TIMEBOOST_net_21578) );
in01s01 g58219_u0 ( .a(FE_OFN595_n_9694), .o(g58219_sb) );
na02s01 TIMEBOOST_cell_51897 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q), .o(TIMEBOOST_net_16166) );
na02s01 g58219_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN595_n_9694), .o(g58219_db) );
in01s01 g58220_u0 ( .a(FE_OFN595_n_9694), .o(g58220_sb) );
na02s01 TIMEBOOST_cell_63006 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q), .o(TIMEBOOST_net_20450) );
na03f02 TIMEBOOST_cell_66661 ( .a(TIMEBOOST_net_13379), .b(n_6554), .c(g62677_sb), .o(n_6186) );
in01s01 g58221_u0 ( .a(FE_OFN597_n_9694), .o(g58221_sb) );
na04m04 TIMEBOOST_cell_46517 ( .a(n_2187), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q), .c(FE_OFN713_n_8140), .d(g61728_sb), .o(n_8364) );
na03f02 TIMEBOOST_cell_73547 ( .a(TIMEBOOST_net_20603), .b(FE_OFN1235_n_6391), .c(g62623_sb), .o(n_6311) );
in01s02 g58222_u0 ( .a(FE_OFN592_n_9694), .o(g58222_sb) );
na02s02 g58222_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q), .b(FE_OFN593_n_9694), .o(g58222_db) );
na03f02 TIMEBOOST_cell_66058 ( .a(TIMEBOOST_net_16760), .b(g62840_sb), .c(FE_OFN1139_g64577_p), .o(n_5293) );
in01s01 g58223_u0 ( .a(FE_OFN595_n_9694), .o(g58223_sb) );
na02s01 g58223_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q), .b(FE_OFN595_n_9694), .o(g58223_db) );
na04s03 TIMEBOOST_cell_72897 ( .a(TIMEBOOST_net_12626), .b(FE_OFN1044_n_2037), .c(g65901_sb), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q), .o(TIMEBOOST_net_22080) );
in01s01 g58224_u0 ( .a(FE_OFN597_n_9694), .o(g58224_sb) );
na02m02 TIMEBOOST_cell_69144 ( .a(n_4498), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q), .o(TIMEBOOST_net_21780) );
na02s01 g58224_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q), .b(FE_OFN597_n_9694), .o(g58224_db) );
na02s01 TIMEBOOST_cell_30991 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_29__Q), .b(n_9834), .o(TIMEBOOST_net_9600) );
in01s01 g58225_u0 ( .a(FE_OFN593_n_9694), .o(g58225_sb) );
na02s02 TIMEBOOST_cell_37884 ( .a(g58123_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q), .o(TIMEBOOST_net_10554) );
na02s02 g58225_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN593_n_9694), .o(g58225_db) );
na02m02 TIMEBOOST_cell_68091 ( .a(TIMEBOOST_net_21253), .b(g66433_db), .o(n_1533) );
na02s04 TIMEBOOST_cell_51979 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q), .b(TIMEBOOST_net_13875), .o(TIMEBOOST_net_16207) );
in01s01 g58227_u0 ( .a(FE_OFN595_n_9694), .o(g58227_sb) );
na03f06 TIMEBOOST_cell_73296 ( .a(TIMEBOOST_net_20929), .b(FE_OFN1126_g64577_p), .c(g59381_sb), .o(n_7677) );
na02s01 g58227_u2 ( .a(FE_OFN595_n_9694), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q), .o(g58227_db) );
na02m01 TIMEBOOST_cell_26431 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN1046_n_16657), .o(TIMEBOOST_net_7320) );
in01s01 g58228_u0 ( .a(FE_OFN592_n_9694), .o(g58228_sb) );
na02m02 TIMEBOOST_cell_51202 ( .a(TIMEBOOST_net_15818), .b(g63162_sb), .o(n_5812) );
na02s01 g58228_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q), .b(FE_OFN592_n_9694), .o(g58228_db) );
na02m02 TIMEBOOST_cell_54071 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_147), .o(TIMEBOOST_net_17253) );
in01s01 g58229_u0 ( .a(FE_OFN540_n_9690), .o(g58229_sb) );
na03f02 TIMEBOOST_cell_66729 ( .a(TIMEBOOST_net_16835), .b(FE_OFN1305_n_13124), .c(g54353_sb), .o(n_13088) );
na02s02 g58229_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q), .b(FE_OFN540_n_9690), .o(g58229_db) );
in01s02 TIMEBOOST_cell_45988 ( .a(TIMEBOOST_net_13948), .o(TIMEBOOST_net_13949) );
in01m01 g58230_u0 ( .a(FE_OFN539_n_9690), .o(g58230_sb) );
na03f02 TIMEBOOST_cell_73548 ( .a(TIMEBOOST_net_22788), .b(g54174_sb), .c(g54174_db), .o(TIMEBOOST_net_11792) );
na03f02 TIMEBOOST_cell_73549 ( .a(TIMEBOOST_net_17068), .b(FE_OFN1233_n_6391), .c(g63155_sb), .o(n_5830) );
na03s02 TIMEBOOST_cell_72891 ( .a(g61812_sb), .b(g61812_db), .c(n_1603), .o(n_8168) );
in01s02 g58231_u0 ( .a(FE_OFN1801_n_9690), .o(g58231_sb) );
na02s01 TIMEBOOST_cell_29373 ( .a(parchk_pci_ad_out_in_1196), .b(configuration_wb_err_data_599), .o(TIMEBOOST_net_8791) );
na02m02 TIMEBOOST_cell_53843 ( .a(n_4330), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_17139) );
in01s02 g58232_u0 ( .a(FE_OFN540_n_9690), .o(g58232_sb) );
na02f02 TIMEBOOST_cell_42830 ( .a(TIMEBOOST_net_12309), .b(g58795_sb), .o(n_9112) );
na03f02 TIMEBOOST_cell_73550 ( .a(TIMEBOOST_net_17067), .b(FE_OFN1233_n_6391), .c(g62941_sb), .o(n_5999) );
na02s01 TIMEBOOST_cell_38445 ( .a(TIMEBOOST_net_10834), .b(g57982_db), .o(n_9110) );
in01s01 g58233_u0 ( .a(FE_OFN543_n_9690), .o(g58233_sb) );
na02m02 TIMEBOOST_cell_48030 ( .a(TIMEBOOST_net_14232), .b(FE_OFN250_n_9789), .o(TIMEBOOST_net_10773) );
na02s01 g58233_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q), .b(FE_OFN543_n_9690), .o(g58233_db) );
in01s01 g58234_u0 ( .a(FE_OFN543_n_9690), .o(g58234_sb) );
na02s01 g58234_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q), .b(FE_OFN543_n_9690), .o(g58234_db) );
na02s02 TIMEBOOST_cell_38273 ( .a(TIMEBOOST_net_10748), .b(g58062_db), .o(n_9090) );
in01s01 g58235_u0 ( .a(FE_OFN1800_n_9690), .o(g58235_sb) );
na03f02 TIMEBOOST_cell_24140 ( .a(FE_OFN1398_n_8567), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .c(n_9341), .o(n_9343) );
na02f02 TIMEBOOST_cell_40084 ( .a(FE_OFN1186_n_3476), .b(configuration_pci_err_addr_476), .o(TIMEBOOST_net_11654) );
in01s01 g58236_u0 ( .a(FE_OFN540_n_9690), .o(g58236_sb) );
in01s01 TIMEBOOST_cell_63556 ( .a(TIMEBOOST_net_20736), .o(wbs_adr_i_24_) );
na03f02 TIMEBOOST_cell_73551 ( .a(TIMEBOOST_net_17556), .b(FE_OFN2063_n_6391), .c(g62339_sb), .o(n_6920) );
na03f02 TIMEBOOST_cell_73552 ( .a(TIMEBOOST_net_17073), .b(FE_OFN1235_n_6391), .c(g62465_sb), .o(n_6665) );
in01s01 g58237_u0 ( .a(FE_OFN542_n_9690), .o(g58237_sb) );
na03s02 TIMEBOOST_cell_48861 ( .a(g58225_sb), .b(g58225_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q), .o(TIMEBOOST_net_14648) );
in01s01 g58238_u0 ( .a(FE_OFN542_n_9690), .o(g58238_sb) );
na02f02 TIMEBOOST_cell_70655 ( .a(TIMEBOOST_net_22535), .b(g62853_sb), .o(n_5263) );
na02f02 TIMEBOOST_cell_70599 ( .a(TIMEBOOST_net_22507), .b(g62797_sb), .o(n_5391) );
in01m01 g58239_u0 ( .a(FE_OFN539_n_9690), .o(g58239_sb) );
na02m02 TIMEBOOST_cell_68934 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_21675) );
na02f02 TIMEBOOST_cell_49930 ( .a(TIMEBOOST_net_15182), .b(g63113_sb), .o(n_5029) );
in01s02 g58240_u0 ( .a(FE_OFN1801_n_9690), .o(g58240_sb) );
na02m02 TIMEBOOST_cell_4288 ( .a(g52473_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_704) );
na03f02 TIMEBOOST_cell_73221 ( .a(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .b(n_16452), .c(n_7725), .o(TIMEBOOST_net_376) );
na02m04 TIMEBOOST_cell_37122 ( .a(n_2305), .b(n_2756), .o(TIMEBOOST_net_10173) );
na02m02 TIMEBOOST_cell_69005 ( .a(TIMEBOOST_net_21710), .b(g64871_sb), .o(TIMEBOOST_net_12542) );
na02s01 g58241_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q), .b(FE_OFN542_n_9690), .o(g58241_db) );
na03m02 TIMEBOOST_cell_68692 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN684_n_4417), .c(g64898_sb), .o(TIMEBOOST_net_21554) );
in01s01 g58242_u0 ( .a(FE_OFN1802_n_9690), .o(g58242_sb) );
na02s01 TIMEBOOST_cell_47642 ( .a(TIMEBOOST_net_14038), .b(TIMEBOOST_net_9652), .o(TIMEBOOST_net_12829) );
in01s01 g58243_u0 ( .a(FE_OFN542_n_9690), .o(g58243_sb) );
na02s01 g58243_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q), .b(FE_OFN542_n_9690), .o(g58243_db) );
na02s01 TIMEBOOST_cell_44176 ( .a(TIMEBOOST_net_12982), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9529) );
in01s01 g58244_u0 ( .a(FE_OFN540_n_9690), .o(g58244_sb) );
na02m02 TIMEBOOST_cell_69423 ( .a(TIMEBOOST_net_21919), .b(g64951_sb), .o(TIMEBOOST_net_12687) );
na03f02 TIMEBOOST_cell_72879 ( .a(g64346_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q), .c(TIMEBOOST_net_14493), .o(TIMEBOOST_net_8343) );
na02s01 TIMEBOOST_cell_25309 ( .a(pci_ad_i_4_), .b(parchk_pci_ad_reg_in_1208), .o(TIMEBOOST_net_6759) );
na03m02 TIMEBOOST_cell_72764 ( .a(TIMEBOOST_net_21524), .b(g65095_sb), .c(TIMEBOOST_net_21780), .o(TIMEBOOST_net_21032) );
na02s01 g58245_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q), .b(FE_OFN540_n_9690), .o(g58245_db) );
na03m02 TIMEBOOST_cell_66057 ( .a(TIMEBOOST_net_16579), .b(FE_OFN1655_n_9502), .c(g58418_sb), .o(n_8998) );
na02m02 TIMEBOOST_cell_68477 ( .a(TIMEBOOST_net_21446), .b(FE_OFN951_n_2055), .o(TIMEBOOST_net_16200) );
na02m02 TIMEBOOST_cell_69063 ( .a(TIMEBOOST_net_21739), .b(g64129_sb), .o(n_4033) );
na02f02 TIMEBOOST_cell_50554 ( .a(TIMEBOOST_net_15494), .b(g62946_sb), .o(n_5989) );
na02m02 TIMEBOOST_cell_69963 ( .a(TIMEBOOST_net_22189), .b(g60686_sb), .o(TIMEBOOST_net_13086) );
na02s01 TIMEBOOST_cell_38407 ( .a(TIMEBOOST_net_10815), .b(g58080_db), .o(n_9714) );
na02s01 g58248_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q), .b(FE_OFN542_n_9690), .o(g58248_db) );
na02m02 TIMEBOOST_cell_69688 ( .a(FE_OFN1680_n_4655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q), .o(TIMEBOOST_net_22052) );
na03m02 TIMEBOOST_cell_71920 ( .a(n_3752), .b(g64849_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q), .o(TIMEBOOST_net_23168) );
na02s01 g58249_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q), .b(FE_OFN543_n_9690), .o(g58249_db) );
na02m08 TIMEBOOST_cell_63780 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(TIMEBOOST_net_20876) );
na03f02 TIMEBOOST_cell_72529 ( .a(TIMEBOOST_net_21398), .b(g64147_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q), .o(TIMEBOOST_net_20473) );
in01m02 g58251_u0 ( .a(FE_OFN541_n_9690), .o(g58251_sb) );
na03f04 TIMEBOOST_cell_70140 ( .a(FE_OFN923_n_4740), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q), .c(pci_target_unit_fifos_pciw_cbe_in_153), .o(TIMEBOOST_net_22278) );
na02m04 g58251_u2 ( .a(FE_OFN541_n_9690), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q), .o(g58251_db) );
na03f02 TIMEBOOST_cell_34900 ( .a(TIMEBOOST_net_9447), .b(FE_OFN1407_n_8567), .c(g57265_sb), .o(n_11487) );
in01s01 g58252_u0 ( .a(FE_OFN543_n_9690), .o(g58252_sb) );
na02m01 TIMEBOOST_cell_4280 ( .a(g52471_da), .b(FE_OFN1023_n_11877), .o(TIMEBOOST_net_700) );
na02m01 g52470_u1 ( .a(wbs_adr_i_24_), .b(g52470_sb), .o(g52470_da) );
na02s01 TIMEBOOST_cell_62475 ( .a(TIMEBOOST_net_20184), .b(g54205_sb), .o(TIMEBOOST_net_14106) );
na02s04 TIMEBOOST_cell_37124 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_10174) );
in01s01 g58254_u0 ( .a(FE_OFN1803_n_9690), .o(g58254_sb) );
na03f02 TIMEBOOST_cell_73370 ( .a(TIMEBOOST_net_16704), .b(FE_OFN1301_n_5763), .c(g62065_sb), .o(n_7744) );
na02s01 TIMEBOOST_cell_63724 ( .a(g61992_sb), .b(g61992_db), .o(TIMEBOOST_net_20848) );
in01s01 g58255_u0 ( .a(FE_OFN543_n_9690), .o(g58255_sb) );
in01s01 TIMEBOOST_cell_64273 ( .a(TIMEBOOST_net_21128), .o(TIMEBOOST_net_21129) );
na02s01 g58255_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q), .b(FE_OFN543_n_9690), .o(g58255_db) );
in01s01 g58256_u0 ( .a(FE_OFN539_n_9690), .o(g58256_sb) );
na03f02 TIMEBOOST_cell_73569 ( .a(FE_OFN1234_n_6391), .b(TIMEBOOST_net_13394), .c(g63005_sb), .o(n_5872) );
in01s01 TIMEBOOST_cell_63575 ( .a(TIMEBOOST_net_20754), .o(TIMEBOOST_net_20755) );
in01s01 g58257_u0 ( .a(FE_OFN539_n_9690), .o(g58257_sb) );
in01s01 g58258_u0 ( .a(FE_OFN1801_n_9690), .o(g58258_sb) );
na03f02 TIMEBOOST_cell_73371 ( .a(TIMEBOOST_net_16716), .b(FE_OFN1301_n_5763), .c(g62037_sb), .o(n_7779) );
na02s01 g58258_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q), .b(FE_OFN1801_n_9690), .o(g58258_db) );
na02s01 TIMEBOOST_cell_48084 ( .a(TIMEBOOST_net_14259), .b(FE_OFN209_n_9126), .o(n_9095) );
na04f04 TIMEBOOST_cell_67681 ( .a(n_3232), .b(n_2830), .c(n_2857), .d(n_3424), .o(n_5643) );
na02f02 TIMEBOOST_cell_62904 ( .a(TIMEBOOST_net_12916), .b(n_2111), .o(TIMEBOOST_net_20399) );
in01s01 g58260_u0 ( .a(FE_OFN584_n_9692), .o(g58260_sb) );
na02s01 g58260_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q), .b(FE_OFN584_n_9692), .o(g58260_db) );
na02s01 TIMEBOOST_cell_37126 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q), .o(TIMEBOOST_net_10175) );
in01f02 g58261_u0 ( .a(FE_OFN1698_n_5751), .o(g58261_sb) );
na03f02 TIMEBOOST_cell_67976 ( .a(TIMEBOOST_net_8839), .b(FE_OFN1183_n_3476), .c(g60670_sb), .o(n_5648) );
na02f02 TIMEBOOST_cell_69895 ( .a(TIMEBOOST_net_22155), .b(g63547_db), .o(n_4610) );
in01s01 g58262_u0 ( .a(FE_OFN519_n_9697), .o(g58262_sb) );
in01s01 g58263_u0 ( .a(FE_OFN1801_n_9690), .o(g58263_sb) );
na03f02 TIMEBOOST_cell_66563 ( .a(TIMEBOOST_net_17091), .b(FE_OFN1208_n_6356), .c(g62470_sb), .o(n_6651) );
na03f02 TIMEBOOST_cell_73372 ( .a(TIMEBOOST_net_16693), .b(FE_OFN1300_n_5763), .c(g62032_sb), .o(n_7783) );
in01m01 g58264_u0 ( .a(FE_OFN1632_n_9531), .o(g58264_sb) );
na02s01 TIMEBOOST_cell_53965 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q), .o(TIMEBOOST_net_17200) );
na02f02 TIMEBOOST_cell_50216 ( .a(TIMEBOOST_net_15325), .b(g62620_sb), .o(n_6318) );
in01s01 TIMEBOOST_cell_67778 ( .a(TIMEBOOST_net_21204), .o(TIMEBOOST_net_21205) );
in01s01 g58265_u0 ( .a(FE_OFN1649_n_9428), .o(g58265_sb) );
na02s02 TIMEBOOST_cell_37900 ( .a(g58123_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q), .o(TIMEBOOST_net_10562) );
na03m02 TIMEBOOST_cell_66296 ( .a(n_3970), .b(g62844_sb), .c(g62844_db), .o(n_5283) );
in01m01 g58266_u0 ( .a(FE_OFN579_n_9531), .o(g58266_sb) );
in01s01 g58267_u0 ( .a(FE_OFN1651_n_9428), .o(g58267_sb) );
na02m02 TIMEBOOST_cell_54529 ( .a(TIMEBOOST_net_7584), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_17482) );
na04s02 TIMEBOOST_cell_46584 ( .a(TIMEBOOST_net_10788), .b(g65846_sb), .c(g61918_sb), .d(g61918_db), .o(n_7985) );
in01s01 g58268_u0 ( .a(FE_OFN602_n_9687), .o(g58268_sb) );
na02m10 TIMEBOOST_cell_49537 ( .a(g53892_sb), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in_417), .o(TIMEBOOST_net_14986) );
na02s01 g58268_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q), .b(FE_OFN602_n_9687), .o(g58268_db) );
na02m02 TIMEBOOST_cell_63171 ( .a(TIMEBOOST_net_20532), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_15488) );
in01s01 g58269_u0 ( .a(FE_OFN602_n_9687), .o(g58269_sb) );
na02m02 TIMEBOOST_cell_68672 ( .a(g65050_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q), .o(TIMEBOOST_net_21544) );
na02s01 g58269_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q), .b(FE_OFN602_n_9687), .o(g58269_db) );
in01s01 g58270_u0 ( .a(FE_OFN602_n_9687), .o(g58270_sb) );
na02m20 TIMEBOOST_cell_52193 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_140), .o(TIMEBOOST_net_16314) );
na02m01 TIMEBOOST_cell_52913 ( .a(n_6986), .b(n_13447), .o(TIMEBOOST_net_16674) );
in01m02 g58271_u0 ( .a(FE_OFN569_n_9528), .o(g58271_sb) );
na03m02 TIMEBOOST_cell_72777 ( .a(n_4465), .b(n_4323), .c(TIMEBOOST_net_12688), .o(TIMEBOOST_net_20971) );
na03f02 TIMEBOOST_cell_70318 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q), .b(FE_OFN1150_n_13249), .c(TIMEBOOST_net_12998), .o(TIMEBOOST_net_22367) );
in01s01 g58272_u0 ( .a(FE_OFN1690_n_9528), .o(g58272_sb) );
na02s02 TIMEBOOST_cell_71926 ( .a(TIMEBOOST_net_20201), .b(FE_OFN953_n_2055), .o(TIMEBOOST_net_23171) );
in01m01 g58273_u0 ( .a(FE_OFN1687_n_9528), .o(g58273_sb) );
na02m02 TIMEBOOST_cell_63121 ( .a(TIMEBOOST_net_20507), .b(FE_OFN569_n_9528), .o(TIMEBOOST_net_11462) );
na02m02 TIMEBOOST_cell_68960 ( .a(g65066_sb), .b(n_3608), .o(TIMEBOOST_net_21688) );
in01m02 g58274_u0 ( .a(FE_OFN1688_n_9528), .o(g58274_sb) );
na02m01 TIMEBOOST_cell_38926 ( .a(n_3785), .b(FE_OFN1680_n_4655), .o(TIMEBOOST_net_11075) );
na03f02 TIMEBOOST_cell_72531 ( .a(n_504), .b(n_2104), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q), .o(TIMEBOOST_net_22270) );
na02m04 TIMEBOOST_cell_68784 ( .a(g64897_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_21600) );
in01m01 g58275_u0 ( .a(FE_OFN1687_n_9528), .o(g58275_sb) );
na03f02 TIMEBOOST_cell_73160 ( .a(TIMEBOOST_net_16637), .b(FE_OFN2128_n_16497), .c(g54334_sb), .o(n_12982) );
na02f02 TIMEBOOST_cell_38969 ( .a(TIMEBOOST_net_11096), .b(FE_OFN1151_n_13249), .o(TIMEBOOST_net_345) );
in01s01 g58276_u0 ( .a(FE_OFN568_n_9528), .o(g58276_sb) );
na02s02 g58276_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN568_n_9528), .o(g58276_db) );
na02m02 TIMEBOOST_cell_44700 ( .a(TIMEBOOST_net_13244), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_11581) );
in01s01 g58277_u0 ( .a(FE_OFN568_n_9528), .o(g58277_sb) );
na02m01 TIMEBOOST_cell_38928 ( .a(n_3774), .b(FE_OFN1677_n_4655), .o(TIMEBOOST_net_11076) );
na02s02 g58277_u2 ( .a(FE_OFN215_n_9856), .b(FE_OFN568_n_9528), .o(g58277_db) );
in01s01 g58278_u0 ( .a(FE_OFN1691_n_9528), .o(g58278_sb) );
na02m02 TIMEBOOST_cell_69004 ( .a(FE_OFN612_n_4501), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q), .o(TIMEBOOST_net_21710) );
na02s02 g58278_u2 ( .a(FE_OFN217_n_9889), .b(FE_OFN1691_n_9528), .o(g58278_db) );
na02s02 TIMEBOOST_cell_39133 ( .a(TIMEBOOST_net_11178), .b(g58177_db), .o(n_9612) );
in01m02 g58279_u0 ( .a(FE_OFN1687_n_9528), .o(g58279_sb) );
no03f04 TIMEBOOST_cell_47254 ( .a(FE_RN_238_0), .b(TIMEBOOST_net_13542), .c(n_12453), .o(n_12799) );
no03f06 TIMEBOOST_cell_47255 ( .a(FE_RN_244_0), .b(TIMEBOOST_net_13543), .c(n_12453), .o(n_12795) );
in01m02 g58280_u0 ( .a(FE_OFN1690_n_9528), .o(g58280_sb) );
no03f02 TIMEBOOST_cell_47256 ( .a(FE_RN_247_0), .b(TIMEBOOST_net_8598), .c(n_12453), .o(n_12790) );
na03f02 TIMEBOOST_cell_73775 ( .a(TIMEBOOST_net_13722), .b(n_13987), .c(FE_OFN1589_n_13736), .o(n_16238) );
in01m01 g58281_u0 ( .a(FE_OFN1689_n_9528), .o(g58281_sb) );
na02m06 TIMEBOOST_cell_69007 ( .a(TIMEBOOST_net_21711), .b(g64762_sb), .o(TIMEBOOST_net_14426) );
na02m02 TIMEBOOST_cell_68873 ( .a(TIMEBOOST_net_21644), .b(TIMEBOOST_net_20196), .o(TIMEBOOST_net_17006) );
na02s01 TIMEBOOST_cell_53462 ( .a(TIMEBOOST_net_16948), .b(g58235_sb), .o(n_9556) );
in01m01 g58282_u0 ( .a(FE_OFN569_n_9528), .o(g58282_sb) );
na02s02 TIMEBOOST_cell_63120 ( .a(FE_OFN201_n_9230), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q), .o(TIMEBOOST_net_20507) );
na02m04 TIMEBOOST_cell_68474 ( .a(g64809_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q), .o(TIMEBOOST_net_21445) );
na03m04 TIMEBOOST_cell_65779 ( .a(n_13732), .b(n_16452), .c(n_4822), .o(TIMEBOOST_net_16433) );
in01s01 g58283_u0 ( .a(FE_OFN1690_n_9528), .o(g58283_sb) );
na03m04 TIMEBOOST_cell_72449 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q), .b(g58767_sb), .c(TIMEBOOST_net_14045), .o(n_9865) );
na02s02 g58283_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1690_n_9528), .o(g58283_db) );
na04f04 TIMEBOOST_cell_73297 ( .a(n_3958), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q), .c(FE_OFN2105_g64577_p), .d(g62817_sb), .o(n_5342) );
in01m02 g58284_u0 ( .a(FE_OFN1692_n_9528), .o(g58284_sb) );
in01s01 g58285_u0 ( .a(FE_OFN1690_n_9528), .o(g58285_sb) );
na03f02 TIMEBOOST_cell_73437 ( .a(TIMEBOOST_net_23333), .b(FE_OFN1222_n_6391), .c(g62365_sb), .o(n_6871) );
na03m02 TIMEBOOST_cell_64575 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q), .b(FE_OFN670_n_4505), .c(n_3744), .o(TIMEBOOST_net_16169) );
in01s01 g58286_u0 ( .a(FE_OFN1687_n_9528), .o(g58286_sb) );
na02s01 TIMEBOOST_cell_37132 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_10178) );
in01s01 g58287_u0 ( .a(FE_OFN1687_n_9528), .o(g58287_sb) );
na02m01 TIMEBOOST_cell_4276 ( .a(g52470_da), .b(FE_OFN1025_n_11877), .o(TIMEBOOST_net_698) );
na02s02 g58287_u2 ( .a(FE_OFN227_n_9841), .b(FE_OFN1687_n_9528), .o(g58287_db) );
na03f02 TIMEBOOST_cell_73712 ( .a(TIMEBOOST_net_13553), .b(n_11977), .c(FE_OFN1749_n_12004), .o(n_12675) );
in01m01 g58288_u0 ( .a(FE_OFN1688_n_9528), .o(g58288_sb) );
na02m02 TIMEBOOST_cell_4274 ( .a(g52469_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_697) );
na03m02 TIMEBOOST_cell_66347 ( .a(TIMEBOOST_net_8878), .b(g54189_sb), .c(g54189_db), .o(n_13358) );
in01m02 g58289_u0 ( .a(FE_OFN1687_n_9528), .o(g58289_sb) );
na02m20 TIMEBOOST_cell_54073 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q), .b(pci_target_unit_fifos_pciw_cbe_in_152), .o(TIMEBOOST_net_17254) );
na03m02 TIMEBOOST_cell_72779 ( .a(n_4470), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q), .c(TIMEBOOST_net_12559), .o(TIMEBOOST_net_20530) );
in01m01 g58290_u0 ( .a(FE_OFN1690_n_9528), .o(g58290_sb) );
na02m02 g58290_u2 ( .a(FE_OFN233_n_9876), .b(FE_OFN1690_n_9528), .o(g58290_db) );
na03f02 TIMEBOOST_cell_66158 ( .a(TIMEBOOST_net_17358), .b(FE_OFN1180_n_3476), .c(g60641_sb), .o(n_5688) );
in01s01 g58291_u0 ( .a(FE_OFN1690_n_9528), .o(g58291_sb) );
na03f04 TIMEBOOST_cell_66883 ( .a(TIMEBOOST_net_17184), .b(n_7213), .c(n_13127), .o(TIMEBOOST_net_13545) );
na02m02 TIMEBOOST_cell_68464 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q), .b(FE_OFN671_n_4505), .o(TIMEBOOST_net_21440) );
in01f02 g58292_u0 ( .a(FE_OFN1690_n_9528), .o(g58292_sb) );
na02f02 TIMEBOOST_cell_50596 ( .a(TIMEBOOST_net_15515), .b(g62436_sb), .o(n_6724) );
na02f01 g58292_u2 ( .a(FE_OFN235_n_9834), .b(FE_OFN1690_n_9528), .o(g58292_db) );
na02f02 TIMEBOOST_cell_38799 ( .a(TIMEBOOST_net_11011), .b(g58407_db), .o(n_9433) );
in01m01 g58293_u0 ( .a(FE_OFN1689_n_9528), .o(g58293_sb) );
na02m02 TIMEBOOST_cell_52294 ( .a(TIMEBOOST_net_16364), .b(g58381_sb), .o(n_9450) );
na03f02 TIMEBOOST_cell_66565 ( .a(n_8526), .b(wishbone_slave_unit_fifos_outGreyCount_0_), .c(n_8668), .o(n_8717) );
na03f02 TIMEBOOST_cell_73608 ( .a(TIMEBOOST_net_17465), .b(FE_OFN1285_n_4097), .c(g63187_sb), .o(n_5778) );
in01m01 g58294_u0 ( .a(FE_OFN1691_n_9528), .o(g58294_sb) );
na03f02 TIMEBOOST_cell_73454 ( .a(TIMEBOOST_net_21037), .b(FE_OFN1268_n_4095), .c(g62420_sb), .o(n_6757) );
na03f02 TIMEBOOST_cell_73373 ( .a(TIMEBOOST_net_16710), .b(FE_OFN1301_n_5763), .c(g62041_sb), .o(n_7773) );
in01s02 g58295_u0 ( .a(FE_OFN568_n_9528), .o(g58295_sb) );
na02m01 TIMEBOOST_cell_4290 ( .a(g52467_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_705) );
na02s02 g58295_u2 ( .a(FE_OFN241_n_9830), .b(FE_OFN568_n_9528), .o(g58295_db) );
in01s01 TIMEBOOST_cell_63553 ( .a(TIMEBOOST_net_20732), .o(TIMEBOOST_net_20733) );
in01m02 g58296_u0 ( .a(FE_OFN569_n_9528), .o(g58296_sb) );
na03f02 TIMEBOOST_cell_71502 ( .a(n_3005), .b(g52402_sb), .c(FE_OFN1697_n_5751), .o(TIMEBOOST_net_22959) );
na02f02 TIMEBOOST_cell_50624 ( .a(TIMEBOOST_net_15529), .b(g62542_sb), .o(n_6483) );
in01s01 TIMEBOOST_cell_63537 ( .a(TIMEBOOST_net_20716), .o(TIMEBOOST_net_20717) );
in01s01 g58297_u0 ( .a(FE_OFN568_n_9528), .o(g58297_sb) );
na02m02 TIMEBOOST_cell_69412 ( .a(g64943_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q), .o(TIMEBOOST_net_21914) );
na02f02 TIMEBOOST_cell_70963 ( .a(TIMEBOOST_net_22689), .b(g62579_sb), .o(n_6395) );
na03m02 TIMEBOOST_cell_73609 ( .a(TIMEBOOST_net_17436), .b(FE_OFN1278_n_4097), .c(g62910_sb), .o(n_6058) );
in01m01 g58298_u0 ( .a(FE_OFN569_n_9528), .o(g58298_sb) );
in01s01 TIMEBOOST_cell_73916 ( .a(wbm_dat_i_0_), .o(TIMEBOOST_net_23481) );
in01m01 g58299_u0 ( .a(FE_OFN1691_n_9528), .o(g58299_sb) );
in01s01 TIMEBOOST_cell_73937 ( .a(TIMEBOOST_net_23501), .o(TIMEBOOST_net_23502) );
na02f01 TIMEBOOST_cell_48983 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q), .b(n_12595), .o(TIMEBOOST_net_14709) );
na03f02 TIMEBOOST_cell_47175 ( .a(g53914_sb), .b(TIMEBOOST_net_13449), .c(FE_OFN1327_n_13547), .o(n_13470) );
in01m02 g58300_u0 ( .a(FE_OFN1689_n_9528), .o(g58300_sb) );
na02m02 TIMEBOOST_cell_54328 ( .a(TIMEBOOST_net_17381), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_15515) );
na02m01 TIMEBOOST_cell_37134 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q), .o(TIMEBOOST_net_10179) );
in01m01 g58301_u0 ( .a(FE_OFN1691_n_9528), .o(g58301_sb) );
na02m01 TIMEBOOST_cell_69792 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q), .o(TIMEBOOST_net_22104) );
in01s08 TIMEBOOST_cell_62384 ( .a(TIMEBOOST_net_20137), .o(FE_OFN554_n_9864) );
in01s02 g58302_u0 ( .a(FE_OFN568_n_9528), .o(g58302_sb) );
na03f02 TIMEBOOST_cell_65695 ( .a(TIMEBOOST_net_12869), .b(FE_OFN2126_n_16497), .c(g54335_sb), .o(n_12981) );
na03f02 TIMEBOOST_cell_72525 ( .a(TIMEBOOST_net_21390), .b(g64096_sb), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_22469) );
na02s01 TIMEBOOST_cell_47597 ( .a(TIMEBOOST_net_6793), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_14016) );
in01m02 g58303_u0 ( .a(FE_OFN1689_n_9528), .o(g58303_sb) );
na03f02 TIMEBOOST_cell_70732 ( .a(TIMEBOOST_net_16983), .b(FE_OCPN1911_FE_OFN1152_n_13249), .c(n_2110), .o(TIMEBOOST_net_22574) );
in01m01 g58304_u0 ( .a(FE_OFN1689_n_9528), .o(g58304_sb) );
na02s02 TIMEBOOST_cell_43310 ( .a(TIMEBOOST_net_12549), .b(g58211_sb), .o(n_9053) );
na02s02 TIMEBOOST_cell_4272 ( .a(g52465_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_696) );
na02f06 TIMEBOOST_cell_47680 ( .a(TIMEBOOST_net_14057), .b(n_1379), .o(TIMEBOOST_net_199) );
in01s01 g58305_u0 ( .a(FE_OFN569_n_9528), .o(g58305_sb) );
na03f02 TIMEBOOST_cell_73374 ( .a(TIMEBOOST_net_16705), .b(FE_OFN1301_n_5763), .c(g62052_sb), .o(n_7757) );
na04m02 TIMEBOOST_cell_67272 ( .a(g61707_sb), .b(g65697_db), .c(TIMEBOOST_net_20260), .d(TIMEBOOST_net_8194), .o(n_8413) );
in01m02 g58306_u0 ( .a(FE_OFN1687_n_9528), .o(g58306_sb) );
na03f02 TIMEBOOST_cell_65652 ( .a(TIMEBOOST_net_16633), .b(g64134_sb), .c(g64134_db), .o(TIMEBOOST_net_13070) );
na02m04 g58306_u2 ( .a(FE_OFN1687_n_9528), .b(FE_OFN254_n_9825), .o(g58306_db) );
na03s08 TIMEBOOST_cell_72420 ( .a(TIMEBOOST_net_14011), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q), .c(wbu_addr_in_266), .o(n_9853) );
in01m01 g58307_u0 ( .a(FE_OFN1657_n_9502), .o(g58307_sb) );
na02m02 TIMEBOOST_cell_68875 ( .a(TIMEBOOST_net_21645), .b(g64932_db), .o(TIMEBOOST_net_17007) );
na04s02 TIMEBOOST_cell_72880 ( .a(TIMEBOOST_net_12490), .b(g65779_sb), .c(g61767_sb), .d(g61767_db), .o(n_8277) );
in01s01 g58308_u0 ( .a(FE_OFN572_n_9502), .o(g58308_sb) );
na04f04 TIMEBOOST_cell_67968 ( .a(n_3060), .b(n_2926), .c(n_2859), .d(n_2865), .o(n_4168) );
na03m02 TIMEBOOST_cell_72815 ( .a(g65321_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q), .c(TIMEBOOST_net_16249), .o(TIMEBOOST_net_17555) );
in01s01 g58309_u0 ( .a(FE_OFN1654_n_9502), .o(g58309_sb) );
na02s01 g58309_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q), .b(g58309_sb), .o(g58309_da) );
na02m04 TIMEBOOST_cell_71878 ( .a(FE_OFN681_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q), .o(TIMEBOOST_net_23147) );
in01m02 g58310_u0 ( .a(FE_OFN1655_n_9502), .o(g58310_sb) );
na02m10 TIMEBOOST_cell_43643 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57), .b(pci_target_unit_pcit_if_strd_addr_in_693), .o(TIMEBOOST_net_12716) );
na02s02 TIMEBOOST_cell_43633 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q), .b(FE_OFN540_n_9690), .o(TIMEBOOST_net_12711) );
in01m01 g58311_u0 ( .a(FE_OFN572_n_9502), .o(g58311_sb) );
na02f01 TIMEBOOST_cell_70350 ( .a(TIMEBOOST_net_9983), .b(FE_OFN1100_g64577_p), .o(TIMEBOOST_net_22383) );
na04f02 TIMEBOOST_cell_67879 ( .a(g64792_sb), .b(n_4447), .c(n_28), .d(FE_OFN667_n_4495), .o(n_4472) );
in01s01 g58312_u0 ( .a(FE_OFN1656_n_9502), .o(g58312_sb) );
na02m01 TIMEBOOST_cell_43639 ( .a(n_6), .b(FE_OFN1628_n_4438), .o(TIMEBOOST_net_12714) );
na02s01 g58312_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN1656_n_9502), .o(g58312_db) );
na03m02 TIMEBOOST_cell_72537 ( .a(g64785_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q), .c(TIMEBOOST_net_10333), .o(TIMEBOOST_net_17481) );
in01m02 g58313_u0 ( .a(FE_OFN572_n_9502), .o(g58313_sb) );
na04f04 TIMEBOOST_cell_35026 ( .a(n_9894), .b(g57035_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q), .d(FE_OFN1407_n_8567), .o(n_11697) );
na02m02 g58313_u2 ( .a(FE_OFN217_n_9889), .b(FE_OFN572_n_9502), .o(g58313_db) );
na04f04 TIMEBOOST_cell_35027 ( .a(n_9693), .b(g57315_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q), .d(FE_OFN1376_n_8567), .o(n_11436) );
in01s01 g58314_u0 ( .a(FE_OFN1654_n_9502), .o(g58314_sb) );
na03m02 TIMEBOOST_cell_72882 ( .a(TIMEBOOST_net_12627), .b(FE_OFN1043_n_2037), .c(g65827_sb), .o(n_1889) );
na02s02 g58314_u2 ( .a(FE_OFN219_n_9853), .b(FE_OFN1654_n_9502), .o(g58314_db) );
na02m01 TIMEBOOST_cell_43645 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60), .b(pci_target_unit_pcit_if_strd_addr_in_696), .o(TIMEBOOST_net_12717) );
in01m01 g58315_u0 ( .a(FE_OFN572_n_9502), .o(g58315_sb) );
na03f02 TIMEBOOST_cell_67004 ( .a(FE_OFN1588_n_13736), .b(TIMEBOOST_net_16524), .c(FE_OCP_RBN1995_n_13971), .o(n_14300) );
in01s03 TIMEBOOST_cell_45961 ( .a(pci_target_unit_fifos_pcir_data_in_188), .o(TIMEBOOST_net_13922) );
in01m01 g58316_u0 ( .a(FE_OFN572_n_9502), .o(g58316_sb) );
na02m01 TIMEBOOST_cell_43635 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q), .o(TIMEBOOST_net_12712) );
na03f04 TIMEBOOST_cell_67001 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_16518), .c(FE_OFN1587_n_13736), .o(g53301_p) );
in01s02 g58317_u0 ( .a(FE_OFN1657_n_9502), .o(g58317_sb) );
na02s01 TIMEBOOST_cell_37140 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q), .b(pci_target_unit_fifos_pcir_data_in_165), .o(TIMEBOOST_net_10182) );
in01s01 g58318_u0 ( .a(FE_OFN1656_n_9502), .o(g58318_sb) );
na02m01 TIMEBOOST_cell_4300 ( .a(g52463_da), .b(FE_OFN1022_n_11877), .o(TIMEBOOST_net_710) );
na02s02 g58318_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1656_n_9502), .o(g58318_db) );
in01m01 g58319_u0 ( .a(FE_OFN572_n_9502), .o(g58319_sb) );
na04f04 TIMEBOOST_cell_35028 ( .a(n_9674), .b(g57256_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q), .d(FE_OFN1376_n_8567), .o(n_11497) );
na02m02 g58319_u2 ( .a(FE_OFN223_n_9844), .b(FE_OFN572_n_9502), .o(g58319_db) );
na04f04 TIMEBOOST_cell_35029 ( .a(n_9719), .b(g57215_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q), .d(FE_OFN1384_n_8567), .o(n_11543) );
in01s01 g58320_u0 ( .a(FE_OFN572_n_9502), .o(g58320_sb) );
na02m08 TIMEBOOST_cell_43629 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q), .o(TIMEBOOST_net_12709) );
na02s01 g58320_u2 ( .a(FE_OFN225_n_9122), .b(FE_OFN572_n_9502), .o(g58320_db) );
na02m02 TIMEBOOST_cell_43631 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_122), .o(TIMEBOOST_net_12710) );
in01m01 g58321_u0 ( .a(FE_OFN1654_n_9502), .o(g58321_sb) );
na02f02 TIMEBOOST_cell_62868 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q), .b(FE_OFN712_n_8140), .o(TIMEBOOST_net_20381) );
na02m01 TIMEBOOST_cell_68506 ( .a(g65710_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_21461) );
na02f01 TIMEBOOST_cell_53553 ( .a(FE_OFN1094_g64577_p), .b(g62733_sb), .o(TIMEBOOST_net_16994) );
in01s01 g58322_u0 ( .a(FE_OFN1654_n_9502), .o(g58322_sb) );
na03m06 TIMEBOOST_cell_66786 ( .a(TIMEBOOST_net_16669), .b(FE_OFN1119_g64577_p), .c(g63043_sb), .o(n_5166) );
na02m10 TIMEBOOST_cell_45771 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q), .o(TIMEBOOST_net_13780) );
in01m01 g58323_u0 ( .a(FE_OFN1655_n_9502), .o(g58323_sb) );
na04s02 TIMEBOOST_cell_72918 ( .a(g61734_sb), .b(g61734_db), .c(g65691_db), .d(TIMEBOOST_net_10338), .o(n_8351) );
na02f02 TIMEBOOST_cell_50340 ( .a(TIMEBOOST_net_15387), .b(g62353_sb), .o(n_6895) );
in01m01 g58324_u0 ( .a(FE_OFN572_n_9502), .o(g58324_sb) );
na02s01 TIMEBOOST_cell_53327 ( .a(TIMEBOOST_net_6822), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q), .o(TIMEBOOST_net_16881) );
in01s01 g58325_u0 ( .a(FE_OFN572_n_9502), .o(g58325_sb) );
na04f04 TIMEBOOST_cell_35222 ( .a(n_10942), .b(n_9286), .c(n_10099), .d(n_9287), .o(n_17041) );
na03f02 TIMEBOOST_cell_67003 ( .a(FE_OFN1588_n_13736), .b(TIMEBOOST_net_16526), .c(FE_OCP_RBN1995_n_13971), .o(n_14260) );
na02s01 TIMEBOOST_cell_68238 ( .a(pci_inta_oe_o), .b(g63590_sb), .o(TIMEBOOST_net_21327) );
in01s01 g58326_u0 ( .a(FE_OFN1657_n_9502), .o(g58326_sb) );
na02s01 g58326_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q), .b(g58326_sb), .o(g58326_da) );
na02f02 TIMEBOOST_cell_70537 ( .a(TIMEBOOST_net_22476), .b(g63182_sb), .o(n_4945) );
na03m02 TIMEBOOST_cell_71924 ( .a(FE_OFN662_n_4392), .b(g65076_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q), .o(TIMEBOOST_net_23170) );
in01s01 g58327_u0 ( .a(FE_OFN572_n_9502), .o(g58327_sb) );
na04f02 TIMEBOOST_cell_35224 ( .a(n_10660), .b(n_10931), .c(n_10661), .d(n_12441), .o(n_12774) );
na02m02 TIMEBOOST_cell_4296 ( .a(g52461_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_708) );
in01s01 g58328_u0 ( .a(FE_OFN572_n_9502), .o(g58328_sb) );
na02s01 TIMEBOOST_cell_49286 ( .a(TIMEBOOST_net_14860), .b(TIMEBOOST_net_10864), .o(TIMEBOOST_net_10015) );
in01s01 g58329_u0 ( .a(FE_OFN1656_n_9502), .o(g58329_sb) );
na02s01 g58329_u2 ( .a(FE_OFN241_n_9830), .b(FE_OFN1656_n_9502), .o(g58329_db) );
in01s01 g58330_u0 ( .a(FE_OFN1657_n_9502), .o(g58330_sb) );
na04f04 TIMEBOOST_cell_35030 ( .a(n_9028), .b(g57439_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q), .d(FE_OFN1405_n_8567), .o(n_10353) );
na02s01 g58330_u2 ( .a(FE_OFN201_n_9230), .b(FE_OFN1657_n_9502), .o(g58330_db) );
in01m02 g58331_u0 ( .a(FE_OFN1656_n_9502), .o(g58331_sb) );
na02f02 TIMEBOOST_cell_69975 ( .a(TIMEBOOST_net_22195), .b(FE_OFN713_n_8140), .o(TIMEBOOST_net_15804) );
na02s04 g58331_u2 ( .a(FE_OFN203_n_9228), .b(FE_OFN1656_n_9502), .o(g58331_db) );
in01s01 TIMEBOOST_cell_73881 ( .a(TIMEBOOST_net_23445), .o(TIMEBOOST_net_23446) );
in01m01 g58332_u0 ( .a(FE_OFN1657_n_9502), .o(g58332_sb) );
na03m02 TIMEBOOST_cell_73161 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q), .b(g64322_sb), .c(TIMEBOOST_net_22320), .o(TIMEBOOST_net_13109) );
in01s01 g58333_u0 ( .a(FE_OFN1657_n_9502), .o(g58333_sb) );
na02s02 g58333_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q), .b(g58333_sb), .o(g58333_da) );
na02s01 TIMEBOOST_cell_37781 ( .a(TIMEBOOST_net_10502), .b(g57954_db), .o(n_9854) );
in01m02 g58334_u0 ( .a(FE_OFN1654_n_9502), .o(g58334_sb) );
na04m06 TIMEBOOST_cell_67182 ( .a(n_3739), .b(FE_OFN634_n_4454), .c(g65030_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q), .o(n_3627) );
in01s01 g58335_u0 ( .a(FE_OFN572_n_9502), .o(g58335_sb) );
na03f02 TIMEBOOST_cell_73162 ( .a(n_1880), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q), .c(FE_OFN707_n_8119), .o(TIMEBOOST_net_14813) );
na02s02 g58335_u2 ( .a(FE_OFN243_n_9116), .b(FE_OFN572_n_9502), .o(g58335_db) );
na02m01 TIMEBOOST_cell_43617 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_124), .o(TIMEBOOST_net_12703) );
in01s01 g58336_u0 ( .a(FE_OFN1656_n_9502), .o(g58336_sb) );
na02m01 TIMEBOOST_cell_43619 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_139), .o(TIMEBOOST_net_12704) );
na02s01 g58336_u2 ( .a(FE_OFN245_n_9114), .b(FE_OFN1656_n_9502), .o(g58336_db) );
na04m08 TIMEBOOST_cell_67184 ( .a(g64905_sb), .b(FE_OFN624_n_4409), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q), .d(n_4447), .o(n_4406) );
in01m02 g58337_u0 ( .a(FE_OFN1655_n_9502), .o(g58337_sb) );
na03s01 TIMEBOOST_cell_41702 ( .a(g58440_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q), .c(TIMEBOOST_net_8741), .o(n_9411) );
in01m01 g58338_u0 ( .a(FE_OFN1654_n_9502), .o(g58338_sb) );
na02m02 TIMEBOOST_cell_69137 ( .a(TIMEBOOST_net_21776), .b(TIMEBOOST_net_14414), .o(TIMEBOOST_net_17376) );
na04f04 TIMEBOOST_cell_73503 ( .a(n_2170), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q), .c(FE_OFN706_n_8119), .d(g62006_sb), .o(n_7883) );
na03f02 TIMEBOOST_cell_66920 ( .a(FE_OFN1551_n_12104), .b(TIMEBOOST_net_16492), .c(FE_OCP_RBN1979_n_10273), .o(n_12508) );
in01m02 g58339_u0 ( .a(FE_OFN1657_n_9502), .o(g58339_sb) );
na02s02 g58339_u2 ( .a(FE_OFN252_n_9868), .b(FE_OFN1657_n_9502), .o(g58339_db) );
na02s01 TIMEBOOST_cell_45359 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q), .o(TIMEBOOST_net_13574) );
in01s01 g58340_u0 ( .a(FE_OFN1654_n_9502), .o(g58340_sb) );
na02s02 g58340_u2 ( .a(FE_OFN254_n_9825), .b(FE_OFN1654_n_9502), .o(g58340_db) );
na02s01 TIMEBOOST_cell_43615 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q), .b(FE_OFN539_n_9690), .o(TIMEBOOST_net_12702) );
in01m02 g58341_u0 ( .a(FE_OFN1670_n_9477), .o(g58341_sb) );
na02f02 TIMEBOOST_cell_44688 ( .a(TIMEBOOST_net_13238), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_11623) );
na02f01 TIMEBOOST_cell_62446 ( .a(n_2648), .b(g65994_sb), .o(TIMEBOOST_net_20170) );
in01s01 g58342_u0 ( .a(FE_OFN1666_n_9477), .o(g58342_sb) );
na02m02 TIMEBOOST_cell_4294 ( .a(g52460_da), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_707) );
na03m02 TIMEBOOST_cell_64574 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q), .b(FE_OFN670_n_4505), .c(n_3747), .o(TIMEBOOST_net_16165) );
in01s01 g58343_u0 ( .a(FE_OFN1666_n_9477), .o(g58343_sb) );
na03m06 TIMEBOOST_cell_72720 ( .a(g64918_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q), .c(TIMEBOOST_net_14282), .o(TIMEBOOST_net_17455) );
na04f04 TIMEBOOST_cell_73298 ( .a(n_4733), .b(n_366), .c(FE_OFN1127_g64577_p), .d(g63035_sb), .o(n_7126) );
na03f02 TIMEBOOST_cell_73553 ( .a(TIMEBOOST_net_20583), .b(FE_OFN1235_n_6391), .c(g62656_sb), .o(n_6231) );
in01s01 g58344_u0 ( .a(FE_OFN1668_n_9477), .o(g58344_sb) );
na03m02 TIMEBOOST_cell_72939 ( .a(pci_target_unit_del_sync_addr_in_231), .b(g65213_sb), .c(TIMEBOOST_net_7160), .o(n_2674) );
na03m06 TIMEBOOST_cell_68730 ( .a(TIMEBOOST_net_17214), .b(FE_OFN917_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q), .o(TIMEBOOST_net_21573) );
na02s01 TIMEBOOST_cell_63754 ( .a(FE_OFN1648_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q), .o(TIMEBOOST_net_20863) );
in01s01 g58345_u0 ( .a(FE_OFN1666_n_9477), .o(g58345_sb) );
na04f04 TIMEBOOST_cell_72642 ( .a(TIMEBOOST_net_21483), .b(g53939_sb), .c(wishbone_slave_unit_pcim_if_wbw_cbe_in_416), .d(FE_OFN1083_n_13221), .o(TIMEBOOST_net_23362) );
no03f02 TIMEBOOST_cell_66934 ( .a(FE_OCP_RBN2292_FE_OFN1575_n_12028), .b(TIMEBOOST_net_16499), .c(FE_OCPN1895_FE_OFN1559_n_12042), .o(n_12709) );
in01s01 g58346_u0 ( .a(FE_OFN548_n_9477), .o(g58346_sb) );
na02s01 g58346_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN548_n_9477), .o(g58346_db) );
na03f02 TIMEBOOST_cell_72940 ( .a(pci_target_unit_del_sync_addr_in_217), .b(g65219_sb), .c(TIMEBOOST_net_7140), .o(n_2668) );
in01s01 g58347_u0 ( .a(FE_OFN548_n_9477), .o(g58347_sb) );
na02f10 TIMEBOOST_cell_68093 ( .a(TIMEBOOST_net_21254), .b(n_783), .o(n_11877) );
in01m01 g58348_u0 ( .a(FE_OFN1671_n_9477), .o(g58348_sb) );
na02s01 TIMEBOOST_cell_53237 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in), .o(TIMEBOOST_net_16836) );
na02m02 g58348_u2 ( .a(FE_OFN217_n_9889), .b(FE_OFN1671_n_9477), .o(g58348_db) );
na03f02 TIMEBOOST_cell_73375 ( .a(TIMEBOOST_net_16712), .b(FE_OFN1300_n_5763), .c(g62062_sb), .o(n_7747) );
in01s01 g58349_u0 ( .a(FE_OFN1666_n_9477), .o(g58349_sb) );
na03f02 TIMEBOOST_cell_72941 ( .a(pci_target_unit_del_sync_addr_in_222), .b(g65244_sb), .c(TIMEBOOST_net_7156), .o(n_2638) );
na02s01 g58349_u2 ( .a(FE_OFN219_n_9853), .b(FE_OFN1666_n_9477), .o(g58349_db) );
na03s02 TIMEBOOST_cell_64358 ( .a(g61962_db), .b(g61962_sb), .c(wbs_dat_i_1_), .o(TIMEBOOST_net_14689) );
in01m10 g58350_u0 ( .a(FE_OFN1666_n_9477), .o(g58350_sb) );
na02s01 TIMEBOOST_cell_68498 ( .a(pci_target_unit_del_sync_addr_in_219), .b(g66403_sb), .o(TIMEBOOST_net_21457) );
na03f02 TIMEBOOST_cell_34935 ( .a(TIMEBOOST_net_9524), .b(FE_OFN1390_n_8567), .c(g57531_sb), .o(n_11211) );
na02m02 TIMEBOOST_cell_53626 ( .a(TIMEBOOST_net_17030), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_15539) );
in01m02 g58351_u0 ( .a(FE_OFN1670_n_9477), .o(g58351_sb) );
na02f02 TIMEBOOST_cell_54642 ( .a(TIMEBOOST_net_17538), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_15516) );
in01s01 g58352_u0 ( .a(FE_OFN1666_n_9477), .o(g58352_sb) );
na02f02 TIMEBOOST_cell_70325 ( .a(TIMEBOOST_net_22370), .b(g61697_sb), .o(n_6980) );
na02m01 TIMEBOOST_cell_4286 ( .a(g52458_da), .b(FE_OFN1023_n_11877), .o(TIMEBOOST_net_703) );
in01s01 g58353_u0 ( .a(FE_OFN1668_n_9477), .o(g58353_sb) );
na03f02 TIMEBOOST_cell_72942 ( .a(pci_target_unit_del_sync_addr_in_230), .b(g65217_sb), .c(TIMEBOOST_net_7162), .o(n_2670) );
in01s01 g58354_u0 ( .a(FE_OFN1666_n_9477), .o(g58354_sb) );
na03f02 TIMEBOOST_cell_72943 ( .a(pci_target_unit_del_sync_addr_in_228), .b(g65221_sb), .c(TIMEBOOST_net_7143), .o(n_2666) );
na02s01 g58354_u2 ( .a(FE_OFN225_n_9122), .b(FE_OFN1666_n_9477), .o(g58354_db) );
na03m10 TIMEBOOST_cell_64355 ( .a(n_1196), .b(n_1383), .c(n_1551), .o(TIMEBOOST_net_10177) );
in01s01 g58355_u0 ( .a(FE_OFN1666_n_9477), .o(g58355_sb) );
na02f02 TIMEBOOST_cell_70449 ( .a(TIMEBOOST_net_22432), .b(n_7216), .o(n_7624) );
na03f02 TIMEBOOST_cell_73554 ( .a(TIMEBOOST_net_17513), .b(FE_OFN1236_n_6391), .c(g62601_sb), .o(n_6348) );
in01s01 g58356_u0 ( .a(FE_OFN1666_n_9477), .o(g58356_sb) );
na03m02 TIMEBOOST_cell_72593 ( .a(TIMEBOOST_net_21438), .b(g64779_sb), .c(TIMEBOOST_net_21654), .o(TIMEBOOST_net_17471) );
na02s01 g58356_u2 ( .a(FE_OFN227_n_9841), .b(FE_OFN1666_n_9477), .o(g58356_db) );
na03f02 TIMEBOOST_cell_71168 ( .a(TIMEBOOST_net_17474), .b(n_13221), .c(FE_OFN2070_n_15978), .o(TIMEBOOST_net_22792) );
in01s01 g58357_u0 ( .a(FE_OFN1668_n_9477), .o(g58357_sb) );
na04f04 TIMEBOOST_cell_73094 ( .a(g65919_db), .b(TIMEBOOST_net_12630), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q), .d(FE_OFN719_n_8060), .o(TIMEBOOST_net_15046) );
na03f01 TIMEBOOST_cell_65080 ( .a(n_3770), .b(TIMEBOOST_net_12590), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q), .o(TIMEBOOST_net_16778) );
na02f02 TIMEBOOST_cell_30310 ( .a(TIMEBOOST_net_9259), .b(n_7317), .o(n_8535) );
in01s01 g58358_u0 ( .a(FE_OFN1666_n_9477), .o(g58358_sb) );
na02s01 TIMEBOOST_cell_63118 ( .a(FE_OFN1789_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q), .o(TIMEBOOST_net_20506) );
na03m02 TIMEBOOST_cell_72810 ( .a(TIMEBOOST_net_21614), .b(g64931_sb), .c(TIMEBOOST_net_21841), .o(TIMEBOOST_net_16786) );
na03s02 TIMEBOOST_cell_46415 ( .a(TIMEBOOST_net_12607), .b(g57980_sb), .c(TIMEBOOST_net_12738), .o(TIMEBOOST_net_9418) );
in01s01 g58359_u0 ( .a(FE_OFN1666_n_9477), .o(g58359_sb) );
in01s01 g58360_u0 ( .a(FE_OFN1666_n_9477), .o(g58360_sb) );
na04f04 TIMEBOOST_cell_36036 ( .a(n_662), .b(g63195_sb), .c(TIMEBOOST_net_5664), .d(g53939_db), .o(n_13506) );
na03m02 TIMEBOOST_cell_72816 ( .a(g65317_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q), .c(TIMEBOOST_net_14373), .o(TIMEBOOST_net_17371) );
na02m04 TIMEBOOST_cell_68481 ( .a(TIMEBOOST_net_21448), .b(TIMEBOOST_net_20204), .o(n_9884) );
in01s01 g58361_u0 ( .a(FE_OFN1666_n_9477), .o(g58361_sb) );
na02m10 TIMEBOOST_cell_52669 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q), .o(TIMEBOOST_net_16552) );
in01s01 TIMEBOOST_cell_67726 ( .a(TIMEBOOST_net_21152), .o(TIMEBOOST_net_21153) );
in01s01 g58362_u0 ( .a(FE_OFN1668_n_9477), .o(g58362_sb) );
na02m01 TIMEBOOST_cell_4284 ( .a(g52457_da), .b(FE_OFN1025_n_11877), .o(TIMEBOOST_net_702) );
na02m02 TIMEBOOST_cell_63303 ( .a(TIMEBOOST_net_20598), .b(FE_OFN1687_n_9528), .o(TIMEBOOST_net_12976) );
in01m01 g58363_u0 ( .a(FE_OFN1668_n_9477), .o(g58363_sb) );
na02m01 TIMEBOOST_cell_62790 ( .a(n_4473), .b(n_26), .o(TIMEBOOST_net_20342) );
na02f01 TIMEBOOST_cell_48984 ( .a(TIMEBOOST_net_14709), .b(FE_OFN2127_n_16497), .o(TIMEBOOST_net_323) );
na02s01 TIMEBOOST_cell_38411 ( .a(TIMEBOOST_net_10817), .b(g58020_db), .o(n_9770) );
in01s01 g58364_u0 ( .a(FE_OFN548_n_9477), .o(g58364_sb) );
na03s01 TIMEBOOST_cell_72365 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_70), .b(wishbone_slave_unit_pci_initiator_if_data_source), .c(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_8632) );
na03f01 TIMEBOOST_cell_65070 ( .a(n_3777), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q), .c(FE_OFN612_n_4501), .o(TIMEBOOST_net_14453) );
in01m01 g58365_u0 ( .a(FE_OFN1671_n_9477), .o(g58365_sb) );
na03f02 TIMEBOOST_cell_73438 ( .a(TIMEBOOST_net_20605), .b(FE_OFN1215_n_4151), .c(g62448_sb), .o(n_6701) );
na02m02 TIMEBOOST_cell_69139 ( .a(TIMEBOOST_net_21777), .b(g64963_db), .o(TIMEBOOST_net_17385) );
na02s01 TIMEBOOST_cell_48909 ( .a(FE_OFN535_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q), .o(TIMEBOOST_net_14672) );
in01f02 g58366_u0 ( .a(FE_OFN1670_n_9477), .o(g58366_sb) );
na02m06 TIMEBOOST_cell_69006 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q), .b(FE_OFN1663_n_4490), .o(TIMEBOOST_net_21711) );
na04m10 TIMEBOOST_cell_67801 ( .a(pci_target_unit_pci_target_sm_n_2), .b(pci_target_unit_pci_target_sm_n_3), .c(n_976), .d(g66457_sb), .o(n_1134) );
na02s01 g58367_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q), .b(FE_OFN1669_n_9477), .o(g58367_da) );
na03s01 TIMEBOOST_cell_72572 ( .a(pci_target_unit_del_sync_addr_in_224), .b(g66403_sb), .c(g66407_db), .o(n_2531) );
na02f01 TIMEBOOST_cell_69790 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q), .o(TIMEBOOST_net_22103) );
in01m02 g58368_u0 ( .a(FE_OFN1668_n_9477), .o(g58368_sb) );
na03f02 TIMEBOOST_cell_65323 ( .a(TIMEBOOST_net_8276), .b(n_5633), .c(g62101_sb), .o(n_5601) );
na02s01 TIMEBOOST_cell_49737 ( .a(FE_OFN561_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q), .o(TIMEBOOST_net_15086) );
in01s01 g58369_u0 ( .a(FE_OFN1667_n_9477), .o(g58369_sb) );
na02s01 g58369_u2 ( .a(FE_OFN1667_n_9477), .b(FE_OFN243_n_9116), .o(g58369_db) );
na03s02 TIMEBOOST_cell_64981 ( .a(g65780_db), .b(TIMEBOOST_net_6914), .c(TIMEBOOST_net_8201), .o(n_8400) );
in01s01 g58370_u0 ( .a(FE_OFN548_n_9477), .o(g58370_sb) );
na02f02 TIMEBOOST_cell_68377 ( .a(TIMEBOOST_net_21396), .b(g64203_sb), .o(TIMEBOOST_net_13062) );
na02s01 g58370_u2 ( .a(FE_OFN548_n_9477), .b(FE_OFN245_n_9114), .o(g58370_db) );
na03f02 TIMEBOOST_cell_72781 ( .a(n_4488), .b(n_4280), .c(TIMEBOOST_net_12592), .o(TIMEBOOST_net_20964) );
in01m01 g58371_u0 ( .a(FE_OFN1668_n_9477), .o(g58371_sb) );
na02s02 TIMEBOOST_cell_49447 ( .a(g58239_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q), .o(TIMEBOOST_net_14941) );
na02s01 g58371_u2 ( .a(FE_OFN247_n_9112), .b(FE_OFN1668_n_9477), .o(g58371_db) );
na02f01 TIMEBOOST_cell_52299 ( .a(TIMEBOOST_net_12732), .b(FE_OFN1033_n_4732), .o(TIMEBOOST_net_16367) );
in01s01 g58372_u0 ( .a(FE_OFN1668_n_9477), .o(g58372_sb) );
na03f02 TIMEBOOST_cell_73299 ( .a(TIMEBOOST_net_13056), .b(FE_OFN1122_g64577_p), .c(g63024_sb), .o(n_5198) );
na03f02 TIMEBOOST_cell_73776 ( .a(TIMEBOOST_net_8112), .b(n_13987), .c(FE_OFN1588_n_13736), .o(n_16229) );
in01f02 g58373_u0 ( .a(FE_OFN1670_n_9477), .o(g58373_sb) );
na02m02 TIMEBOOST_cell_53648 ( .a(TIMEBOOST_net_17041), .b(g62549_sb), .o(n_6468) );
na02m02 TIMEBOOST_cell_68483 ( .a(TIMEBOOST_net_21449), .b(g65099_sb), .o(TIMEBOOST_net_17430) );
in01s01 g58374_u0 ( .a(FE_OFN1666_n_9477), .o(g58374_sb) );
na02s01 g58374_u2 ( .a(FE_OFN254_n_9825), .b(FE_OFN1666_n_9477), .o(g58374_db) );
na04f04 TIMEBOOST_cell_73455 ( .a(n_4905), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q), .c(FE_OFN1222_n_6391), .d(g62512_sb), .o(n_7381) );
in01f06 g58375_u0 ( .a(FE_OFN1635_n_9531), .o(g58375_sb) );
na03f02 TIMEBOOST_cell_73300 ( .a(TIMEBOOST_net_13077), .b(FE_OFN1128_g64577_p), .c(g63551_sb), .o(n_4926) );
na02f06 g58375_u2 ( .a(FE_OFN1635_n_9531), .b(FE_OFN207_n_9865), .o(g58375_db) );
na02s01 TIMEBOOST_cell_45793 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q), .o(TIMEBOOST_net_13791) );
in01m01 g58376_u0 ( .a(FE_OFN580_n_9531), .o(g58376_sb) );
na02s01 TIMEBOOST_cell_43621 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q), .o(TIMEBOOST_net_12705) );
na02f06 TIMEBOOST_cell_52696 ( .a(TIMEBOOST_net_16565), .b(n_1973), .o(n_2492) );
na02m02 TIMEBOOST_cell_37087 ( .a(TIMEBOOST_net_10155), .b(g67057_sb), .o(n_1685) );
in01s01 g58377_u0 ( .a(FE_OFN579_n_9531), .o(g58377_sb) );
na03m02 TIMEBOOST_cell_72964 ( .a(pci_target_unit_del_sync_addr_in_234), .b(g65231_sb), .c(TIMEBOOST_net_5417), .o(n_2656) );
in01m02 g58378_u0 ( .a(FE_OFN1632_n_9531), .o(g58378_sb) );
na02m02 TIMEBOOST_cell_43597 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(g65747_sb), .o(TIMEBOOST_net_12693) );
in01m01 g58379_u0 ( .a(FE_OFN580_n_9531), .o(g58379_sb) );
na03f04 TIMEBOOST_cell_66768 ( .a(TIMEBOOST_net_17140), .b(FE_OFN1313_n_6624), .c(g63160_sb), .o(n_5816) );
na03f02 TIMEBOOST_cell_65272 ( .a(TIMEBOOST_net_16932), .b(FE_OFN1055_n_4727), .c(g64260_sb), .o(TIMEBOOST_net_13097) );
in01m02 g58380_u0 ( .a(FE_OFN1634_n_9531), .o(g58380_sb) );
na03f02 TIMEBOOST_cell_34860 ( .a(TIMEBOOST_net_9323), .b(FE_OFN1397_n_8567), .c(g57037_sb), .o(n_10515) );
na02s02 g58380_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN1634_n_9531), .o(g58380_db) );
na02s02 TIMEBOOST_cell_68282 ( .a(g65695_sb), .b(TIMEBOOST_net_21203), .o(TIMEBOOST_net_21349) );
in01m01 g58381_u0 ( .a(FE_OFN1634_n_9531), .o(g58381_sb) );
na03f02 TIMEBOOST_cell_47401 ( .a(FE_OFN1586_n_13736), .b(TIMEBOOST_net_13711), .c(FE_OCP_RBN1999_n_13971), .o(n_14419) );
na02s01 TIMEBOOST_cell_51531 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_15983) );
in01m01 g58382_u0 ( .a(FE_OFN1631_n_9531), .o(g58382_sb) );
na02f02 TIMEBOOST_cell_70579 ( .a(TIMEBOOST_net_22497), .b(g63123_sb), .o(n_5009) );
na02m02 g58382_u1 ( .a(g58382_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q), .o(g58382_da) );
in01s01 g58383_u0 ( .a(FE_OFN579_n_9531), .o(g58383_sb) );
na02s02 TIMEBOOST_cell_44180 ( .a(TIMEBOOST_net_12984), .b(g58244_sb), .o(n_9548) );
na03m02 TIMEBOOST_cell_72783 ( .a(TIMEBOOST_net_21547), .b(g65721_sb), .c(FE_OFN717_n_8176), .o(TIMEBOOST_net_22202) );
na02s02 TIMEBOOST_cell_44181 ( .a(FE_OFN268_n_9880), .b(g58083_sb), .o(TIMEBOOST_net_12985) );
in01m02 g58384_u0 ( .a(FE_OFN580_n_9531), .o(g58384_sb) );
na02m01 TIMEBOOST_cell_69190 ( .a(TIMEBOOST_net_12443), .b(FE_OFN928_n_4730), .o(TIMEBOOST_net_21803) );
in01f01 g58385_u0 ( .a(FE_OFN580_n_9531), .o(g58385_sb) );
na03m02 TIMEBOOST_cell_72638 ( .a(g64900_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q), .c(TIMEBOOST_net_16180), .o(TIMEBOOST_net_17375) );
na04m04 TIMEBOOST_cell_65484 ( .a(n_2194), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q), .c(FE_OFN699_n_7845), .d(g61731_sb), .o(n_8358) );
in01f01 g58386_u0 ( .a(FE_OFN1635_n_9531), .o(g58386_sb) );
in01s01 TIMEBOOST_cell_64272 ( .a(pci_target_unit_fifos_pcir_data_in_186), .o(TIMEBOOST_net_21128) );
na03f02 TIMEBOOST_cell_73222 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_1_), .b(g60407_sb), .c(TIMEBOOST_net_5465), .o(n_4860) );
in01s01 g58387_u0 ( .a(FE_OFN1635_n_9531), .o(g58387_sb) );
na03f02 TIMEBOOST_cell_73376 ( .a(TIMEBOOST_net_16699), .b(FE_OFN1299_n_5763), .c(g62055_sb), .o(n_7754) );
na02s02 g58387_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1635_n_9531), .o(g58387_db) );
na02s01 TIMEBOOST_cell_44182 ( .a(TIMEBOOST_net_12985), .b(g58083_db), .o(n_9712) );
in01m01 g58388_u0 ( .a(FE_OFN580_n_9531), .o(g58388_sb) );
na03m02 TIMEBOOST_cell_72563 ( .a(TIMEBOOST_net_23134), .b(FE_OFN630_n_4454), .c(TIMEBOOST_net_21505), .o(TIMEBOOST_net_17137) );
na02m02 g58388_u2 ( .a(FE_OFN580_n_9531), .b(FE_OFN223_n_9844), .o(g58388_db) );
na02f02 TIMEBOOST_cell_69965 ( .a(TIMEBOOST_net_22190), .b(g64321_sb), .o(TIMEBOOST_net_15057) );
in01s01 g58389_u0 ( .a(FE_OFN580_n_9531), .o(g58389_sb) );
na03f02 TIMEBOOST_cell_66428 ( .a(TIMEBOOST_net_20611), .b(FE_OFN1320_n_6436), .c(g62576_sb), .o(n_7377) );
na02m01 g58389_u2 ( .a(FE_OFN580_n_9531), .b(FE_OFN225_n_9122), .o(g58389_db) );
na02m02 TIMEBOOST_cell_68793 ( .a(TIMEBOOST_net_21604), .b(TIMEBOOST_net_10541), .o(TIMEBOOST_net_17363) );
in01m02 g58390_u0 ( .a(FE_OFN579_n_9531), .o(g58390_sb) );
na03f02 TIMEBOOST_cell_73814 ( .a(TIMEBOOST_net_13778), .b(FE_OFN1775_n_13800), .c(FE_OFN1769_n_14054), .o(n_14510) );
in01s01 TIMEBOOST_cell_73882 ( .a(n_7943), .o(TIMEBOOST_net_23447) );
in01s01 g58391_u0 ( .a(FE_OFN579_n_9531), .o(g58391_sb) );
na02s02 g58391_u2 ( .a(FE_OFN227_n_9841), .b(FE_OFN579_n_9531), .o(g58391_db) );
na03f02 TIMEBOOST_cell_66663 ( .a(TIMEBOOST_net_17115), .b(FE_OFN1314_n_6624), .c(g62571_sb), .o(n_6413) );
in01m02 g58392_u0 ( .a(FE_OFN1632_n_9531), .o(g58392_sb) );
na03f02 TIMEBOOST_cell_66318 ( .a(TIMEBOOST_net_17050), .b(n_6645), .c(g63003_sb), .o(n_5876) );
na02m02 TIMEBOOST_cell_70073 ( .a(TIMEBOOST_net_22244), .b(g61727_sb), .o(n_8366) );
na02f01 TIMEBOOST_cell_68265 ( .a(TIMEBOOST_net_21340), .b(n_14070), .o(TIMEBOOST_net_503) );
in01m02 g58393_u0 ( .a(FE_OFN580_n_9531), .o(g58393_sb) );
na03s01 TIMEBOOST_cell_41706 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q), .b(g58312_sb), .c(g58312_db), .o(n_9025) );
in01s01 g58394_u0 ( .a(FE_OFN1635_n_9531), .o(g58394_sb) );
na02m01 g58394_u2 ( .a(FE_OFN270_n_9836), .b(FE_OFN1635_n_9531), .o(g58394_db) );
in01m01 g58395_u0 ( .a(FE_OFN580_n_9531), .o(g58395_sb) );
na03f01 TIMEBOOST_cell_69196 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(FE_OFN928_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q), .o(TIMEBOOST_net_21806) );
na02f01 g58395_u2 ( .a(FE_OFN235_n_9834), .b(FE_OFN580_n_9531), .o(g58395_db) );
na04f02 TIMEBOOST_cell_67685 ( .a(n_14746), .b(n_14839), .c(g52448_sb), .d(n_3425), .o(n_14844) );
in01m01 g58396_u0 ( .a(FE_OFN580_n_9531), .o(g58396_sb) );
na03f02 TIMEBOOST_cell_66664 ( .a(TIMEBOOST_net_17002), .b(FE_OFN1285_n_4097), .c(g62566_sb), .o(n_6425) );
na02m10 TIMEBOOST_cell_72036 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_149), .o(TIMEBOOST_net_23226) );
in01s01 g58397_u0 ( .a(FE_OFN580_n_9531), .o(g58397_sb) );
na02m02 TIMEBOOST_cell_72261 ( .a(TIMEBOOST_net_23338), .b(g62966_sb), .o(n_5950) );
na02m01 g58397_u2 ( .a(FE_OFN580_n_9531), .b(FE_OFN239_n_9832), .o(g58397_db) );
na02s01 TIMEBOOST_cell_45695 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q), .o(TIMEBOOST_net_13742) );
in01m01 g58398_u0 ( .a(FE_OFN1634_n_9531), .o(g58398_sb) );
na04f04 TIMEBOOST_cell_24820 ( .a(n_10081), .b(n_9280), .c(n_10084), .d(n_9283), .o(n_11846) );
in01s01 TIMEBOOST_cell_73944 ( .a(wbm_dat_i_22_), .o(TIMEBOOST_net_23509) );
na03f02 TIMEBOOST_cell_67005 ( .a(FE_OFN1588_n_13736), .b(TIMEBOOST_net_16525), .c(FE_OCP_RBN1995_n_13971), .o(g53207_p) );
in01s01 g58399_u0 ( .a(FE_OFN1631_n_9531), .o(g58399_sb) );
na02s01 g58399_u2 ( .a(FE_OFN201_n_9230), .b(FE_OFN1631_n_9531), .o(g58399_db) );
na02m02 TIMEBOOST_cell_69141 ( .a(TIMEBOOST_net_21778), .b(TIMEBOOST_net_10634), .o(TIMEBOOST_net_17563) );
in01m01 g58400_u0 ( .a(FE_OFN1634_n_9531), .o(g58400_sb) );
na02s02 g58400_u2 ( .a(FE_OFN203_n_9228), .b(FE_OFN1634_n_9531), .o(g58400_db) );
na04s02 TIMEBOOST_cell_35727 ( .a(g57899_sb), .b(FE_OFN205_n_9140), .c(g57899_db), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q), .o(TIMEBOOST_net_9478) );
in01f01 g58401_u0 ( .a(FE_OFN1631_n_9531), .o(g58401_sb) );
na02m01 TIMEBOOST_cell_52179 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_16307) );
in01s01 TIMEBOOST_cell_67792 ( .a(TIMEBOOST_net_21219), .o(TIMEBOOST_net_21218) );
na02m02 g58401_u2 ( .a(FE_OFN205_n_9140), .b(FE_OFN1631_n_9531), .o(g58401_db) );
in01s01 g58402_u0 ( .a(FE_OFN1631_n_9531), .o(g58402_sb) );
na03m02 TIMEBOOST_cell_72577 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q), .b(FE_OFN660_n_4392), .c(TIMEBOOST_net_21679), .o(TIMEBOOST_net_17548) );
in01f02 g58403_u0 ( .a(FE_OFN579_n_9531), .o(g58403_sb) );
na03f02 TIMEBOOST_cell_73163 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q), .b(g64324_sb), .c(g64324_db), .o(n_3852) );
na02f02 TIMEBOOST_cell_49354 ( .a(TIMEBOOST_net_14894), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_5472) );
in01s01 g58404_u0 ( .a(FE_OFN580_n_9531), .o(g58404_sb) );
na02s01 TIMEBOOST_cell_45697 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q), .o(TIMEBOOST_net_13743) );
na02s02 g58404_u2 ( .a(FE_OFN243_n_9116), .b(FE_OFN580_n_9531), .o(g58404_db) );
in01m01 g58405_u0 ( .a(FE_OFN1634_n_9531), .o(g58405_sb) );
na02f02 TIMEBOOST_cell_70075 ( .a(TIMEBOOST_net_22245), .b(g64973_db), .o(TIMEBOOST_net_20961) );
na02s02 g58405_u2 ( .a(FE_OFN245_n_9114), .b(FE_OFN1634_n_9531), .o(g58405_db) );
na04f10 TIMEBOOST_cell_73223 ( .a(TIMEBOOST_net_14986), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q), .c(FE_OFN1147_n_13249), .d(g54164_sb), .o(g53893_da) );
in01m02 g58406_u0 ( .a(FE_OFN1632_n_9531), .o(g58406_sb) );
in01f02 g58407_u0 ( .a(FE_OFN1635_n_9531), .o(g58407_sb) );
na02f02 TIMEBOOST_cell_50206 ( .a(TIMEBOOST_net_15320), .b(g62691_sb), .o(n_6164) );
na02f02 g58407_u2 ( .a(FE_OFN1635_n_9531), .b(FE_OFN252_n_9868), .o(g58407_db) );
na04m08 TIMEBOOST_cell_67187 ( .a(n_3741), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q), .c(FE_OFN625_n_4409), .d(g65044_sb), .o(n_3623) );
in01s01 g58408_u0 ( .a(FE_OFN579_n_9531), .o(g58408_sb) );
na02m10 TIMEBOOST_cell_45699 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_13744) );
na02m04 TIMEBOOST_cell_72234 ( .a(FE_OFN247_n_9112), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q), .o(TIMEBOOST_net_23325) );
in01s01 g58409_u0 ( .a(FE_OFN1656_n_9502), .o(g58409_sb) );
na02s02 TIMEBOOST_cell_53265 ( .a(FE_OFN564_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q), .o(TIMEBOOST_net_16850) );
na03m02 TIMEBOOST_cell_46590 ( .a(TIMEBOOST_net_12631), .b(g64276_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q), .o(TIMEBOOST_net_12895) );
na03f02 TIMEBOOST_cell_73795 ( .a(TIMEBOOST_net_13749), .b(FE_OFN1601_n_13995), .c(FE_OFN1605_n_13997), .o(n_14441) );
in01s01 g58410_u0 ( .a(FE_OFN519_n_9697), .o(g58410_sb) );
na02m04 TIMEBOOST_cell_72033 ( .a(TIMEBOOST_net_23224), .b(TIMEBOOST_net_14454), .o(TIMEBOOST_net_13363) );
na02s01 g58410_u2 ( .a(FE_OFN519_n_9697), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q), .o(g58410_db) );
na02f02 TIMEBOOST_cell_50612 ( .a(TIMEBOOST_net_15523), .b(g63164_sb), .o(n_5808) );
in01s01 g58411_u0 ( .a(FE_OFN518_n_9697), .o(g58411_sb) );
na02f02 TIMEBOOST_cell_70573 ( .a(TIMEBOOST_net_22494), .b(g62730_sb), .o(n_5519) );
na02s01 g58411_u2 ( .a(FE_OFN518_n_9697), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q), .o(g58411_db) );
na02m02 TIMEBOOST_cell_70937 ( .a(TIMEBOOST_net_22676), .b(g63166_sb), .o(n_5806) );
in01s01 g58412_u0 ( .a(FE_OFN587_n_9692), .o(g58412_sb) );
na02s01 TIMEBOOST_cell_43081 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q), .o(TIMEBOOST_net_12435) );
na02s02 g58412_u2 ( .a(FE_OFN587_n_9692), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q), .o(g58412_db) );
in01s01 g58413_u0 ( .a(FE_OFN589_n_9692), .o(g58413_sb) );
na02m10 TIMEBOOST_cell_68095 ( .a(TIMEBOOST_net_21255), .b(n_2316), .o(TIMEBOOST_net_195) );
na02s01 g58413_u2 ( .a(FE_OFN589_n_9692), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q), .o(g58413_db) );
in01s01 g58414_u0 ( .a(FE_OFN587_n_9692), .o(g58414_sb) );
na04f04 TIMEBOOST_cell_73224 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in), .b(TIMEBOOST_net_7274), .c(FE_OFN1148_n_13249), .d(g54234_sb), .o(n_13441) );
na02f02 TIMEBOOST_cell_71100 ( .a(TIMEBOOST_net_17029), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_22758) );
na02s01 TIMEBOOST_cell_45069 ( .a(g58448_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q), .o(TIMEBOOST_net_13429) );
in01s01 g58415_u0 ( .a(FE_OFN595_n_9694), .o(g58415_sb) );
in01s01 TIMEBOOST_cell_31881 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .o(TIMEBOOST_net_10045) );
na02s01 g58415_u2 ( .a(FE_OFN595_n_9694), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q), .o(g58415_db) );
in01s01 g58416_u0 ( .a(FE_OFN597_n_9694), .o(g58416_sb) );
na02s01 TIMEBOOST_cell_47792 ( .a(TIMEBOOST_net_14113), .b(FE_OFN519_n_9697), .o(TIMEBOOST_net_10350) );
na02s01 g58416_u2 ( .a(FE_OFN597_n_9694), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q), .o(g58416_db) );
in01s01 g58417_u0 ( .a(FE_OFN595_n_9694), .o(g58417_sb) );
na02f02 TIMEBOOST_cell_72227 ( .a(TIMEBOOST_net_23321), .b(g63096_sb), .o(n_5062) );
na02s01 TIMEBOOST_cell_42807 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_12298) );
na02f02 TIMEBOOST_cell_70587 ( .a(TIMEBOOST_net_22501), .b(g62766_sb), .o(n_5463) );
in01m01 g58418_u0 ( .a(FE_OFN1655_n_9502), .o(g58418_sb) );
na02s01 TIMEBOOST_cell_45701 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q), .o(TIMEBOOST_net_13745) );
na03f02 TIMEBOOST_cell_73570 ( .a(TIMEBOOST_net_17510), .b(FE_OFN1231_n_6391), .c(g62909_sb), .o(n_6060) );
na02s02 TIMEBOOST_cell_53267 ( .a(g58308_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q), .o(TIMEBOOST_net_16851) );
in01s01 g58419_u0 ( .a(FE_OFN1651_n_9428), .o(g58419_sb) );
na02s01 TIMEBOOST_cell_45703 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q), .o(TIMEBOOST_net_13746) );
na02m02 TIMEBOOST_cell_50294 ( .a(TIMEBOOST_net_15364), .b(g62661_sb), .o(n_6221) );
in01s01 g58420_u0 ( .a(FE_OFN1650_n_9428), .o(g58420_sb) );
na02m01 TIMEBOOST_cell_47598 ( .a(TIMEBOOST_net_14016), .b(n_2299), .o(TIMEBOOST_net_12301) );
in01s01 g58421_u0 ( .a(FE_OFN523_n_9428), .o(g58421_sb) );
na02s01 g58421_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q), .b(g58421_sb), .o(g58421_da) );
na03m02 TIMEBOOST_cell_73301 ( .a(TIMEBOOST_net_22317), .b(FE_OFN701_n_7845), .c(g61911_sb), .o(n_7999) );
na02f02 TIMEBOOST_cell_70975 ( .a(TIMEBOOST_net_22695), .b(g62665_sb), .o(n_6208) );
in01m10 g58422_u0 ( .a(FE_OFN1648_n_9428), .o(g58422_sb) );
na02s02 TIMEBOOST_cell_63223 ( .a(TIMEBOOST_net_20558), .b(FE_OFN252_n_9868), .o(TIMEBOOST_net_10853) );
in01s01 g58423_u0 ( .a(FE_OFN1650_n_9428), .o(g58423_sb) );
na03f02 TIMEBOOST_cell_73302 ( .a(TIMEBOOST_net_13063), .b(FE_OFN877_g64577_p), .c(g63130_sb), .o(n_4991) );
na02s01 g58423_u2 ( .a(FE_OFN213_n_9124), .b(FE_OFN1650_n_9428), .o(g58423_db) );
in01s01 g58424_u0 ( .a(FE_OFN1650_n_9428), .o(g58424_sb) );
na03s02 TIMEBOOST_cell_72579 ( .a(n_2544), .b(g66398_sb), .c(g66398_db), .o(n_2545) );
na03m02 TIMEBOOST_cell_47143 ( .a(TIMEBOOST_net_13386), .b(g54188_sb), .c(g54188_db), .o(n_13427) );
in01s01 g58425_u0 ( .a(FE_OFN523_n_9428), .o(g58425_sb) );
na02s01 TIMEBOOST_cell_45705 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_13747) );
na02s01 g58425_u2 ( .a(FE_OFN219_n_9853), .b(FE_OFN523_n_9428), .o(g58425_db) );
na02s02 TIMEBOOST_cell_53271 ( .a(g58254_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q), .o(TIMEBOOST_net_16853) );
in01s01 g58426_u0 ( .a(FE_OFN1648_n_9428), .o(g58426_sb) );
na02m02 TIMEBOOST_cell_70389 ( .a(TIMEBOOST_net_22402), .b(g58128_sb), .o(TIMEBOOST_net_20453) );
na02f02 TIMEBOOST_cell_29437 ( .a(configuration_wb_err_addr_553), .b(FE_OFN1174_n_5592), .o(TIMEBOOST_net_8823) );
na02s01 TIMEBOOST_cell_38210 ( .a(g58322_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q), .o(TIMEBOOST_net_10717) );
in01s01 g58427_u0 ( .a(FE_OFN1649_n_9428), .o(g58427_sb) );
na02m02 TIMEBOOST_cell_62825 ( .a(TIMEBOOST_net_20359), .b(FE_OFN1037_n_4732), .o(TIMEBOOST_net_14744) );
na02s01 TIMEBOOST_cell_45707 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q), .o(TIMEBOOST_net_13748) );
in01s01 g58428_u0 ( .a(FE_OFN1650_n_9428), .o(g58428_sb) );
na02f02 TIMEBOOST_cell_53273 ( .a(wbu_addr_in_258), .b(n_2740), .o(TIMEBOOST_net_16854) );
na02s01 g58428_u2 ( .a(FE_OFN221_n_9846), .b(FE_OFN1650_n_9428), .o(g58428_db) );
na02f02 TIMEBOOST_cell_53275 ( .a(n_2226), .b(wbu_addr_in_256), .o(TIMEBOOST_net_16855) );
in01s01 g58429_u0 ( .a(FE_OFN1649_n_9428), .o(g58429_sb) );
na02m10 TIMEBOOST_cell_45715 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q), .o(TIMEBOOST_net_13752) );
na02f04 TIMEBOOST_cell_53277 ( .a(wbu_addr_in_277), .b(n_3471), .o(TIMEBOOST_net_16856) );
in01s01 g58430_u0 ( .a(FE_OFN1648_n_9428), .o(g58430_sb) );
na02s01 TIMEBOOST_cell_45717 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_13753) );
na02s01 g58430_u2 ( .a(FE_OFN1648_n_9428), .b(FE_OFN225_n_9122), .o(g58430_db) );
na02f02 TIMEBOOST_cell_53279 ( .a(wbu_addr_in_261), .b(n_2719), .o(TIMEBOOST_net_16857) );
in01s01 g58431_u0 ( .a(FE_OFN1648_n_9428), .o(g58431_sb) );
na02s01 TIMEBOOST_cell_45719 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q), .o(TIMEBOOST_net_13754) );
na02m02 TIMEBOOST_cell_62578 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q), .b(n_3764), .o(TIMEBOOST_net_20236) );
na02f02 TIMEBOOST_cell_53281 ( .a(wbu_addr_in_260), .b(n_2695), .o(TIMEBOOST_net_16858) );
in01s01 g58432_u0 ( .a(FE_OFN1649_n_9428), .o(g58432_sb) );
na04s02 TIMEBOOST_cell_67189 ( .a(g58046_sb), .b(g58061_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q), .d(FE_OFN272_n_9828), .o(TIMEBOOST_net_9496) );
na03m02 TIMEBOOST_cell_72814 ( .a(n_4452), .b(FE_OFN639_n_4669), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q), .o(TIMEBOOST_net_23288) );
in01s01 g58433_u0 ( .a(FE_OFN1648_n_9428), .o(g58433_sb) );
na02s01 TIMEBOOST_cell_45721 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q), .o(TIMEBOOST_net_13755) );
na02f02 TIMEBOOST_cell_70516 ( .a(TIMEBOOST_net_13094), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_22466) );
in01s01 g58434_u0 ( .a(FE_OFN1650_n_9428), .o(g58434_sb) );
na02s01 g58434_u1 ( .a(g58434_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q), .o(g58434_da) );
na02f04 TIMEBOOST_cell_53283 ( .a(wbu_addr_in_273), .b(n_3332), .o(TIMEBOOST_net_16859) );
na02f02 TIMEBOOST_cell_53285 ( .a(wbu_addr_in_276), .b(n_3465), .o(TIMEBOOST_net_16860) );
in01s01 g58435_u0 ( .a(FE_OFN1648_n_9428), .o(g58435_sb) );
na02m08 TIMEBOOST_cell_38113 ( .a(TIMEBOOST_net_10668), .b(g64273_db), .o(n_3900) );
in01s01 g58436_u0 ( .a(FE_OFN1649_n_9428), .o(g58436_sb) );
in01s01 g58437_u0 ( .a(FE_OFN1650_n_9428), .o(g58437_sb) );
na02f02 TIMEBOOST_cell_53316 ( .a(FE_RN_496_0), .b(TIMEBOOST_net_16875), .o(FE_RN_498_0) );
na02s02 TIMEBOOST_cell_37940 ( .a(g58319_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q), .o(TIMEBOOST_net_10582) );
na02f06 g54489_u1 ( .a(g54489_sb), .b(TIMEBOOST_net_13885), .o(g54489_da) );
in01s02 g58438_u0 ( .a(FE_OFN1651_n_9428), .o(g58438_sb) );
na02f01 TIMEBOOST_cell_62419 ( .a(TIMEBOOST_net_20156), .b(n_16424), .o(TIMEBOOST_net_16141) );
na02s02 g58438_u2 ( .a(FE_OFN201_n_9230), .b(FE_OFN1651_n_9428), .o(g58438_db) );
na02s01 TIMEBOOST_cell_45070 ( .a(TIMEBOOST_net_13429), .b(g58448_db), .o(n_9197) );
in01s01 g58439_u0 ( .a(FE_OFN1650_n_9428), .o(g58439_sb) );
na02f02 TIMEBOOST_cell_70977 ( .a(TIMEBOOST_net_22696), .b(g62443_sb), .o(n_6709) );
na02s01 g58439_u2 ( .a(FE_OFN203_n_9228), .b(FE_OFN1650_n_9428), .o(g58439_db) );
in01s01 g58440_u0 ( .a(FE_OFN1651_n_9428), .o(g58440_sb) );
na03f02 TIMEBOOST_cell_73713 ( .a(n_12010), .b(TIMEBOOST_net_13566), .c(FE_OFN1748_n_12004), .o(n_12512) );
na03f02 TIMEBOOST_cell_73050 ( .a(TIMEBOOST_net_16624), .b(FE_OFN2079_n_8069), .c(g62071_sb), .o(n_7826) );
in01s02 g58441_u0 ( .a(FE_OFN523_n_9428), .o(g58441_sb) );
na03m02 TIMEBOOST_cell_65569 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q), .b(n_4450), .c(TIMEBOOST_net_12823), .o(TIMEBOOST_net_17397) );
na03f02 TIMEBOOST_cell_73225 ( .a(TIMEBOOST_net_23295), .b(TIMEBOOST_net_10918), .c(FE_OFN1276_n_4096), .o(TIMEBOOST_net_22703) );
in01s01 g58442_u0 ( .a(FE_OFN1650_n_9428), .o(g58442_sb) );
na02f02 TIMEBOOST_cell_50682 ( .a(TIMEBOOST_net_15558), .b(g62832_sb), .o(n_5311) );
na02f02 TIMEBOOST_cell_50680 ( .a(TIMEBOOST_net_15557), .b(g62759_sb), .o(n_5472) );
in01s01 g58443_u0 ( .a(FE_OFN1649_n_9428), .o(g58443_sb) );
na02f06 TIMEBOOST_cell_53320 ( .a(TIMEBOOST_net_16877), .b(FE_RN_270_0), .o(TIMEBOOST_net_10222) );
na03f02 TIMEBOOST_cell_66567 ( .a(TIMEBOOST_net_17099), .b(FE_OFN1312_n_6624), .c(g62599_sb), .o(n_6353) );
in01s01 g58444_u0 ( .a(FE_OFN523_n_9428), .o(g58444_sb) );
na03f02 TIMEBOOST_cell_73377 ( .a(TIMEBOOST_net_16715), .b(FE_OFN1301_n_5763), .c(g62050_sb), .o(n_7760) );
na02f01 TIMEBOOST_cell_62988 ( .a(conf_wb_err_addr_in_956), .b(g62116_sb), .o(TIMEBOOST_net_20441) );
in01s01 g58445_u0 ( .a(FE_OFN523_n_9428), .o(g58445_sb) );
na02f04 TIMEBOOST_cell_53319 ( .a(FE_RN_269_0), .b(FE_RN_271_0), .o(TIMEBOOST_net_16877) );
na04m06 TIMEBOOST_cell_72836 ( .a(n_3770), .b(g64780_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q), .d(g64780_db), .o(TIMEBOOST_net_17551) );
na02s01 TIMEBOOST_cell_49285 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q), .b(g58424_sb), .o(TIMEBOOST_net_14860) );
in01s01 g58446_u0 ( .a(FE_OFN1801_n_9690), .o(g58446_sb) );
na02m02 TIMEBOOST_cell_48850 ( .a(TIMEBOOST_net_14642), .b(FE_OFN1691_n_9528), .o(TIMEBOOST_net_11082) );
na02s01 g58446_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q), .b(FE_OFN1801_n_9690), .o(g58446_db) );
na03f04 TIMEBOOST_cell_67009 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_16523), .c(FE_OFN1587_n_13736), .o(g53255_p) );
in01s01 g58447_u0 ( .a(FE_OFN543_n_9690), .o(g58447_sb) );
na02s01 g58447_u2 ( .a(FE_OFN543_n_9690), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q), .o(g58447_db) );
na02s02 TIMEBOOST_cell_51316 ( .a(TIMEBOOST_net_15875), .b(TIMEBOOST_net_10872), .o(TIMEBOOST_net_9489) );
in01s01 g58448_u0 ( .a(FE_OFN548_n_9477), .o(g58448_sb) );
na02f04 TIMEBOOST_cell_53287 ( .a(wbu_addr_in_266), .b(n_3346), .o(TIMEBOOST_net_16861) );
na02s01 g58448_u2 ( .a(FE_OFN548_n_9477), .b(FE_OFN203_n_9228), .o(g58448_db) );
in01s01 g58449_u0 ( .a(FE_OFN1648_n_9428), .o(g58449_sb) );
na03f02 TIMEBOOST_cell_34819 ( .a(TIMEBOOST_net_9381), .b(FE_OFN1404_n_8567), .c(g57090_sb), .o(n_11651) );
in01s01 g58450_u0 ( .a(FE_OFN1648_n_9428), .o(g58450_sb) );
na03f02 TIMEBOOST_cell_66708 ( .a(TIMEBOOST_net_17127), .b(FE_OFN1320_n_6436), .c(g62998_sb), .o(n_5886) );
na02f02 TIMEBOOST_cell_53289 ( .a(wbu_addr_in_263), .b(n_3358), .o(TIMEBOOST_net_16862) );
in01s01 g58451_u0 ( .a(FE_OFN1649_n_9428), .o(g58451_sb) );
na02m10 TIMEBOOST_cell_45777 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q), .o(TIMEBOOST_net_13783) );
in01s01 g58452_u0 ( .a(FE_OFN1651_n_9428), .o(g58452_sb) );
na02m10 TIMEBOOST_cell_45779 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q), .o(TIMEBOOST_net_13784) );
na02s01 g58452_u2 ( .a(FE_OFN252_n_9868), .b(FE_OFN1651_n_9428), .o(g58452_db) );
in01s01 g58453_u0 ( .a(FE_OFN1651_n_9428), .o(g58453_sb) );
na04f04 TIMEBOOST_cell_67689 ( .a(TIMEBOOST_net_16865), .b(FE_OFN2200_n_10256), .c(g52605_sb), .d(TIMEBOOST_net_705), .o(n_11866) );
na04f04 TIMEBOOST_cell_67691 ( .a(TIMEBOOST_net_16860), .b(FE_OFN2200_n_10256), .c(g52611_sb), .d(TIMEBOOST_net_704), .o(n_11860) );
in01s01 g58454_u0 ( .a(FE_OFN1649_n_9428), .o(g58454_sb) );
na02m10 TIMEBOOST_cell_45781 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q), .o(TIMEBOOST_net_13785) );
in01f02 g58455_u0 ( .a(FE_OFN1437_n_9372), .o(g58455_sb) );
in01s01 TIMEBOOST_cell_31882 ( .a(TIMEBOOST_net_10045), .o(TIMEBOOST_net_10046) );
in01s01 TIMEBOOST_cell_46001 ( .a(wbu_sel_in), .o(TIMEBOOST_net_13962) );
na02f06 TIMEBOOST_cell_3652 ( .a(n_15918), .b(n_15908), .o(TIMEBOOST_net_386) );
in01f02 g58456_u0 ( .a(FE_OFN1436_n_9372), .o(g58456_sb) );
na02f08 TIMEBOOST_cell_3653 ( .a(FE_RN_895_0), .b(TIMEBOOST_net_386), .o(n_16520) );
na02s01 TIMEBOOST_cell_48088 ( .a(TIMEBOOST_net_14261), .b(FE_OFN223_n_9844), .o(TIMEBOOST_net_9321) );
in01f02 g58457_u0 ( .a(FE_OFN1440_n_9372), .o(g58457_sb) );
na04f04 TIMEBOOST_cell_73672 ( .a(n_3863), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q), .c(FE_OFN1122_g64577_p), .d(g63103_sb), .o(n_5048) );
na02f06 TIMEBOOST_cell_3656 ( .a(n_2753), .b(n_1355), .o(TIMEBOOST_net_388) );
in01f02 g58458_u0 ( .a(FE_OFN1440_n_9372), .o(g58458_sb) );
na02f08 TIMEBOOST_cell_3657 ( .a(TIMEBOOST_net_388), .b(n_3189), .o(n_3190) );
na02s01 TIMEBOOST_cell_43448 ( .a(TIMEBOOST_net_12618), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_10781) );
in01f02 g58459_u0 ( .a(FE_OFN1439_n_9372), .o(g58459_sb) );
na02s01 TIMEBOOST_cell_43450 ( .a(TIMEBOOST_net_12619), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_10782) );
in01f02 g58460_u0 ( .a(FE_OFN1436_n_9372), .o(g58460_sb) );
na02f04 TIMEBOOST_cell_53291 ( .a(wbu_addr_in_264), .b(n_3133), .o(TIMEBOOST_net_16863) );
in01f02 g58461_u0 ( .a(FE_OFN1436_n_9372), .o(g58461_sb) );
na03f02 TIMEBOOST_cell_47327 ( .a(FE_OFN1572_n_11027), .b(TIMEBOOST_net_13617), .c(FE_OFN1752_n_12086), .o(n_12679) );
na02m10 TIMEBOOST_cell_53193 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68), .b(pci_target_unit_pcit_if_strd_addr_in_704), .o(TIMEBOOST_net_16814) );
na02s01 TIMEBOOST_cell_30999 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_26__Q), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_9604) );
in01f02 g58462_u0 ( .a(FE_OFN1436_n_9372), .o(g58462_sb) );
na02s01 TIMEBOOST_cell_44035 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q), .b(g58265_sb), .o(TIMEBOOST_net_12912) );
na02f02 TIMEBOOST_cell_3665 ( .a(TIMEBOOST_net_392), .b(n_7626), .o(n_8487) );
na03f02 TIMEBOOST_cell_24839 ( .a(n_10865), .b(FE_RN_143_0), .c(n_12562), .o(n_12824) );
in01f02 g58463_u0 ( .a(FE_OFN1441_n_9372), .o(g58463_sb) );
na02f10 TIMEBOOST_cell_3667 ( .a(TIMEBOOST_net_393), .b(g54131_da), .o(n_13679) );
na03f02 TIMEBOOST_cell_72681 ( .a(TIMEBOOST_net_16590), .b(FE_OFN789_n_2678), .c(g65242_sb), .o(n_2640) );
in01f02 g58464_u0 ( .a(FE_OFN1439_n_9372), .o(g58464_sb) );
na02s01 TIMEBOOST_cell_68053 ( .a(TIMEBOOST_net_21234), .b(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_10137) );
na03f06 TIMEBOOST_cell_65704 ( .a(TIMEBOOST_net_16949), .b(FE_OFN2128_n_16497), .c(g54333_sb), .o(n_12983) );
in01f02 g58465_u0 ( .a(FE_OFN1441_n_9372), .o(g58465_sb) );
na03f02 TIMEBOOST_cell_65947 ( .a(TIMEBOOST_net_16405), .b(FE_OFN1171_n_5592), .c(g62137_sb), .o(n_5556) );
in01s01 TIMEBOOST_cell_73968 ( .a(wbm_dat_i_4_), .o(TIMEBOOST_net_23533) );
in01s01 TIMEBOOST_cell_46004 ( .a(TIMEBOOST_net_13965), .o(TIMEBOOST_net_13964) );
in01f02 g58466_u0 ( .a(FE_OFN1437_n_9372), .o(g58466_sb) );
na03f02 TIMEBOOST_cell_34798 ( .a(TIMEBOOST_net_9548), .b(FE_OFN1397_n_8567), .c(g57051_sb), .o(n_10509) );
na03f02 TIMEBOOST_cell_67013 ( .a(FE_OFN1586_n_13736), .b(n_13993), .c(TIMEBOOST_net_13723), .o(n_14415) );
na02s01 TIMEBOOST_cell_3674 ( .a(n_16818), .b(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q), .o(TIMEBOOST_net_397) );
in01f02 g58467_u0 ( .a(FE_OFN1436_n_9372), .o(g58467_sb) );
na03s02 TIMEBOOST_cell_73095 ( .a(TIMEBOOST_net_22059), .b(g65894_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q), .o(TIMEBOOST_net_22199) );
na02f02 TIMEBOOST_cell_3675 ( .a(n_8596), .b(TIMEBOOST_net_397), .o(n_8680) );
na02f01 TIMEBOOST_cell_44554 ( .a(TIMEBOOST_net_13171), .b(g62790_sb), .o(n_5409) );
in01f02 g58468_u0 ( .a(FE_OFN1441_n_9372), .o(g58468_sb) );
na03f02 TIMEBOOST_cell_73485 ( .a(TIMEBOOST_net_22597), .b(g58800_db), .c(TIMEBOOST_net_22779), .o(n_14824) );
na04f04 TIMEBOOST_cell_36867 ( .a(TIMEBOOST_net_9619), .b(FE_OFN2200_n_10256), .c(g52610_sb), .d(TIMEBOOST_net_709), .o(n_11861) );
na03f02 TIMEBOOST_cell_34698 ( .a(n_4065), .b(g62735_sb), .c(TIMEBOOST_net_7700), .o(n_5509) );
in01f02 g58469_u0 ( .a(FE_OFN1439_n_9372), .o(g58469_sb) );
na04f02 TIMEBOOST_cell_25255 ( .a(n_14296), .b(n_14011), .c(n_13862), .d(n_14567), .o(n_14612) );
na02m02 TIMEBOOST_cell_69704 ( .a(g65382_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q), .o(TIMEBOOST_net_22060) );
na03m02 TIMEBOOST_cell_72744 ( .a(n_4479), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q), .c(TIMEBOOST_net_12546), .o(TIMEBOOST_net_17067) );
in01f02 g58470_u0 ( .a(FE_OFN1439_n_9372), .o(g58470_sb) );
na02m02 TIMEBOOST_cell_69692 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q), .b(FE_OFN1678_n_4655), .o(TIMEBOOST_net_22054) );
na02s01 TIMEBOOST_cell_17995 ( .a(g58773_sb), .b(wbu_addr_in_264), .o(TIMEBOOST_net_5361) );
in01f02 g58471_u0 ( .a(FE_OFN1440_n_9372), .o(g58471_sb) );
na02s01 TIMEBOOST_cell_37146 ( .a(n_9904), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q), .o(TIMEBOOST_net_10185) );
na02s01 TIMEBOOST_cell_48171 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q), .b(FE_OFN585_n_9692), .o(TIMEBOOST_net_14303) );
na03f01 TIMEBOOST_cell_68206 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q), .b(FE_OFN276_n_9941), .c(TIMEBOOST_net_8590), .o(TIMEBOOST_net_21311) );
in01f02 g58472_u0 ( .a(FE_OFN1440_n_9372), .o(g58472_sb) );
in01s01 TIMEBOOST_cell_63554 ( .a(TIMEBOOST_net_20734), .o(wbs_adr_i_19_) );
na04m04 TIMEBOOST_cell_67468 ( .a(TIMEBOOST_net_20353), .b(FE_OFN1628_n_4438), .c(g65015_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q), .o(TIMEBOOST_net_13369) );
no04f80 TIMEBOOST_cell_64291 ( .a(FE_RN_731_0), .b(parchk_pci_ad_out_in_1174), .c(parchk_pci_ad_out_in_1173), .d(FE_RN_732_0), .o(n_585) );
in01f02 g58473_u0 ( .a(FE_OFN1441_n_9372), .o(g58473_sb) );
na03f02 TIMEBOOST_cell_73226 ( .a(TIMEBOOST_net_14593), .b(FE_OFN2081_n_8176), .c(g61751_sb), .o(n_8313) );
na02m01 TIMEBOOST_cell_69148 ( .a(n_4452), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q), .o(TIMEBOOST_net_21782) );
na02f08 TIMEBOOST_cell_3688 ( .a(n_4743), .b(n_2742), .o(TIMEBOOST_net_404) );
in01f02 g58474_u0 ( .a(FE_OFN1439_n_9372), .o(g58474_sb) );
na03f01 TIMEBOOST_cell_21132 ( .a(pci_target_unit_fifos_pcir_whole_waddr_94), .b(n_8503), .c(FE_OFN2079_n_8069), .o(n_8505) );
na02f08 TIMEBOOST_cell_3689 ( .a(TIMEBOOST_net_404), .b(n_7110), .o(n_8465) );
na02f02 TIMEBOOST_cell_3690 ( .a(n_4743), .b(n_2308), .o(TIMEBOOST_net_405) );
in01f02 g58475_u0 ( .a(FE_OFN1436_n_9372), .o(g58475_sb) );
na02s01 TIMEBOOST_cell_31015 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_22__Q), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_9612) );
na02f08 TIMEBOOST_cell_3691 ( .a(TIMEBOOST_net_405), .b(n_7110), .o(n_8512) );
na02m02 TIMEBOOST_cell_70159 ( .a(TIMEBOOST_net_22287), .b(g64221_sb), .o(n_3948) );
in01f02 g58476_u0 ( .a(FE_OFN1438_n_9372), .o(g58476_sb) );
na02m02 TIMEBOOST_cell_69431 ( .a(TIMEBOOST_net_21923), .b(TIMEBOOST_net_16238), .o(TIMEBOOST_net_17147) );
na02s02 TIMEBOOST_cell_52405 ( .a(FE_OFN243_n_9116), .b(g58132_sb), .o(TIMEBOOST_net_16420) );
in01f02 g58477_u0 ( .a(FE_OFN1440_n_9372), .o(g58477_sb) );
in01s01 TIMEBOOST_cell_45940 ( .a(TIMEBOOST_net_13901), .o(TIMEBOOST_net_13900) );
na02f04 TIMEBOOST_cell_3695 ( .a(TIMEBOOST_net_407), .b(n_13625), .o(n_13821) );
na02s01 TIMEBOOST_cell_3696 ( .a(n_7530), .b(n_7044), .o(TIMEBOOST_net_408) );
in01f02 g58478_u0 ( .a(FE_OFN1438_n_9372), .o(g58478_sb) );
na02s01 TIMEBOOST_cell_51707 ( .a(n_384), .b(n_255), .o(TIMEBOOST_net_16071) );
na02f04 TIMEBOOST_cell_3697 ( .a(TIMEBOOST_net_408), .b(n_13625), .o(n_13810) );
na02f10 TIMEBOOST_cell_17964 ( .a(TIMEBOOST_net_5345), .b(FE_RN_209_0), .o(n_1535) );
in01f02 g58479_u0 ( .a(FE_OFN1436_n_9372), .o(g58479_sb) );
in01s01 TIMEBOOST_cell_67774 ( .a(TIMEBOOST_net_21200), .o(TIMEBOOST_net_21201) );
in01f02 g58480_u0 ( .a(FE_OFN1440_n_9372), .o(g58480_sb) );
no03f04 TIMEBOOST_cell_73695 ( .a(n_4649), .b(n_12595), .c(n_4877), .o(g59347_p) );
na02f06 g54176_u1 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_396), .b(g54176_sb), .o(g54176_da) );
in01f02 g58481_u0 ( .a(FE_OFN1438_n_9372), .o(g58481_sb) );
na02f02 TIMEBOOST_cell_71361 ( .a(TIMEBOOST_net_22888), .b(n_5232), .o(n_13414) );
na02s01 TIMEBOOST_cell_31001 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_20__Q), .b(FE_OFN221_n_9846), .o(TIMEBOOST_net_9605) );
in01f02 g58482_u0 ( .a(FE_OFN1439_n_9372), .o(g58482_sb) );
na02f02 TIMEBOOST_cell_3705 ( .a(TIMEBOOST_net_412), .b(n_13828), .o(n_14087) );
in01f02 g58483_u0 ( .a(FE_OFN1440_n_9372), .o(g58483_sb) );
na02s01 TIMEBOOST_cell_48322 ( .a(TIMEBOOST_net_14378), .b(FE_OFN596_n_9694), .o(TIMEBOOST_net_12549) );
in01f02 g58484_u0 ( .a(FE_OFN1440_n_9372), .o(g58484_sb) );
na02s02 TIMEBOOST_cell_63368 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q), .b(g58321_sb), .o(TIMEBOOST_net_20631) );
na02f80 TIMEBOOST_cell_3709 ( .a(TIMEBOOST_net_414), .b(n_8489), .o(n_8567) );
na04f02 TIMEBOOST_cell_73504 ( .a(TIMEBOOST_net_11632), .b(TIMEBOOST_net_5472), .c(n_8757), .d(TIMEBOOST_net_6034), .o(n_14810) );
in01f02 g58485_u0 ( .a(FE_OFN1437_n_9372), .o(g58485_sb) );
na02m02 TIMEBOOST_cell_44067 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q), .o(TIMEBOOST_net_12928) );
na02f02 TIMEBOOST_cell_3711 ( .a(TIMEBOOST_net_415), .b(n_4619), .o(n_7214) );
na02s01 g57798_u1 ( .a(g57797_sb), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(g57798_da) );
in01f02 g58486_u0 ( .a(FE_OFN1440_n_9372), .o(g58486_sb) );
na04s02 TIMEBOOST_cell_73096 ( .a(TIMEBOOST_net_14486), .b(g65812_db), .c(g61863_sb), .d(g61863_db), .o(n_8111) );
na02f02 TIMEBOOST_cell_3713 ( .a(n_16444), .b(TIMEBOOST_net_416), .o(n_9154) );
in01m01 TIMEBOOST_cell_64271 ( .a(TIMEBOOST_net_21127), .o(TIMEBOOST_net_21126) );
in01s01 g58487_u0 ( .a(FE_OFN1668_n_9477), .o(g58487_sb) );
na02m04 TIMEBOOST_cell_68743 ( .a(TIMEBOOST_net_21579), .b(g64922_sb), .o(TIMEBOOST_net_9706) );
na02f02 TIMEBOOST_cell_53293 ( .a(wbu_addr_in_274), .b(n_3351), .o(TIMEBOOST_net_16864) );
na02s04 TIMEBOOST_cell_45603 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q), .o(TIMEBOOST_net_13696) );
in01s01 g58488_u0 ( .a(FE_OFN1651_n_9428), .o(g58488_sb) );
na03f02 TIMEBOOST_cell_73303 ( .a(TIMEBOOST_net_13108), .b(FE_OFN1127_g64577_p), .c(g63054_sb), .o(n_7122) );
na02m02 TIMEBOOST_cell_69083 ( .a(TIMEBOOST_net_21749), .b(g64156_sb), .o(n_4009) );
na02f04 TIMEBOOST_cell_53295 ( .a(wbu_addr_in_270), .b(n_3167), .o(TIMEBOOST_net_16865) );
in01f01 g58489_u0 ( .a(n_9144), .o(g58489_sb) );
na02f06 TIMEBOOST_cell_37113 ( .a(n_5641), .b(TIMEBOOST_net_10168), .o(TIMEBOOST_net_625) );
na02s02 TIMEBOOST_cell_68267 ( .a(TIMEBOOST_net_21341), .b(g65698_db), .o(n_2203) );
na02s01 TIMEBOOST_cell_51601 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q), .o(TIMEBOOST_net_16018) );
no02f02 g58490_u0 ( .a(n_397), .b(n_9144), .o(g58490_p) );
ao12f02 g58490_u1 ( .a(g58490_p), .b(n_397), .c(n_9144), .o(n_8917) );
no02s01 g58554_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN601_n_9687), .o(n_8971) );
no02s01 g58555_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN562_n_9895), .o(n_8970) );
no02s01 g58556_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN554_n_9864), .o(n_8968) );
no02s01 g58557_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN519_n_9697), .o(n_8967) );
no02s01 g58558_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN587_n_9692), .o(n_8966) );
no02s01 g58559_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN532_n_9823), .o(n_8965) );
no02s01 g58560_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN595_n_9694), .o(n_8964) );
no02s01 g58561_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN529_n_9899), .o(n_8963) );
no02s01 g58562_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN606_n_9904), .o(n_8962) );
no02f06 g58563_u0 ( .a(n_3024), .b(n_522), .o(n_3025) );
no02f01 g58564_u0 ( .a(n_2479), .b(FE_OFN778_n_4152), .o(n_3028) );
no02s01 g58565_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN1803_n_9690), .o(n_8961) );
no02s01 g58566_u0 ( .a(FE_OFN256_n_8969), .b(FE_OFN577_n_9902), .o(n_8960) );
na02f01 TIMEBOOST_cell_26107 ( .a(pci_target_unit_pcit_if_strd_addr_in_702), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7158) );
no02f02 g58568_u0 ( .a(n_4713), .b(FE_OFN1145_n_15261), .o(n_5754) );
na02f02 g58569_u0 ( .a(n_14967), .b(n_8493), .o(g58569_p) );
in01f02 g58569_u1 ( .a(g58569_p), .o(n_10787) );
no02f08 g58570_u0 ( .a(n_3073), .b(n_784), .o(n_3074) );
no02f02 g58571_u0 ( .a(n_2631), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8661) );
na02f04 g58572_u0 ( .a(n_1085), .b(n_9144), .o(n_9143) );
in01s01 TIMEBOOST_cell_67766 ( .a(TIMEBOOST_net_21192), .o(TIMEBOOST_net_21193) );
in01f02 g58574_u0 ( .a(FE_OFN1398_n_8567), .o(g58574_sb) );
na02m02 TIMEBOOST_cell_71971 ( .a(TIMEBOOST_net_23193), .b(g64962_sb), .o(TIMEBOOST_net_17408) );
na02s06 TIMEBOOST_cell_27113 ( .a(n_14753), .b(n_14839), .o(TIMEBOOST_net_7661) );
na02f01 TIMEBOOST_cell_26637 ( .a(FE_OFN2069_n_15978), .b(conf_wb_err_addr_in_952), .o(TIMEBOOST_net_7423) );
in01f02 g58576_u0 ( .a(FE_OFN1369_n_8567), .o(g58576_sb) );
na03f02 TIMEBOOST_cell_73571 ( .a(TIMEBOOST_net_17072), .b(FE_OFN1230_n_6391), .c(g62533_sb), .o(n_6506) );
na02s01 TIMEBOOST_cell_25312 ( .a(TIMEBOOST_net_6760), .b(n_2373), .o(TIMEBOOST_net_531) );
na02f02 g58578_u0 ( .a(n_2351), .b(n_8572), .o(n_8574) );
oa12f02 g58580_u0 ( .a(n_8680), .b(FE_OFN1437_n_9372), .c(wishbone_slave_unit_pcim_if_del_bc_in_383), .o(n_8796) );
na02m08 TIMEBOOST_cell_54013 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_132), .o(TIMEBOOST_net_17224) );
in01f02 g58582_u1 ( .a(g58582_p), .o(n_8571) );
oa12f02 g58583_u0 ( .a(n_8749), .b(n_8750), .c(n_3022), .o(n_8752) );
oa12f02 g58584_u0 ( .a(n_8749), .b(n_8750), .c(n_67), .o(n_8751) );
ao12f02 g58585_u0 ( .a(n_4715), .b(conf_wb_err_addr_in_967), .c(FE_OFN1145_n_15261), .o(n_5753) );
in01f01 g58586_u0 ( .a(FE_OFN1394_n_8567), .o(g58586_sb) );
na02m01 TIMEBOOST_cell_47579 ( .a(n_8831), .b(g58783_sb), .o(TIMEBOOST_net_14007) );
na02f02 TIMEBOOST_cell_50198 ( .a(TIMEBOOST_net_15316), .b(g60660_sb), .o(n_5660) );
na03m02 TIMEBOOST_cell_72706 ( .a(g64331_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q), .c(TIMEBOOST_net_16194), .o(TIMEBOOST_net_17325) );
in01f02 g58587_u0 ( .a(FE_OFN2185_n_8567), .o(g58587_sb) );
na02s01 TIMEBOOST_cell_48569 ( .a(FE_OFN225_n_9122), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q), .o(TIMEBOOST_net_14502) );
na03m02 TIMEBOOST_cell_67599 ( .a(TIMEBOOST_net_14649), .b(FE_OFN247_n_9112), .c(TIMEBOOST_net_14848), .o(TIMEBOOST_net_9453) );
in01f02 g58588_u0 ( .a(FE_OFN2184_n_8567), .o(g58588_sb) );
na02s02 TIMEBOOST_cell_48565 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q), .o(TIMEBOOST_net_14500) );
na03m08 TIMEBOOST_cell_72728 ( .a(TIMEBOOST_net_16913), .b(FE_OFN648_n_4497), .c(g65670_sb), .o(n_1959) );
na02s01 TIMEBOOST_cell_49430 ( .a(TIMEBOOST_net_14932), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_12978) );
in01f02 g58589_u0 ( .a(FE_OFN1403_n_8567), .o(g58589_sb) );
na02f02 TIMEBOOST_cell_69181 ( .a(TIMEBOOST_net_21798), .b(g64279_sb), .o(n_3894) );
in01s01 TIMEBOOST_cell_67762 ( .a(TIMEBOOST_net_21188), .o(TIMEBOOST_net_21189) );
in01f02 g58590_u0 ( .a(FE_OFN1403_n_8567), .o(g58590_sb) );
na02s02 TIMEBOOST_cell_48525 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q), .b(g65977_sb), .o(TIMEBOOST_net_14480) );
na03m02 TIMEBOOST_cell_66062 ( .a(n_3988), .b(g62788_sb), .c(TIMEBOOST_net_7672), .o(n_5414) );
in01f02 g58591_u0 ( .a(FE_OFN1403_n_8567), .o(g58591_sb) );
na02s02 TIMEBOOST_cell_49462 ( .a(TIMEBOOST_net_14948), .b(FE_OFN572_n_9502), .o(TIMEBOOST_net_11192) );
na02m01 TIMEBOOST_cell_27135 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_7672) );
in01f01 g58592_u0 ( .a(FE_OFN1394_n_8567), .o(g58592_sb) );
na02m08 g52475_u1 ( .a(TIMEBOOST_net_20733), .b(g52470_sb), .o(g52475_da) );
na03f02 TIMEBOOST_cell_66731 ( .a(TIMEBOOST_net_16822), .b(FE_OFN1306_n_13124), .c(g54357_sb), .o(n_13085) );
na04f10 TIMEBOOST_cell_46116 ( .a(n_2883), .b(n_1617), .c(TIMEBOOST_net_370), .d(n_15406), .o(n_13124) );
in01f02 g58593_u0 ( .a(FE_OFN1403_n_8567), .o(g58593_sb) );
in01s01 TIMEBOOST_cell_45955 ( .a(TIMEBOOST_net_13916), .o(TIMEBOOST_net_13867) );
na02f02 g53812_u0 ( .a(n_13467), .b(n_1794), .o(n_13673) );
na02f02 TIMEBOOST_cell_72263 ( .a(TIMEBOOST_net_23339), .b(g62645_sb), .o(n_6259) );
in01f01 g58594_u0 ( .a(FE_OFN1394_n_8567), .o(g58594_sb) );
na02s02 TIMEBOOST_cell_63787 ( .a(TIMEBOOST_net_20879), .b(g57999_sb), .o(TIMEBOOST_net_9469) );
na02m04 TIMEBOOST_cell_70210 ( .a(n_1953), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q), .o(TIMEBOOST_net_22313) );
na02f01 TIMEBOOST_cell_70428 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_22422) );
in01f02 g58595_u0 ( .a(FE_OFN2184_n_8567), .o(g58595_sb) );
na03s01 TIMEBOOST_cell_41743 ( .a(g58445_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q), .c(g58445_db), .o(n_9408) );
na03m02 TIMEBOOST_cell_72581 ( .a(TIMEBOOST_net_21439), .b(g64748_sb), .c(TIMEBOOST_net_21632), .o(TIMEBOOST_net_17361) );
na02m04 TIMEBOOST_cell_68936 ( .a(n_4645), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q), .o(TIMEBOOST_net_21676) );
in01f02 g58596_u0 ( .a(FE_OFN2185_n_8567), .o(g58596_sb) );
na02s02 TIMEBOOST_cell_71309 ( .a(TIMEBOOST_net_22862), .b(g58207_sb), .o(TIMEBOOST_net_20599) );
na03f02 TIMEBOOST_cell_66460 ( .a(TIMEBOOST_net_17125), .b(FE_OFN1311_n_6624), .c(g62477_sb), .o(n_6634) );
in01f02 g58597_u0 ( .a(FE_OFN1398_n_8567), .o(g58597_sb) );
na03f02 TIMEBOOST_cell_25083 ( .a(n_11823), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q), .c(n_12088), .o(n_12513) );
na03f02 TIMEBOOST_cell_66061 ( .a(n_3886), .b(g63071_sb), .c(TIMEBOOST_net_7684), .o(n_5108) );
in01f02 g58598_u0 ( .a(n_8747), .o(g58598_sb) );
na02m02 TIMEBOOST_cell_54522 ( .a(TIMEBOOST_net_17478), .b(g62489_sb), .o(n_6607) );
na03f02 TIMEBOOST_cell_66554 ( .a(g53931_sb), .b(FE_OFN1331_n_13547), .c(TIMEBOOST_net_16802), .o(n_13514) );
na04f04 TIMEBOOST_cell_24556 ( .a(n_9224), .b(g57165_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q), .d(FE_OFN1417_n_8567), .o(n_10836) );
no02f02 g58599_u0 ( .a(n_440), .b(n_14971), .o(g58599_p) );
ao12f02 g58599_u1 ( .a(g58599_p), .b(n_440), .c(n_14971), .o(n_8842) );
in01f02 g58600_u0 ( .a(n_14971), .o(g58600_sb) );
na02s01 TIMEBOOST_cell_62902 ( .a(TIMEBOOST_net_12803), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q), .o(TIMEBOOST_net_20398) );
in01f02 g58601_u0 ( .a(n_14971), .o(g58601_sb) );
na03s02 TIMEBOOST_cell_67891 ( .a(g61899_sb), .b(g61920_db), .c(n_1655), .o(n_7981) );
na02s01 TIMEBOOST_cell_48185 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_14310) );
na03f03 TIMEBOOST_cell_73683 ( .a(FE_RN_739_0), .b(n_2927), .c(n_4654), .o(n_5724) );
na03m02 TIMEBOOST_cell_71946 ( .a(FE_OFN682_n_4460), .b(g64818_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q), .o(TIMEBOOST_net_23181) );
oa12f02 g58603_u0 ( .a(n_8954), .b(FE_OFN1398_n_8567), .c(n_8953), .o(n_9340) );
oa12f02 g58604_u0 ( .a(n_8682), .b(n_8747), .c(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_8794) );
in01m02 g58605_u0 ( .a(FE_OFN1144_n_15261), .o(g58605_sb) );
na02s02 TIMEBOOST_cell_39182 ( .a(g58048_sb), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_11203) );
in01s01 TIMEBOOST_cell_73927 ( .a(TIMEBOOST_net_23491), .o(TIMEBOOST_net_23492) );
in01f02 g58606_u0 ( .a(FE_OFN2182_n_8567), .o(g58606_sb) );
na03f02 TIMEBOOST_cell_47403 ( .a(FE_OFN1588_n_13736), .b(TIMEBOOST_net_13713), .c(FE_OCP_RBN1995_n_13971), .o(n_14274) );
na02f02 TIMEBOOST_cell_38260 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(g65807_sb), .o(TIMEBOOST_net_10742) );
in01f01 g58607_u0 ( .a(FE_OFN1394_n_8567), .o(g58607_sb) );
na04f02 TIMEBOOST_cell_67191 ( .a(g64085_sb), .b(pci_target_unit_fifos_pciw_addr_data_in_124), .c(g64085_db), .d(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_20571) );
na02s01 TIMEBOOST_cell_43444 ( .a(TIMEBOOST_net_12616), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_10779) );
na03m02 TIMEBOOST_cell_72699 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q), .b(g64358_sb), .c(g64358_db), .o(n_4723) );
in01f02 g58608_u0 ( .a(FE_OFN1403_n_8567), .o(g58608_sb) );
in01s02 TIMEBOOST_cell_45920 ( .a(TIMEBOOST_net_13880), .o(TIMEBOOST_net_13881) );
in01s01 TIMEBOOST_cell_73932 ( .a(wbm_dat_i_17_), .o(TIMEBOOST_net_23497) );
in01s01 TIMEBOOST_cell_46006 ( .a(TIMEBOOST_net_13967), .o(TIMEBOOST_net_13966) );
in01f02 g58609_u0 ( .a(FE_OFN2185_n_8567), .o(g58609_sb) );
na02f01 TIMEBOOST_cell_53584 ( .a(TIMEBOOST_net_17009), .b(FE_OFN1225_n_6391), .o(TIMEBOOST_net_15519) );
in01f01 g58610_u0 ( .a(FE_OFN1394_n_8567), .o(g58610_sb) );
na02f02 TIMEBOOST_cell_38261 ( .a(TIMEBOOST_net_10742), .b(g65807_db), .o(n_1905) );
na03f02 TIMEBOOST_cell_25001 ( .a(n_10676), .b(FE_RN_471_0), .c(n_12578), .o(n_12840) );
in01m01 g58611_u0 ( .a(n_6986), .o(g58611_sb) );
na03f02 TIMEBOOST_cell_73714 ( .a(n_12010), .b(TIMEBOOST_net_13546), .c(FE_OFN1749_n_12004), .o(n_12684) );
in01f06 g58612_u0 ( .a(n_16534), .o(n_8686) );
in01f02 g58613_u0 ( .a(n_16536), .o(n_8745) );
in01f02 g58616_u0 ( .a(FE_OFN1369_n_8567), .o(g58616_sb) );
in01s01 TIMEBOOST_cell_45921 ( .a(TIMEBOOST_net_13931), .o(TIMEBOOST_net_13882) );
na02f01 TIMEBOOST_cell_71620 ( .a(TIMEBOOST_net_13596), .b(FE_OCPN1827_n_14995), .o(TIMEBOOST_net_23018) );
in01f02 g58617_u0 ( .a(FE_OFN1369_n_8567), .o(g58617_sb) );
in01s01 TIMEBOOST_cell_45922 ( .a(TIMEBOOST_net_13882), .o(TIMEBOOST_net_13883) );
na03m02 TIMEBOOST_cell_72892 ( .a(g61746_sb), .b(g61746_db), .c(n_1916), .o(n_8325) );
in01f02 g58618_u0 ( .a(FE_OFN1369_n_8567), .o(g58618_sb) );
na02f02 TIMEBOOST_cell_71271 ( .a(TIMEBOOST_net_22843), .b(g62338_sb), .o(n_6922) );
in01f02 g58619_u0 ( .a(FE_OFN1369_n_8567), .o(g58619_sb) );
na03m02 TIMEBOOST_cell_72446 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q), .b(g65875_sb), .c(g65875_db), .o(n_2059) );
na02s01 TIMEBOOST_cell_47794 ( .a(TIMEBOOST_net_14114), .b(FE_OFN529_n_9899), .o(TIMEBOOST_net_10353) );
in01f02 g58620_u0 ( .a(FE_OFN1398_n_8567), .o(g58620_sb) );
na03f02 TIMEBOOST_cell_25087 ( .a(n_11823), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q), .c(n_12072), .o(n_12494) );
na02m02 TIMEBOOST_cell_71138 ( .a(g62000_sb), .b(g62000_db), .o(TIMEBOOST_net_22777) );
in01f02 g58621_u0 ( .a(FE_OFN1398_n_8567), .o(g58621_sb) );
na03f02 TIMEBOOST_cell_25089 ( .a(n_12084), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q), .c(n_11823), .o(n_12509) );
na02f02 TIMEBOOST_cell_27159 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_7684) );
in01f02 g58622_u0 ( .a(n_8747), .o(g58622_sb) );
na04f04 TIMEBOOST_cell_24557 ( .a(n_9198), .b(g57597_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q), .d(FE_OFN1416_n_8567), .o(n_10795) );
na04f04 TIMEBOOST_cell_24646 ( .a(n_9898), .b(g57242_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q), .d(FE_OFN2173_n_8567), .o(n_11516) );
in01f04 g58624_u0 ( .a(n_15517), .o(n_8792) );
in01f08 g58628_u0 ( .a(n_15515), .o(n_8790) );
in01f02 g58630_u0 ( .a(n_8747), .o(g58630_sb) );
na03s01 TIMEBOOST_cell_52727 ( .a(g58160_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q), .c(g58160_db), .o(TIMEBOOST_net_16581) );
na02f06 TIMEBOOST_cell_4004 ( .a(n_1805), .b(FE_OFN2121_n_2687), .o(TIMEBOOST_net_562) );
in01f02 g58631_u0 ( .a(n_8747), .o(g58631_sb) );
na02f08 TIMEBOOST_cell_4005 ( .a(TIMEBOOST_net_562), .b(FE_OFN2052_n_6965), .o(TIMEBOOST_net_331) );
na02s02 TIMEBOOST_cell_52729 ( .a(FE_OFN217_n_9889), .b(g58102_sb), .o(TIMEBOOST_net_16582) );
in01f02 g58632_u0 ( .a(n_8747), .o(g58632_sb) );
na02m08 TIMEBOOST_cell_52731 ( .a(pci_target_unit_pcit_if_strd_addr_in_694), .b(n_2503), .o(TIMEBOOST_net_16583) );
na04m02 TIMEBOOST_cell_73097 ( .a(TIMEBOOST_net_20373), .b(TIMEBOOST_net_8720), .c(n_8272), .d(g61877_sb), .o(n_8076) );
in01f01 g58633_u0 ( .a(n_8747), .o(g58633_sb) );
na02s01 TIMEBOOST_cell_4010 ( .a(FE_OFN1778_parchk_pci_ad_reg_in_1222), .b(g65858_sb), .o(TIMEBOOST_net_565) );
in01f02 g58634_u0 ( .a(n_8747), .o(g58634_sb) );
na02m02 TIMEBOOST_cell_48916 ( .a(TIMEBOOST_net_14675), .b(FE_OFN579_n_9531), .o(TIMEBOOST_net_12790) );
na02f02 TIMEBOOST_cell_70233 ( .a(TIMEBOOST_net_22324), .b(FE_OFN714_n_8140), .o(TIMEBOOST_net_14916) );
na02s01 TIMEBOOST_cell_4012 ( .a(parchk_pci_ad_reg_in_1223), .b(g65858_sb), .o(TIMEBOOST_net_566) );
in01f01 g58635_u0 ( .a(n_8747), .o(g58635_sb) );
na04m02 TIMEBOOST_cell_73098 ( .a(TIMEBOOST_net_17265), .b(g65837_sb), .c(g61904_sb), .d(g61904_db), .o(n_8014) );
in01m02 g58636_u0 ( .a(FE_OFN1700_n_5751), .o(g58636_sb) );
na02f02 TIMEBOOST_cell_70893 ( .a(TIMEBOOST_net_22654), .b(g60655_sb), .o(n_5668) );
in01s01 TIMEBOOST_cell_63559 ( .a(TIMEBOOST_net_20739), .o(TIMEBOOST_net_20738) );
ao12f02 g58637_u0 ( .a(n_8732), .b(n_3158), .c(n_1077), .o(n_8734) );
ao12f02 g58638_u0 ( .a(n_8732), .b(n_3156), .c(n_1260), .o(n_8733) );
ao12f02 g58639_u0 ( .a(n_8732), .b(n_2988), .c(n_1261), .o(n_8731) );
in01f02 g58640_u0 ( .a(n_14971), .o(g58640_sb) );
na02s01 TIMEBOOST_cell_37653 ( .a(TIMEBOOST_net_10438), .b(g57962_db), .o(n_9842) );
na03f02 TIMEBOOST_cell_66762 ( .a(TIMEBOOST_net_17143), .b(FE_OFN1322_n_6436), .c(g62901_sb), .o(n_6075) );
in01f02 g58641_u0 ( .a(n_16076), .o(n_8897) );
in01f02 g58645_u0 ( .a(n_16550), .o(n_8896) );
in01f02 g58652_u0 ( .a(n_14971), .o(g58652_sb) );
na02s02 TIMEBOOST_cell_38547 ( .a(TIMEBOOST_net_10885), .b(g58203_db), .o(n_9054) );
na03f02 TIMEBOOST_cell_73445 ( .a(TIMEBOOST_net_16749), .b(FE_OFN1192_n_6935), .c(g62719_sb), .o(n_6138) );
in01f02 g58653_u0 ( .a(n_14971), .o(g58653_sb) );
na02f04 TIMEBOOST_cell_38966 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q), .b(n_13447), .o(TIMEBOOST_net_11095) );
in01s01 TIMEBOOST_cell_73883 ( .a(TIMEBOOST_net_23447), .o(TIMEBOOST_net_23448) );
na03m04 TIMEBOOST_cell_73034 ( .a(TIMEBOOST_net_21717), .b(g65007_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q), .o(TIMEBOOST_net_16774) );
in01f02 g58654_u0 ( .a(n_14971), .o(g58654_sb) );
na02m04 TIMEBOOST_cell_72010 ( .a(g65279_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q), .o(TIMEBOOST_net_23213) );
na03m02 TIMEBOOST_cell_72602 ( .a(g65371_da), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q), .c(TIMEBOOST_net_10378), .o(TIMEBOOST_net_17020) );
na02f06 TIMEBOOST_cell_47795 ( .a(n_1519), .b(n_763), .o(TIMEBOOST_net_14115) );
in01f02 g58655_u0 ( .a(n_14971), .o(g58655_sb) );
na02f02 TIMEBOOST_cell_70806 ( .a(TIMEBOOST_net_16706), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_22611) );
na03f02 TIMEBOOST_cell_69780 ( .a(FE_OFN928_n_4730), .b(pci_target_unit_fifos_pciw_addr_data_in_142), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q), .o(TIMEBOOST_net_22098) );
no03f06 TIMEBOOST_cell_21393 ( .a(FE_RN_839_0), .b(FE_RN_462_0), .c(FE_RN_837_0), .o(TIMEBOOST_net_593) );
no02f02 g58656_u0 ( .a(n_676), .b(n_7094), .o(g58656_p) );
ao12f02 g58656_u1 ( .a(g58656_p), .b(n_676), .c(n_7094), .o(n_7724) );
no02f02 g58691_u0 ( .a(n_983), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8658) );
no02f10 g58692_u0 ( .a(n_8747), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_), .o(g58692_p) );
in01f10 g58692_u1 ( .a(g58692_p), .o(n_8657) );
no02f02 g58693_u0 ( .a(n_2965), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8656) );
na02f01 g58694_u0 ( .a(n_8566), .b(n_8728), .o(n_8730) );
no02f02 g58695_u0 ( .a(n_8566), .b(n_8728), .o(g58695_p) );
in01f02 g58695_u1 ( .a(g58695_p), .o(n_8727) );
no02f02 g58696_u0 ( .a(n_2422), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8655) );
na02f04 g58697_u0 ( .a(FE_OFN1398_n_8567), .b(n_8953), .o(n_8954) );
na02f02 TIMEBOOST_cell_71142 ( .a(TIMEBOOST_net_20988), .b(g52397_sb), .o(TIMEBOOST_net_22779) );
in01s01 TIMEBOOST_cell_67759 ( .a(pci_target_unit_fifos_pcir_data_in_161), .o(TIMEBOOST_net_21186) );
na02s01 TIMEBOOST_cell_31003 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_14__Q), .b(FE_OFN213_n_9124), .o(TIMEBOOST_net_9606) );
na02f03 g58702_u0 ( .a(FE_OFN2185_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q), .o(n_8950) );
in01s04 g58706_u0 ( .a(FE_OFN256_n_8969), .o(n_8892) );
na02s02 g58708_u0 ( .a(n_8780), .b(n_8832), .o(n_8969) );
na02f02 g58709_u0 ( .a(FE_OFN2184_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q), .o(n_8949) );
na02f02 g58710_u0 ( .a(FE_OFN1402_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q), .o(n_8890) );
na02f03 g58711_u0 ( .a(FE_OFN1403_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q), .o(n_8889) );
na02f02 g58712_u0 ( .a(FE_OFN1403_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q), .o(n_8888) );
na02f02 g58713_u0 ( .a(FE_OFN1402_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q), .o(n_8947) );
na02f02 g58714_u0 ( .a(FE_OFN2184_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q), .o(n_8946) );
na02f02 g58715_u0 ( .a(FE_OFN1402_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q), .o(n_8945) );
na02f02 g58716_u0 ( .a(FE_OFN2184_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q), .o(n_8944) );
na02s02 TIMEBOOST_cell_48093 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q), .b(pci_target_unit_fifos_pcir_data_in_174), .o(TIMEBOOST_net_14264) );
na02f02 g58718_u0 ( .a(FE_OFN1402_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q), .o(n_8943) );
na02f02 g58723_u0 ( .a(FE_OFN2184_n_8567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q), .o(n_8887) );
na02f02 g58724_u0 ( .a(n_8747), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_8682) );
na02f04 g58725_u0 ( .a(n_16332), .b(FE_OFN2093_n_2301), .o(n_8572) );
na03f02 TIMEBOOST_cell_66064 ( .a(n_4029), .b(g62784_sb), .c(TIMEBOOST_net_7697), .o(n_5424) );
na02s01 TIMEBOOST_cell_39184 ( .a(FE_OFN258_n_9862), .b(g58040_sb), .o(TIMEBOOST_net_11204) );
no02f02 g58728_u0 ( .a(n_3496), .b(FE_OFN1144_n_15261), .o(n_4715) );
na02f02 TIMEBOOST_cell_18238 ( .a(TIMEBOOST_net_5482), .b(n_4661), .o(n_6985) );
no02s02 g58730_u0 ( .a(FE_OCP_DRV_N1950_n_8660), .b(wishbone_slave_unit_del_sync_comp_cycle_count_0_), .o(n_8652) );
no02f02 g58731_u0 ( .a(n_2996), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8651) );
no02f02 g58732_u0 ( .a(n_2731), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8650) );
no02f02 g58733_u0 ( .a(n_3184), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8649) );
no02f02 g58734_u0 ( .a(n_3209), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8648) );
no02f02 g58735_u0 ( .a(n_1422), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8647) );
no02f02 g58736_u0 ( .a(n_2023), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8646) );
no02s02 g58737_u0 ( .a(n_2326), .b(FE_OCP_DRV_N2262_n_8660), .o(n_8645) );
no02f02 g58738_u0 ( .a(n_1656), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8644) );
no02f02 g58739_u0 ( .a(n_2008), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8643) );
no02f02 g58740_u0 ( .a(n_2302), .b(FE_OCP_DRV_N1950_n_8660), .o(n_8642) );
no02f08 g58741_u0 ( .a(FE_OFN1344_n_8567), .b(n_8489), .o(n_9144) );
no02f08 g58742_u0 ( .a(n_1110), .b(FE_OFN1398_n_8567), .o(g58742_p) );
in01f04 g58742_u1 ( .a(g58742_p), .o(n_9341) );
na02f08 g58744_u0 ( .a(n_16577), .b(n_16573), .o(g58744_p) );
in01f08 g58744_u1 ( .a(g58744_p), .o(n_8866) );
no02f08 g58745_u0 ( .a(n_8784), .b(n_16573), .o(n_8860) );
ao12f02 g58748_u0 ( .a(n_8782), .b(n_8831), .c(wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q), .o(n_9140) );
na03f02 TIMEBOOST_cell_73572 ( .a(TIMEBOOST_net_17511), .b(FE_OFN1232_n_6391), .c(g62553_sb), .o(n_6458) );
ao12f02 g58751_u0 ( .a(n_8732), .b(n_1264), .c(n_3159), .o(n_8726) );
ao12f02 g58752_u0 ( .a(n_8732), .b(n_1259), .c(n_3076), .o(n_8725) );
ao12f02 g58753_u0 ( .a(n_8732), .b(n_1475), .c(n_2998), .o(n_8724) );
oa12f02 g58754_u0 ( .a(n_8597), .b(FE_OFN1437_n_9372), .c(wishbone_slave_unit_pcim_if_del_bc_in_382), .o(n_8723) );
na03f02 TIMEBOOST_cell_47369 ( .a(FE_OFN1583_n_12306), .b(TIMEBOOST_net_13679), .c(FE_OFN1760_n_10780), .o(n_17036) );
ao12f02 g58756_u0 ( .a(n_8732), .b(n_2223), .c(n_2958), .o(n_8721) );
ao12f02 g58757_u0 ( .a(n_5750), .b(conf_wb_err_addr_in_970), .c(FE_OFN1145_n_15261), .o(n_7341) );
ao12f02 g58758_u0 ( .a(n_3501), .b(conf_wb_err_addr_in_963), .c(FE_OFN1145_n_15261), .o(n_4714) );
no02m01 g58759_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_8_), .b(n_2179), .o(g58759_p) );
ao12f01 g58759_u1 ( .a(g58759_p), .b(pci_target_unit_del_sync_comp_cycle_count_8_), .c(n_2179), .o(n_2479) );
no02f04 g58760_u0 ( .a(conf_wb_err_addr_in_971), .b(n_3359), .o(g58760_p) );
ao12f02 g58760_u1 ( .a(g58760_p), .b(conf_wb_err_addr_in_971), .c(n_3359), .o(n_4713) );
no02m01 g58761_u0 ( .a(n_882), .b(n_2175), .o(g58761_p) );
ao12m01 g58761_u1 ( .a(g58761_p), .b(n_882), .c(n_2175), .o(n_2631) );
ao12f02 g58762_u0 ( .a(n_3502), .b(conf_wb_err_addr_in_955), .c(FE_OFN1144_n_15261), .o(n_4712) );
no02f04 g58763_u0 ( .a(wbu_addr_in_279), .b(n_3489), .o(g58763_p) );
ao12f02 g58763_u1 ( .a(g58763_p), .b(wbu_addr_in_279), .c(n_3489), .o(n_4890) );
no02f04 g58764_u0 ( .a(n_3488), .b(wbm_adr_o_30_), .o(g58764_p) );
ao12f02 g58764_u1 ( .a(g58764_p), .b(wbm_adr_o_30_), .c(n_3488), .o(n_4889) );
na02s01 TIMEBOOST_cell_18373 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_5550) );
in01m20 TIMEBOOST_cell_35516 ( .a(conf_wb_err_addr_in_955), .o(TIMEBOOST_net_10107) );
in01m01 g58767_u0 ( .a(FE_OFN2054_n_8831), .o(g58767_sb) );
na04m04 TIMEBOOST_cell_72708 ( .a(TIMEBOOST_net_12476), .b(FE_OFN2108_n_2047), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q), .d(g65683_sb), .o(TIMEBOOST_net_22322) );
na02f01 TIMEBOOST_cell_38968 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_11096) );
in01f06 g58768_u0 ( .a(n_8884), .o(g58768_sb) );
in01s01 TIMEBOOST_cell_67761 ( .a(pci_target_unit_fifos_pcir_data_in_171), .o(TIMEBOOST_net_21188) );
in01s01 g58769_u0 ( .a(n_8884), .o(g58769_sb) );
na03f02 TIMEBOOST_cell_73802 ( .a(FE_OFN1773_n_13800), .b(TIMEBOOST_net_13784), .c(FE_OFN1769_n_14054), .o(n_14500) );
na03m02 TIMEBOOST_cell_68872 ( .a(g65272_sb), .b(n_4498), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q), .o(TIMEBOOST_net_21644) );
in01m01 g58770_u0 ( .a(n_8831), .o(g58770_sb) );
na03m04 TIMEBOOST_cell_72765 ( .a(n_4645), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q), .c(TIMEBOOST_net_22006), .o(TIMEBOOST_net_13365) );
na03m02 TIMEBOOST_cell_69394 ( .a(n_4447), .b(g64945_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q), .o(TIMEBOOST_net_21905) );
na02f10 TIMEBOOST_cell_62418 ( .a(pciu_pref_en_in_320), .b(configuration_wb_err_data_571), .o(TIMEBOOST_net_20156) );
in01f10 g58771_u0 ( .a(FE_OFN2055_n_8831), .o(g58771_sb) );
na03f40 TIMEBOOST_cell_24021 ( .a(g57794_sb), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .c(g57794_db), .o(n_9173) );
no03f10 TIMEBOOST_cell_130 ( .a(FE_RN_37_0), .b(FE_RN_36_0), .c(n_16310), .o(n_16311) );
in01s01 g58772_u0 ( .a(FE_OFN2054_n_8831), .o(g58772_sb) );
na02f01 TIMEBOOST_cell_70912 ( .a(TIMEBOOST_net_16730), .b(FE_OFN1179_n_3476), .o(TIMEBOOST_net_22664) );
na02m02 TIMEBOOST_cell_38970 ( .a(g58311_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q), .o(TIMEBOOST_net_11097) );
na02f02 TIMEBOOST_cell_52926 ( .a(TIMEBOOST_net_16680), .b(g63010_sb), .o(n_5227) );
in01s01 g58773_u0 ( .a(FE_OFN2054_n_8831), .o(g58773_sb) );
na04f04 TIMEBOOST_cell_73486 ( .a(TIMEBOOST_net_17355), .b(g52402_sb), .c(g59240_sb), .d(wbm_adr_o_6_), .o(TIMEBOOST_net_22988) );
na04f02 TIMEBOOST_cell_73304 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q), .b(FE_OFN1133_g64577_p), .c(n_3880), .d(g63078_sb), .o(n_5096) );
in01f04 g58774_u0 ( .a(n_8831), .o(g58774_sb) );
na02m02 TIMEBOOST_cell_69183 ( .a(TIMEBOOST_net_21799), .b(g64268_sb), .o(n_3905) );
na02f02 TIMEBOOST_cell_70835 ( .a(TIMEBOOST_net_22625), .b(g62045_sb), .o(n_7767) );
na03m20 TIMEBOOST_cell_34 ( .a(g54038_db), .b(g54038_sb), .c(output_backup_par_out_reg_Q), .o(n_13335) );
in01s01 g58775_u0 ( .a(n_8831), .o(g58775_sb) );
na02m02 TIMEBOOST_cell_39749 ( .a(TIMEBOOST_net_11486), .b(g58339_db), .o(n_9481) );
in01f40 g58776_u0 ( .a(n_8884), .o(g58776_sb) );
na02m02 TIMEBOOST_cell_50542 ( .a(TIMEBOOST_net_15488), .b(g62954_sb), .o(n_5973) );
na04m02 TIMEBOOST_cell_67893 ( .a(g61866_sb), .b(g61866_db), .c(TIMEBOOST_net_14485), .d(g65814_db), .o(n_8105) );
in01s01 g58777_u0 ( .a(n_8884), .o(g58777_sb) );
na03f02 TIMEBOOST_cell_47325 ( .a(FE_OFN1752_n_12086), .b(TIMEBOOST_net_13615), .c(FE_OFN2209_n_11027), .o(n_12745) );
na02m01 TIMEBOOST_cell_53967 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q), .o(TIMEBOOST_net_17201) );
in01m01 g58778_u0 ( .a(n_8884), .o(g58778_sb) );
na02m04 TIMEBOOST_cell_68938 ( .a(n_4444), .b(n_156), .o(TIMEBOOST_net_21677) );
in01s01 g58779_u0 ( .a(FE_OFN2054_n_8831), .o(g58779_sb) );
na02m04 TIMEBOOST_cell_54066 ( .a(TIMEBOOST_net_17250), .b(FE_OFN1049_n_16657), .o(TIMEBOOST_net_14722) );
na04m06 TIMEBOOST_cell_72835 ( .a(n_3741), .b(g64866_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q), .d(g64866_db), .o(TIMEBOOST_net_17550) );
na02f02 TIMEBOOST_cell_54286 ( .a(TIMEBOOST_net_17360), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_15325) );
na03f02 TIMEBOOST_cell_70014 ( .a(n_1607), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q), .c(FE_OFN716_n_8176), .o(TIMEBOOST_net_22215) );
in01s01 TIMEBOOST_cell_67772 ( .a(TIMEBOOST_net_21198), .o(TIMEBOOST_net_21199) );
na03m02 TIMEBOOST_cell_70158 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q), .b(FE_OFN1076_n_4740), .c(pci_target_unit_fifos_pciw_addr_data_in_146), .o(TIMEBOOST_net_22287) );
in01m01 g58782_u0 ( .a(n_8884), .o(g58782_sb) );
na04m02 TIMEBOOST_cell_65193 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q), .b(n_8272), .c(g61994_sb), .d(n_2165), .o(n_7907) );
na04m02 TIMEBOOST_cell_73099 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q), .b(g65816_sb), .c(TIMEBOOST_net_13438), .d(g65816_db), .o(TIMEBOOST_net_9803) );
na02m01 TIMEBOOST_cell_29343 ( .a(n_3780), .b(FE_OFN1676_n_4655), .o(TIMEBOOST_net_8776) );
in01m01 g58783_u0 ( .a(n_8831), .o(g58783_sb) );
na02s02 TIMEBOOST_cell_39761 ( .a(TIMEBOOST_net_11492), .b(g57941_db), .o(n_9129) );
na02s01 TIMEBOOST_cell_37605 ( .a(TIMEBOOST_net_10414), .b(g58146_db), .o(n_9648) );
na03f02 TIMEBOOST_cell_66040 ( .a(n_4073), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q), .c(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_11386) );
na02f01 TIMEBOOST_cell_44560 ( .a(TIMEBOOST_net_13174), .b(g63557_sb), .o(n_4920) );
na02s01 TIMEBOOST_cell_18113 ( .a(pci_target_unit_del_sync_be_out_reg_1__Q), .b(FE_OFN786_n_2678), .o(TIMEBOOST_net_5420) );
in01s01 g58785_u0 ( .a(FE_OFN2055_n_8831), .o(g58785_sb) );
na02m02 TIMEBOOST_cell_62678 ( .a(g65739_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q), .o(TIMEBOOST_net_20286) );
na03f02 TIMEBOOST_cell_46797 ( .a(TIMEBOOST_net_8788), .b(FE_OFN1165_n_5615), .c(g62089_sb), .o(n_5618) );
na02s01 TIMEBOOST_cell_31005 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_27__Q), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_9607) );
in01s01 g58786_u0 ( .a(FE_OFN2055_n_8831), .o(g58786_sb) );
na02f01 TIMEBOOST_cell_20253 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_6490) );
in01s01 g58787_u0 ( .a(n_8884), .o(g58787_sb) );
na04f04 TIMEBOOST_cell_36617 ( .a(n_2328), .b(FE_OFN1330_n_13547), .c(g59763_sb), .d(n_16763), .o(n_7625) );
na02m02 g58406_u2 ( .a(FE_OFN247_n_9112), .b(FE_OFN1632_n_9531), .o(g58406_db) );
na02m10 TIMEBOOST_cell_45439 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_13614) );
in01f10 g58788_u0 ( .a(FE_OFN2054_n_8831), .o(g58788_sb) );
na02s06 TIMEBOOST_cell_63808 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q), .o(TIMEBOOST_net_20890) );
in01s01 TIMEBOOST_cell_73976 ( .a(wbm_dat_i_8_), .o(TIMEBOOST_net_23541) );
in01s01 TIMEBOOST_cell_67790 ( .a(TIMEBOOST_net_21217), .o(TIMEBOOST_net_21216) );
in01f04 g58789_u0 ( .a(n_8831), .o(g58789_sb) );
na03f02 TIMEBOOST_cell_65337 ( .a(TIMEBOOST_net_16310), .b(n_5633), .c(g62132_sb), .o(n_5563) );
in01f40 g58790_u0 ( .a(FE_OFN2055_n_8831), .o(g58790_sb) );
na02m10 TIMEBOOST_cell_45389 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_13589) );
na02f02 TIMEBOOST_cell_49942 ( .a(TIMEBOOST_net_15188), .b(g63069_sb), .o(n_5112) );
in01m01 g58791_u0 ( .a(FE_OFN2054_n_8831), .o(g58791_sb) );
na03f02 TIMEBOOST_cell_66351 ( .a(TIMEBOOST_net_17145), .b(FE_OFN1234_n_6391), .c(g62936_sb), .o(n_6009) );
in01s01 g58792_u0 ( .a(n_8884), .o(g58792_sb) );
na02f02 TIMEBOOST_cell_50536 ( .a(TIMEBOOST_net_15485), .b(g63168_sb), .o(n_5802) );
na02f02 TIMEBOOST_cell_44990 ( .a(TIMEBOOST_net_13389), .b(g54203_db), .o(g53942_db) );
na02s01 TIMEBOOST_cell_47641 ( .a(g61962_sb), .b(wbs_dat_i_14_), .o(TIMEBOOST_net_14038) );
in01s01 g58793_u0 ( .a(n_8831), .o(g58793_sb) );
na02m10 TIMEBOOST_cell_69574 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_135), .o(TIMEBOOST_net_21995) );
in01s01 TIMEBOOST_cell_73884 ( .a(n_8323), .o(TIMEBOOST_net_23449) );
na02s02 TIMEBOOST_cell_45005 ( .a(g58394_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q), .o(TIMEBOOST_net_13397) );
in01s01 g58794_u0 ( .a(n_8831), .o(g58794_sb) );
na02m10 TIMEBOOST_cell_52999 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q), .b(wishbone_slave_unit_pcim_sm_data_in_645), .o(TIMEBOOST_net_16717) );
in01s01 g58795_u0 ( .a(FE_OFN2055_n_8831), .o(g58795_sb) );
in01s01 TIMEBOOST_cell_31900 ( .a(TIMEBOOST_net_10064), .o(TIMEBOOST_net_10063) );
na03m02 TIMEBOOST_cell_73100 ( .a(TIMEBOOST_net_10660), .b(g65818_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q), .o(TIMEBOOST_net_22195) );
na02m02 TIMEBOOST_cell_49738 ( .a(TIMEBOOST_net_15086), .b(TIMEBOOST_net_11193), .o(TIMEBOOST_net_9434) );
na02m01 TIMEBOOST_cell_18107 ( .a(pci_target_unit_pcit_if_strd_addr_in_716), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_5417) );
na02f02 TIMEBOOST_cell_70837 ( .a(TIMEBOOST_net_22626), .b(g62039_sb), .o(n_7776) );
in01s01 g58797_u0 ( .a(FE_OFN2054_n_8831), .o(g58797_sb) );
na02f01 TIMEBOOST_cell_48123 ( .a(pciu_pciif_stop_reg_in), .b(g65994_sb), .o(TIMEBOOST_net_14279) );
na03f02 TIMEBOOST_cell_73101 ( .a(TIMEBOOST_net_22051), .b(g65387_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q), .o(TIMEBOOST_net_16772) );
in01s01 g58798_u0 ( .a(FE_OFN2055_n_8831), .o(g58798_sb) );
na04m04 TIMEBOOST_cell_72547 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(g65737_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q), .d(g65737_db), .o(TIMEBOOST_net_22041) );
na02s02 g58798_u2 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q), .b(n_8831), .o(g58798_db) );
in01m02 g58799_u0 ( .a(FE_OFN1700_n_5751), .o(g58799_sb) );
na02s02 TIMEBOOST_cell_52420 ( .a(TIMEBOOST_net_16427), .b(g58005_sb), .o(TIMEBOOST_net_9521) );
in01m02 g58800_u0 ( .a(FE_OFN1697_n_5751), .o(g58800_sb) );
na03m04 TIMEBOOST_cell_72504 ( .a(TIMEBOOST_net_21356), .b(n_3780), .c(TIMEBOOST_net_21466), .o(TIMEBOOST_net_17056) );
in01f02 g58801_u0 ( .a(FE_OFN2153_n_16439), .o(g58801_sb) );
na02s02 TIMEBOOST_cell_53996 ( .a(TIMEBOOST_net_17215), .b(FE_OFN951_n_2055), .o(TIMEBOOST_net_14334) );
na02f01 TIMEBOOST_cell_70900 ( .a(TIMEBOOST_net_17357), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_22658) );
in01f02 g58802_u0 ( .a(FE_OFN2153_n_16439), .o(g58802_sb) );
na02s02 TIMEBOOST_cell_52406 ( .a(TIMEBOOST_net_16420), .b(g58132_db), .o(n_9073) );
in01f02 g58803_u0 ( .a(FE_OFN2157_n_16439), .o(g58803_sb) );
na02f02 TIMEBOOST_cell_70901 ( .a(TIMEBOOST_net_22658), .b(g60639_sb), .o(n_5691) );
na02m02 TIMEBOOST_cell_71935 ( .a(TIMEBOOST_net_23175), .b(n_4470), .o(TIMEBOOST_net_16293) );
in01f02 g58804_u0 ( .a(FE_OFN2157_n_16439), .o(g58804_sb) );
na03f02 TIMEBOOST_cell_24729 ( .a(TIMEBOOST_net_674), .b(g59798_db), .c(g52405_db), .o(n_14814) );
na03f02 TIMEBOOST_cell_70742 ( .a(TIMEBOOST_net_5685), .b(n_3486), .c(FE_OFN1700_n_5751), .o(TIMEBOOST_net_22579) );
na04f02 TIMEBOOST_cell_67193 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(g64105_sb), .c(TIMEBOOST_net_10434), .d(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q), .o(TIMEBOOST_net_20460) );
in01f02 g58805_u0 ( .a(FE_OFN2153_n_16439), .o(g58805_sb) );
na02m01 TIMEBOOST_cell_48707 ( .a(TIMEBOOST_net_12475), .b(FE_OFN2109_n_2047), .o(TIMEBOOST_net_14571) );
in01f02 g58806_u0 ( .a(FE_OFN2153_n_16439), .o(g58806_sb) );
na03f01 TIMEBOOST_cell_69132 ( .a(TIMEBOOST_net_14058), .b(n_5769), .c(n_16271), .o(TIMEBOOST_net_21774) );
na03f02 TIMEBOOST_cell_73456 ( .a(TIMEBOOST_net_20523), .b(FE_OFN1264_n_4095), .c(g62944_sb), .o(n_5993) );
in01f02 g58807_u0 ( .a(FE_OFN2153_n_16439), .o(g58807_sb) );
na02s01 TIMEBOOST_cell_70269 ( .a(TIMEBOOST_net_22342), .b(g58019_db), .o(TIMEBOOST_net_14973) );
na04f04 TIMEBOOST_cell_73305 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q), .b(FE_OFN1121_g64577_p), .c(n_3923), .d(g63033_sb), .o(n_5181) );
in01f02 g58808_u0 ( .a(FE_OFN2153_n_16439), .o(g58808_sb) );
na03s02 TIMEBOOST_cell_35793 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q), .b(g58391_sb), .c(g58391_db), .o(n_9441) );
na03s02 TIMEBOOST_cell_35847 ( .a(n_2066), .b(g61702_sb), .c(g61702_db), .o(n_8423) );
na04f04 TIMEBOOST_cell_73657 ( .a(TIMEBOOST_net_15874), .b(n_7508), .c(TIMEBOOST_net_403), .d(n_13922), .o(n_14619) );
in01f02 g58809_u0 ( .a(FE_OFN2158_n_16439), .o(g58809_sb) );
na03m02 TIMEBOOST_cell_72982 ( .a(TIMEBOOST_net_16611), .b(FE_OFN1056_n_4727), .c(g64229_sb), .o(TIMEBOOST_net_8799) );
na02f20 TIMEBOOST_cell_47542 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q), .b(TIMEBOOST_net_13988), .o(TIMEBOOST_net_12254) );
in01f02 g58810_u0 ( .a(FE_OFN2153_n_16439), .o(g58810_sb) );
na02s01 TIMEBOOST_cell_62474 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_86), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_20184) );
in01f02 g58811_u0 ( .a(FE_OFN2158_n_16439), .o(g58811_sb) );
na03f02 TIMEBOOST_cell_73747 ( .a(TIMEBOOST_net_16511), .b(FE_OFN1755_n_12681), .c(FE_OCP_RBN1973_n_12381), .o(n_15935) );
na03f02 TIMEBOOST_cell_66940 ( .a(FE_OFN1752_n_12086), .b(TIMEBOOST_net_16506), .c(FE_OFN2210_n_11027), .o(n_12618) );
in01f02 g58812_u0 ( .a(FE_OFN2153_n_16439), .o(g58812_sb) );
in01s01 TIMEBOOST_cell_63595 ( .a(TIMEBOOST_net_20775), .o(TIMEBOOST_net_20774) );
na02s01 TIMEBOOST_cell_47631 ( .a(g61962_sb), .b(wbs_dat_i_15_), .o(TIMEBOOST_net_14033) );
na02s01 TIMEBOOST_cell_38470 ( .a(g58237_sb), .b(FE_OFN221_n_9846), .o(TIMEBOOST_net_10847) );
in01f02 g58813_u0 ( .a(FE_OFN2153_n_16439), .o(g58813_sb) );
na02m02 TIMEBOOST_cell_68673 ( .a(TIMEBOOST_net_21544), .b(TIMEBOOST_net_10494), .o(TIMEBOOST_net_17049) );
na02m02 TIMEBOOST_cell_68745 ( .a(TIMEBOOST_net_21580), .b(TIMEBOOST_net_14207), .o(TIMEBOOST_net_17502) );
na03m02 TIMEBOOST_cell_69798 ( .a(n_3761), .b(FE_OFN643_n_4677), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q), .o(TIMEBOOST_net_22107) );
in01f02 g58814_u0 ( .a(FE_OFN2157_n_16439), .o(g58814_sb) );
na03m02 TIMEBOOST_cell_64563 ( .a(FE_OFN669_n_4505), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q), .c(n_3783), .o(TIMEBOOST_net_10333) );
na02s01 TIMEBOOST_cell_38471 ( .a(TIMEBOOST_net_10847), .b(g58241_db), .o(n_9550) );
na03f02 TIMEBOOST_cell_73030 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(FE_OFN1035_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q), .o(TIMEBOOST_net_22194) );
in01f02 g58815_u0 ( .a(FE_OFN2153_n_16439), .o(g58815_sb) );
na02f08 TIMEBOOST_cell_71392 ( .a(TIMEBOOST_net_11793), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_22904) );
in01f02 g58816_u0 ( .a(FE_OFN2158_n_16439), .o(g58816_sb) );
na02m10 TIMEBOOST_cell_45469 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q), .o(TIMEBOOST_net_13629) );
na02s01 TIMEBOOST_cell_47629 ( .a(g61962_sb), .b(wbs_dat_i_0_), .o(TIMEBOOST_net_14032) );
in01f02 g58817_u0 ( .a(FE_OFN2156_n_16439), .o(g58817_sb) );
na02f01 TIMEBOOST_cell_26476 ( .a(TIMEBOOST_net_7342), .b(g63085_sb), .o(n_5084) );
in01f02 g58818_u0 ( .a(FE_OFN2157_n_16439), .o(g58818_sb) );
na03m02 TIMEBOOST_cell_65863 ( .a(TIMEBOOST_net_17297), .b(FE_OFN719_n_8060), .c(g61762_sb), .o(n_8288) );
na02f20 TIMEBOOST_cell_47545 ( .a(conf_wb_err_bc_in_846), .b(conf_wb_err_bc_in), .o(TIMEBOOST_net_13990) );
in01f02 g58819_u0 ( .a(FE_OFN2158_n_16439), .o(g58819_sb) );
na03f02 TIMEBOOST_cell_70636 ( .a(n_4043), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q), .c(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_22526) );
in01s01 TIMEBOOST_cell_64270 ( .a(TIMEBOOST_net_21126), .o(pci_target_unit_fifos_pcir_data_in_170) );
in01f02 g58820_u0 ( .a(FE_OFN2153_n_16439), .o(g58820_sb) );
na03f02 TIMEBOOST_cell_73573 ( .a(TIMEBOOST_net_20579), .b(FE_OFN1235_n_6391), .c(g62406_sb), .o(n_6788) );
na03f02 TIMEBOOST_cell_73748 ( .a(TIMEBOOST_net_13589), .b(FE_OCP_RBN1980_n_10273), .c(FE_OFN1553_n_12104), .o(n_12715) );
in01f02 g58821_u0 ( .a(FE_OFN2153_n_16439), .o(g58821_sb) );
na03f02 TIMEBOOST_cell_24751 ( .a(TIMEBOOST_net_5560), .b(n_10155), .c(n_10792), .o(n_10793) );
in01s01 TIMEBOOST_cell_64269 ( .a(TIMEBOOST_net_21124), .o(TIMEBOOST_net_21125) );
in01f02 g58822_u0 ( .a(FE_OFN2153_n_16439), .o(g58822_sb) );
na03m02 TIMEBOOST_cell_72967 ( .a(wbu_latency_tim_val_in_249), .b(g58611_sb), .c(g59092_sb), .o(TIMEBOOST_net_20910) );
na02m04 TIMEBOOST_cell_25713 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q), .b(FE_OFN905_n_4736), .o(TIMEBOOST_net_6961) );
na02m10 TIMEBOOST_cell_54075 ( .a(pci_target_unit_pcit_if_strd_addr_in_707), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71), .o(TIMEBOOST_net_17255) );
in01f02 g58823_u0 ( .a(FE_OFN2156_n_16439), .o(g58823_sb) );
na03f02 TIMEBOOST_cell_73610 ( .a(n_4735), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_22896) );
na03f02 TIMEBOOST_cell_73457 ( .a(TIMEBOOST_net_20530), .b(FE_OFN1269_n_4095), .c(g62349_sb), .o(n_6902) );
in01f02 g58824_u0 ( .a(FE_OFN2158_n_16439), .o(g58824_sb) );
na03m02 TIMEBOOST_cell_72872 ( .a(TIMEBOOST_net_21697), .b(g64132_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q), .o(TIMEBOOST_net_13093) );
in01s01 TIMEBOOST_cell_67794 ( .a(TIMEBOOST_net_21220), .o(TIMEBOOST_net_21221) );
in01f02 g58825_u0 ( .a(FE_OFN2153_n_16439), .o(g58825_sb) );
na03f02 TIMEBOOST_cell_66556 ( .a(g53915_sb), .b(FE_OFN1331_n_13547), .c(TIMEBOOST_net_16797), .o(n_13527) );
in01f02 g58826_u0 ( .a(FE_OFN2155_n_16439), .o(g58826_sb) );
na02s01 TIMEBOOST_cell_48177 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q), .o(TIMEBOOST_net_14306) );
na03f01 TIMEBOOST_cell_69686 ( .a(FE_OFN1677_n_4655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q), .c(n_4447), .o(TIMEBOOST_net_22051) );
in01f02 g58827_u0 ( .a(FE_OFN2155_n_16439), .o(g58827_sb) );
na04f04 TIMEBOOST_cell_24671 ( .a(n_9034), .b(g57413_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q), .d(FE_OFN2169_n_8567), .o(n_10363) );
na03m02 TIMEBOOST_cell_72595 ( .a(n_3744), .b(FE_OFN654_n_4508), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q), .o(TIMEBOOST_net_22016) );
in01f02 g58828_u0 ( .a(FE_OFN2155_n_16439), .o(g58828_sb) );
na04f04 TIMEBOOST_cell_24673 ( .a(n_9219), .b(g57405_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q), .d(FE_OFN2182_n_8567), .o(n_10829) );
na02f01 TIMEBOOST_cell_71976 ( .a(n_3785), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q), .o(TIMEBOOST_net_23196) );
in01f02 g58829_u0 ( .a(FE_OFN2155_n_16439), .o(g58829_sb) );
na04f04 TIMEBOOST_cell_24675 ( .a(n_9548), .b(g57387_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q), .d(FE_OFN2191_n_8567), .o(n_11357) );
na02s01 TIMEBOOST_cell_45309 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q), .o(TIMEBOOST_net_13549) );
in01f02 g58830_u0 ( .a(FE_OFN2157_n_16439), .o(g58830_sb) );
na03m04 TIMEBOOST_cell_73102 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q), .c(TIMEBOOST_net_16339), .o(TIMEBOOST_net_17514) );
na03m10 TIMEBOOST_cell_64560 ( .a(FE_OFN225_n_9122), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q), .c(FE_OFN527_n_9899), .o(TIMEBOOST_net_10616) );
in01f02 g58831_u0 ( .a(FE_OFN2156_n_16439), .o(g58831_sb) );
in01f06 TIMEBOOST_cell_64268 ( .a(pci_target_unit_fifos_pcir_data_in_160), .o(TIMEBOOST_net_21124) );
na03f02 TIMEBOOST_cell_73306 ( .a(TIMEBOOST_net_17318), .b(FE_OFN1129_g64577_p), .c(g63036_sb), .o(n_5176) );
na03f02 TIMEBOOST_cell_65664 ( .a(TIMEBOOST_net_16357), .b(g64223_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q), .o(TIMEBOOST_net_17324) );
in01f02 g58832_u0 ( .a(FE_OFN2155_n_16439), .o(g58832_sb) );
na04f04 TIMEBOOST_cell_24677 ( .a(n_9046), .b(g57377_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q), .d(FE_OFN2169_n_8567), .o(n_10378) );
na03f02 TIMEBOOST_cell_66952 ( .a(FE_OFN1752_n_12086), .b(TIMEBOOST_net_16508), .c(FE_OFN2209_n_11027), .o(n_12751) );
na02m06 TIMEBOOST_cell_26357 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q), .b(n_13447), .o(TIMEBOOST_net_7283) );
in01f02 g58833_u0 ( .a(FE_OFN2156_n_16439), .o(g58833_sb) );
na02m10 TIMEBOOST_cell_45621 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q), .o(TIMEBOOST_net_13705) );
na03m02 TIMEBOOST_cell_69084 ( .a(FE_OFN1012_n_4734), .b(pci_target_unit_fifos_pciw_control_in_157), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q), .o(TIMEBOOST_net_21750) );
in01f02 g58834_u0 ( .a(FE_OFN2156_n_16439), .o(g58834_sb) );
na02m01 TIMEBOOST_cell_62814 ( .a(n_3755), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q), .o(TIMEBOOST_net_20354) );
na03m06 TIMEBOOST_cell_72661 ( .a(TIMEBOOST_net_23158), .b(FE_OFN927_n_4730), .c(g64286_sb), .o(n_3887) );
na02m01 TIMEBOOST_cell_26361 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_), .b(n_6986), .o(TIMEBOOST_net_7285) );
in01f02 g58835_u0 ( .a(FE_OFN2153_n_16439), .o(g58835_sb) );
na02m02 TIMEBOOST_cell_52392 ( .a(TIMEBOOST_net_16413), .b(g61744_sb), .o(n_8329) );
na02s01 TIMEBOOST_cell_53041 ( .a(configuration_pci_err_data_529), .b(wbm_dat_o_28_), .o(TIMEBOOST_net_16738) );
in01f02 g58836_u0 ( .a(FE_OFN2157_n_16439), .o(g58836_sb) );
na04f06 TIMEBOOST_cell_24685 ( .a(n_3062), .b(n_2913), .c(FE_OFN2260_n_2775), .d(n_2836), .o(n_4170) );
na02m01 TIMEBOOST_cell_26362 ( .a(TIMEBOOST_net_7285), .b(n_4662), .o(TIMEBOOST_net_668) );
in01f02 g58837_u0 ( .a(FE_OFN1437_n_9372), .o(g58837_sb) );
na03f04 TIMEBOOST_cell_46304 ( .a(g64354_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q), .c(TIMEBOOST_net_8231), .o(TIMEBOOST_net_9127) );
na02f02 TIMEBOOST_cell_71775 ( .a(TIMEBOOST_net_23095), .b(FE_OFN1771_n_14054), .o(n_14449) );
in01f02 g58838_u0 ( .a(FE_OFN1438_n_9372), .o(g58838_sb) );
na02m02 TIMEBOOST_cell_44844 ( .a(TIMEBOOST_net_13316), .b(g60663_sb), .o(n_5656) );
na02f03 TIMEBOOST_cell_3717 ( .a(TIMEBOOST_net_418), .b(n_9173), .o(n_8877) );
na03m06 TIMEBOOST_cell_64950 ( .a(TIMEBOOST_net_20271), .b(FE_OFN2108_n_2047), .c(g65773_sb), .o(n_1912) );
in01f02 g58839_u0 ( .a(FE_OFN1438_n_9372), .o(g58839_sb) );
na03m01 TIMEBOOST_cell_72568 ( .a(pci_target_unit_del_sync_addr_in_220), .b(g66402_sb), .c(g66404_db), .o(n_2536) );
in01f02 g58840_u0 ( .a(FE_OFN1438_n_9372), .o(g58840_sb) );
na02f02 TIMEBOOST_cell_70555 ( .a(TIMEBOOST_net_22485), .b(g63018_sb), .o(n_5212) );
na02s02 TIMEBOOST_cell_3721 ( .a(TIMEBOOST_net_420), .b(n_15515), .o(n_8852) );
na03f02 TIMEBOOST_cell_35105 ( .a(TIMEBOOST_net_10026), .b(FE_OFN2155_n_16439), .c(g58828_sb), .o(n_8611) );
in01f02 g58841_u0 ( .a(FE_OFN1438_n_9372), .o(g58841_sb) );
na03s01 TIMEBOOST_cell_41933 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q), .b(g58374_sb), .c(g58374_db), .o(n_9455) );
na02f08 TIMEBOOST_cell_3723 ( .a(TIMEBOOST_net_421), .b(n_16161), .o(n_16167) );
na02s01 TIMEBOOST_cell_49739 ( .a(g58426_sb), .b(n_15567), .o(TIMEBOOST_net_15087) );
in01f02 g58842_u0 ( .a(FE_OFN21_n_9372), .o(g58842_sb) );
na03f06 TIMEBOOST_cell_21392 ( .a(n_16156), .b(pci_target_unit_wishbone_master_burst_chopped), .c(n_15388), .o(n_15389) );
na03f02 TIMEBOOST_cell_34800 ( .a(TIMEBOOST_net_9550), .b(FE_OFN1390_n_8567), .c(g57286_sb), .o(n_11467) );
na02m04 TIMEBOOST_cell_42849 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_149), .o(TIMEBOOST_net_12319) );
in01f01 g58843_u0 ( .a(FE_OFN1700_n_5751), .o(g58843_sb) );
na04f02 TIMEBOOST_cell_67527 ( .a(n_4741), .b(g62821_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q), .d(FE_OFN1097_g64577_p), .o(n_7130) );
na02s01 TIMEBOOST_cell_3997 ( .a(TIMEBOOST_net_558), .b(n_4177), .o(n_4711) );
in01s02 g58855_u0 ( .a(pci_target_unit_wishbone_master_reset_rty_cnt), .o(n_8732) );
no02f02 g58859_u0 ( .a(FE_OFN1437_n_9372), .b(wishbone_slave_unit_pcim_if_del_bc_in), .o(n_8598) );
in01f02 g58860_u0 ( .a(n_8596), .o(n_8597) );
no02f02 g58861_u0 ( .a(n_8569), .b(TIMEBOOST_net_20753), .o(n_8596) );
in01s02 g58863_u0 ( .a(n_8782), .o(n_8832) );
no02s02 g58865_u0 ( .a(n_8831), .b(n_1323), .o(n_8782) );
no02s01 g58866_u0 ( .a(n_8665), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__Q), .o(n_8780) );
no02f04 g58871_u0 ( .a(n_3206), .b(FE_OFN1144_n_15261), .o(n_3502) );
no02f02 g58872_u0 ( .a(n_3210), .b(FE_OFN1144_n_15261), .o(n_3501) );
no02f02 g58873_u0 ( .a(n_4707), .b(FE_OFN1145_n_15261), .o(n_5750) );
na02m01 TIMEBOOST_cell_71830 ( .a(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q), .o(TIMEBOOST_net_23123) );
no02f01 g58875_u0 ( .a(n_665), .b(n_8569), .o(n_8568) );
na03f02 TIMEBOOST_cell_73307 ( .a(TIMEBOOST_net_8799), .b(FE_OFN2105_g64577_p), .c(g63014_sb), .o(n_5221) );
na02f02 g58_u0 ( .a(n_15527), .b(n_15539), .o(n_15540) );
no02s01 g59072_u0 ( .a(n_3211), .b(FE_OFN778_n_4152), .o(n_3497) );
na03f02 TIMEBOOST_cell_67090 ( .a(FE_OFN1593_n_13741), .b(n_13873), .c(TIMEBOOST_net_13798), .o(n_14403) );
in01f02 g59074_u0 ( .a(n_16332), .o(n_8538) );
oa12f02 g59081_u0 ( .a(n_8668), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .c(n_8590), .o(n_8669) );
in01f01 g59082_u0 ( .a(n_8590), .o(g59082_sb) );
na02s02 TIMEBOOST_cell_28171 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q), .b(g65860_sb), .o(TIMEBOOST_net_8190) );
na04f04 TIMEBOOST_cell_24619 ( .a(n_9452), .b(g57518_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q), .d(FE_OFN2188_n_8567), .o(n_11222) );
ao12f02 g59083_u0 ( .a(n_7720), .b(wishbone_slave_unit_del_sync_comp_done_reg_clr), .c(TIMEBOOST_net_20761), .o(n_8496) );
ao12f02 g59084_u0 ( .a(n_2877), .b(n_7704), .c(n_709), .o(n_8495) );
no02f04 g59086_u0 ( .a(conf_wb_err_addr_in_967), .b(n_3008), .o(g59086_p) );
ao12f02 g59086_u1 ( .a(g59086_p), .b(conf_wb_err_addr_in_967), .c(n_3008), .o(n_3496) );
oa12f02 g59087_u0 ( .a(n_3492), .b(n_3491), .c(wbu_addr_in_275), .o(n_4708) );
oa12f02 g59088_u0 ( .a(n_8492), .b(n_16876), .c(n_8564), .o(n_8565) );
in01f02 g59089_u0 ( .a(n_8590), .o(g59089_sb) );
na02m01 TIMEBOOST_cell_37180 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q), .o(TIMEBOOST_net_10202) );
na03f01 TIMEBOOST_cell_73308 ( .a(TIMEBOOST_net_17323), .b(FE_OFN1116_g64577_p), .c(g62823_sb), .o(n_5332) );
in01f04 g59090_u0 ( .a(FE_OCPN1847_n_14981), .o(g59090_sb) );
na03f02 TIMEBOOST_cell_34843 ( .a(TIMEBOOST_net_9462), .b(FE_OFN1411_n_8567), .c(g57080_sb), .o(n_11662) );
na03m02 TIMEBOOST_cell_69814 ( .a(TIMEBOOST_net_14460), .b(g64920_sb), .c(n_4394), .o(TIMEBOOST_net_22115) );
na03f02 TIMEBOOST_cell_67992 ( .a(TIMEBOOST_net_13236), .b(FE_OFN1244_n_4092), .c(g62422_sb), .o(n_6752) );
in01m01 g59092_u0 ( .a(n_4662), .o(g59092_sb) );
in01s01 TIMEBOOST_cell_45923 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_), .o(TIMEBOOST_net_13884) );
na02f06 TIMEBOOST_cell_3647 ( .a(TIMEBOOST_net_383), .b(n_7108), .o(n_8514) );
in01f01 g59093_u0 ( .a(FE_OFN1705_n_4868), .o(g59093_sb) );
na02f08 TIMEBOOST_cell_3725 ( .a(TIMEBOOST_net_422), .b(n_16459), .o(n_17031) );
na02s04 TIMEBOOST_cell_68110 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_100), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_21263) );
na02m06 TIMEBOOST_cell_54077 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q), .b(pci_target_unit_fifos_pciw_cbe_in_153), .o(TIMEBOOST_net_17256) );
oa12s02 g59094_u0 ( .a(n_8664), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .c(FE_OCPN1847_n_14981), .o(n_8765) );
no02f01 g59095_u0 ( .a(n_425), .b(n_8590), .o(g59095_p) );
ao12f01 g59095_u1 ( .a(g59095_p), .b(n_425), .c(n_8590), .o(n_8588) );
in01f01 g59096_u0 ( .a(FE_OFN1698_n_5751), .o(g59096_sb) );
na02f01 TIMEBOOST_cell_39534 ( .a(TIMEBOOST_net_9128), .b(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_11379) );
na02f10 TIMEBOOST_cell_48659 ( .a(n_16021), .b(n_15055), .o(TIMEBOOST_net_14547) );
in01m01 g59097_u0 ( .a(n_14389), .o(g59097_sb) );
na03f02 TIMEBOOST_cell_66236 ( .a(TIMEBOOST_net_20597), .b(FE_OFN1250_n_4093), .c(g62707_sb), .o(n_6152) );
na02f02 TIMEBOOST_cell_50964 ( .a(TIMEBOOST_net_15699), .b(g62608_sb), .o(n_6337) );
in01f04 g59098_u0 ( .a(FE_OCPN1847_n_14981), .o(g59098_sb) );
na03f02 TIMEBOOST_cell_34845 ( .a(TIMEBOOST_net_9470), .b(FE_OFN1381_n_8567), .c(g57142_sb), .o(n_10465) );
na02m02 TIMEBOOST_cell_53851 ( .a(n_4283), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q), .o(TIMEBOOST_net_17143) );
in01f06 g59099_u0 ( .a(n_16577), .o(n_8784) );
in01f02 g59102_u0 ( .a(n_16537), .o(n_8712) );
in01f02 g59105_u0 ( .a(n_16573), .o(n_8711) );
in01f01 g59109_u0 ( .a(FE_OCPN1847_n_14981), .o(g59109_sb) );
na02s01 TIMEBOOST_cell_49740 ( .a(TIMEBOOST_net_15087), .b(TIMEBOOST_net_11189), .o(TIMEBOOST_net_9342) );
na04f04 TIMEBOOST_cell_73309 ( .a(n_3876), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q), .c(FE_OFN1119_g64577_p), .d(g63080_sb), .o(n_5092) );
in01f04 g59110_u0 ( .a(FE_OCPN1847_n_14981), .o(g59110_sb) );
in01s01 TIMEBOOST_cell_63571 ( .a(TIMEBOOST_net_20751), .o(TIMEBOOST_net_20750) );
na03f02 TIMEBOOST_cell_66291 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q), .b(g63199_sb), .c(g63199_db), .o(n_5766) );
no02f02 TIMEBOOST_cell_3186 ( .a(FE_RN_603_0), .b(FE_RN_604_0), .o(TIMEBOOST_net_153) );
in01f02 g59111_u0 ( .a(FE_OCPN1847_n_14981), .o(g59111_sb) );
na02m04 TIMEBOOST_cell_45073 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_411), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_13431) );
no02f02 TIMEBOOST_cell_3187 ( .a(TIMEBOOST_net_153), .b(FE_RN_605_0), .o(FE_RN_606_0) );
na02s01 TIMEBOOST_cell_39733 ( .a(TIMEBOOST_net_11478), .b(g57895_db), .o(n_9229) );
in01f02 g59112_u0 ( .a(FE_OCPN1847_n_14981), .o(g59112_sb) );
in01s01 TIMEBOOST_cell_64267 ( .a(TIMEBOOST_net_21122), .o(TIMEBOOST_net_21123) );
na02f06 TIMEBOOST_cell_3189 ( .a(TIMEBOOST_net_154), .b(n_2558), .o(n_4778) );
na04f04 TIMEBOOST_cell_73227 ( .a(n_1568), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q), .c(FE_OFN713_n_8140), .d(g61940_sb), .o(n_7943) );
in01f02 g59113_u0 ( .a(FE_OCPN1847_n_14981), .o(g59113_sb) );
no02f02 TIMEBOOST_cell_3191 ( .a(TIMEBOOST_net_155), .b(FE_RN_626_0), .o(FE_RN_631_0) );
na02m02 TIMEBOOST_cell_39939 ( .a(TIMEBOOST_net_11581), .b(g62565_sb), .o(n_6427) );
in01s01 TIMEBOOST_cell_67763 ( .a(pci_target_unit_fifos_pcir_data_in_162), .o(TIMEBOOST_net_21190) );
na02m04 TIMEBOOST_cell_68734 ( .a(g65022_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q), .o(TIMEBOOST_net_21575) );
na03f02 TIMEBOOST_cell_70474 ( .a(FE_OFN1695_n_3368), .b(wbu_cache_line_size_in_206), .c(n_3293), .o(TIMEBOOST_net_22445) );
na02s02 TIMEBOOST_cell_39779 ( .a(TIMEBOOST_net_11501), .b(g58003_db), .o(n_9105) );
na03f02 TIMEBOOST_cell_73378 ( .a(TIMEBOOST_net_16702), .b(FE_OFN1300_n_5763), .c(g62044_sb), .o(n_7768) );
na03f02 TIMEBOOST_cell_73442 ( .a(TIMEBOOST_net_17006), .b(FE_OFN1250_n_4093), .c(g62904_sb), .o(n_6069) );
na03f01 TIMEBOOST_cell_67814 ( .a(parchk_pci_ad_reg_in_1220), .b(g67051_sb), .c(TIMEBOOST_net_14100), .o(n_1499) );
in01f04 g59118_u0 ( .a(FE_OCPN1847_n_14981), .o(g59118_sb) );
na03s02 TIMEBOOST_cell_72465 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q), .b(g65865_sb), .c(g65912_db), .o(n_1569) );
na02m02 TIMEBOOST_cell_53893 ( .a(TIMEBOOST_net_7592), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q), .o(TIMEBOOST_net_17164) );
na03s01 TIMEBOOST_cell_64720 ( .a(pci_target_unit_del_sync_addr_in_217), .b(g66406_sb), .c(g66430_db), .o(n_2496) );
na02m06 TIMEBOOST_cell_49539 ( .a(wishbone_slave_unit_pcim_if_wbw_cbe_in), .b(n_691), .o(TIMEBOOST_net_14987) );
na03f02 TIMEBOOST_cell_73715 ( .a(n_12010), .b(TIMEBOOST_net_13564), .c(FE_OFN1746_n_12004), .o(n_12521) );
in01f02 g59121_u0 ( .a(FE_OFN1144_n_15261), .o(g59121_sb) );
na02f02 TIMEBOOST_cell_68158 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q), .b(FE_OFN2054_n_8831), .o(TIMEBOOST_net_21287) );
in01f02 g59122_u0 ( .a(n_8590), .o(g59122_sb) );
na03f02 TIMEBOOST_cell_73051 ( .a(TIMEBOOST_net_22028), .b(FE_OFN710_n_8232), .c(g61795_sb), .o(n_8208) );
na02s01 TIMEBOOST_cell_25608 ( .a(TIMEBOOST_net_6908), .b(n_8746), .o(n_8818) );
in01f02 g59123_u0 ( .a(FE_OFN1697_n_5751), .o(g59123_sb) );
na02s01 TIMEBOOST_cell_38517 ( .a(TIMEBOOST_net_10870), .b(g58202_db), .o(n_9584) );
na03f02 TIMEBOOST_cell_66733 ( .a(TIMEBOOST_net_17116), .b(FE_OFN1314_n_6624), .c(g62988_sb), .o(n_5906) );
na02f02 TIMEBOOST_cell_3633 ( .a(TIMEBOOST_net_376), .b(n_13814), .o(n_7726) );
no02f06 g59124_u0 ( .a(wbu_addr_in_267), .b(n_3203), .o(g59124_p) );
ao12f04 g59124_u1 ( .a(g59124_p), .b(wbu_addr_in_267), .c(n_3203), .o(n_4210) );
no02f04 g59125_u0 ( .a(wbm_adr_o_26_), .b(n_3191), .o(g59125_p) );
ao12f02 g59125_u1 ( .a(g59125_p), .b(wbm_adr_o_26_), .c(n_3191), .o(n_4209) );
in01s01 g59126_u0 ( .a(wbs_rty_o), .o(g59126_sb) );
na02m06 TIMEBOOST_cell_68572 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q), .b(FE_OFN633_n_4454), .o(TIMEBOOST_net_21494) );
na02s01 g59126_u2 ( .a(wbs_rty_o), .b(n_15313), .o(g59126_db) );
no02m04 g59127_u0 ( .a(conf_wb_err_addr_in_959), .b(n_3015), .o(g59127_p) );
ao12m02 g59127_u1 ( .a(g59127_p), .b(conf_wb_err_addr_in_959), .c(n_3015), .o(n_3493) );
no02f02 g59128_u0 ( .a(n_1407), .b(n_4704), .o(g59128_p) );
ao12f02 g59128_u1 ( .a(g59128_p), .b(n_1407), .c(n_4704), .o(n_7095) );
na02m02 TIMEBOOST_cell_48327 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q), .b(g65298_sb), .o(TIMEBOOST_net_14381) );
in01f80 g59133_u0 ( .a(FE_OFN2054_n_8831), .o(n_8665) );
in01f80 g59141_u0 ( .a(n_8665), .o(n_8884) );
no02f04 g59161_u0 ( .a(n_8760), .b(FE_OCP_RBN2003_FE_OFN1026_n_16760), .o(n_14689) );
in01f10 g59169_u0 ( .a(n_8569), .o(n_9372) );
in01s02 TIMEBOOST_cell_62387 ( .a(TIMEBOOST_net_20140), .o(TIMEBOOST_net_20139) );
na02f06 g59175_u0 ( .a(n_1095), .b(n_8590), .o(n_8668) );
na02f04 g59176_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .b(FE_OCPN1847_n_14981), .o(n_8664) );
na02f02 g59177_u0 ( .a(n_3491), .b(wbu_addr_in_275), .o(n_3492) );
no02s01 g59180_u0 ( .a(n_3185), .b(FE_OFN778_n_4152), .o(n_3490) );
no02f01 g59181_u0 ( .a(n_2327), .b(FE_OFN778_n_4152), .o(n_2774) );
na02f02 g59182_u0 ( .a(n_8493), .b(n_1064), .o(n_8494) );
na02f02 g59183_u0 ( .a(n_8493), .b(n_7114), .o(n_8492) );
na02m02 TIMEBOOST_cell_50400 ( .a(TIMEBOOST_net_15417), .b(g62414_sb), .o(n_6770) );
na03m02 TIMEBOOST_cell_73103 ( .a(TIMEBOOST_net_10718), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q), .c(TIMEBOOST_net_16340), .o(TIMEBOOST_net_17423) );
na02f02 TIMEBOOST_cell_70623 ( .a(TIMEBOOST_net_22519), .b(g62860_sb), .o(n_5246) );
no02f06 g59187_u0 ( .a(n_3193), .b(n_1286), .o(n_3489) );
na02s01 TIMEBOOST_cell_25619 ( .a(g61705_sb), .b(g61713_db), .o(TIMEBOOST_net_6914) );
no02f08 g59189_u0 ( .a(n_3190), .b(n_876), .o(n_3488) );
na02f02 TIMEBOOST_cell_70603 ( .a(TIMEBOOST_net_22509), .b(g63015_sb), .o(n_5218) );
ao12f01 g59194_u0 ( .a(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q), .b(n_7715), .c(n_169), .o(n_7720) );
no02m02 g59196_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_15_), .b(n_2491), .o(g59196_p) );
ao12m02 g59196_u1 ( .a(g59196_p), .b(pci_target_unit_del_sync_comp_cycle_count_15_), .c(n_2491), .o(n_3211) );
oa12f02 g59197_u0 ( .a(n_3201), .b(n_3200), .c(wbu_addr_in_271), .o(n_3487) );
no02f02 g59198_u0 ( .a(n_261), .b(n_3179), .o(g59198_p) );
ao12f02 g59198_u1 ( .a(g59198_p), .b(n_261), .c(n_3179), .o(n_4208) );
no02f04 g59199_u0 ( .a(conf_wb_err_addr_in_963), .b(n_2492), .o(g59199_p) );
ao12f02 g59199_u1 ( .a(g59199_p), .b(conf_wb_err_addr_in_963), .c(n_2492), .o(n_3210) );
ao12f02 g59200_u0 ( .a(n_4207), .b(conf_wb_err_addr_in_966), .c(FE_OFN1142_n_15261), .o(n_4886) );
no02f04 g59201_u0 ( .a(conf_wb_err_addr_in_970), .b(n_3353), .o(g59201_p) );
ao12f02 g59201_u1 ( .a(g59201_p), .b(conf_wb_err_addr_in_970), .c(n_3353), .o(n_4707) );
oa12f02 g59202_u0 ( .a(n_3198), .b(n_3197), .c(wbm_adr_o_18_), .o(n_3486) );
oa12f02 g59203_u0 ( .a(n_3196), .b(n_3195), .c(wbm_adr_o_22_), .o(n_3485) );
oa12f02 g59204_u0 ( .a(n_5739), .b(FE_OFN987_n_2696), .c(n_7717), .o(n_7719) );
oa12f02 g59205_u0 ( .a(n_5737), .b(FE_OFN985_n_2697), .c(n_7717), .o(n_7718) );
no02f04 g59206_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q), .b(n_2490), .o(g59206_p) );
ao12f02 g59206_u1 ( .a(g59206_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q), .c(n_2490), .o(n_3209) );
ao12f02 g59208_u0 ( .a(n_3199), .b(conf_wb_err_addr_in_947), .c(FE_OFN1143_n_15261), .o(n_3484) );
in01f02 g59209_u0 ( .a(n_8487), .o(n_8528) );
in01f04 g59211_u0 ( .a(n_2179), .o(n_2180) );
na02m02 TIMEBOOST_cell_53042 ( .a(TIMEBOOST_net_16738), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_15316) );
oa12f01 g59213_u0 ( .a(n_1493), .b(FE_OFN562_n_9895), .c(n_8561), .o(n_8563) );
oa12f02 g59214_u0 ( .a(n_1806), .b(FE_OFN601_n_9687), .c(n_8561), .o(n_8562) );
oa12f02 g59215_u0 ( .a(n_1800), .b(FE_OFN554_n_9864), .c(n_8561), .o(n_8560) );
oa12f02 g59216_u0 ( .a(n_1821), .b(FE_OFN519_n_9697), .c(n_8561), .o(n_8559) );
oa12f02 g59217_u0 ( .a(n_1540), .b(FE_OFN587_n_9692), .c(n_8561), .o(n_8558) );
oa12f02 g59218_u0 ( .a(n_1542), .b(FE_OFN532_n_9823), .c(n_8561), .o(n_8557) );
oa12f02 g59219_u0 ( .a(n_1814), .b(FE_OFN595_n_9694), .c(n_8561), .o(n_8556) );
oa12f02 g59220_u0 ( .a(n_1820), .b(FE_OFN529_n_9899), .c(n_8561), .o(n_8555) );
oa12f02 g59221_u0 ( .a(n_1230), .b(FE_OFN1795_n_9904), .c(n_8561), .o(n_8554) );
oa12f01 g59222_u0 ( .a(n_1822), .b(FE_OFN1800_n_9690), .c(n_8561), .o(n_8553) );
oa12f01 g59223_u0 ( .a(n_1810), .b(FE_OFN577_n_9902), .c(n_8561), .o(n_8552) );
in01f08 g59224_u0 ( .a(n_2175), .o(n_2176) );
in01m01 g59226_u0 ( .a(n_6986), .o(g59226_sb) );
na02f02 g59226_u1 ( .a(wbu_latency_tim_val_in_245), .b(g59226_sb), .o(g59226_da) );
na02m02 TIMEBOOST_cell_40037 ( .a(TIMEBOOST_net_11630), .b(g62564_sb), .o(n_6430) );
in01s01 TIMEBOOST_cell_63596 ( .a(TIMEBOOST_net_20776), .o(TIMEBOOST_net_20749) );
no02f06 g59227_u0 ( .a(wbu_addr_in_263), .b(n_3202), .o(g59227_p) );
ao12f02 g59227_u1 ( .a(g59227_p), .b(wbu_addr_in_263), .c(n_3202), .o(n_3358) );
no02f01 g59228_u0 ( .a(conf_wb_err_addr_in_955), .b(n_3014), .o(g59228_p) );
ao12f02 g59228_u1 ( .a(g59228_p), .b(conf_wb_err_addr_in_955), .c(n_3014), .o(n_3206) );
no02f04 g59229_u0 ( .a(n_3189), .b(wbm_adr_o_14_), .o(g59229_p) );
ao12f02 g59229_u1 ( .a(g59229_p), .b(wbm_adr_o_14_), .c(n_3189), .o(n_3357) );
in01f02 g59230_u0 ( .a(FE_OFN1699_n_5751), .o(g59230_sb) );
na02f01 TIMEBOOST_cell_3639 ( .a(TIMEBOOST_net_379), .b(n_8538), .o(n_8575) );
in01m02 g59231_u0 ( .a(FE_OFN1698_n_5751), .o(g59231_sb) );
na02s01 TIMEBOOST_cell_45591 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q), .o(TIMEBOOST_net_13690) );
na02f01 TIMEBOOST_cell_48100 ( .a(TIMEBOOST_net_14267), .b(FE_OFN787_n_2678), .o(TIMEBOOST_net_12650) );
na02f02 TIMEBOOST_cell_3641 ( .a(TIMEBOOST_net_380), .b(n_8572), .o(n_8573) );
in01s01 TIMEBOOST_cell_67765 ( .a(pci_target_unit_fifos_pcir_data_in_172), .o(TIMEBOOST_net_21192) );
na03f02 TIMEBOOST_cell_73458 ( .a(TIMEBOOST_net_17518), .b(FE_OFN1206_n_6356), .c(g62590_sb), .o(n_6372) );
na02s02 TIMEBOOST_cell_39715 ( .a(TIMEBOOST_net_11469), .b(g58416_db), .o(n_9202) );
in01f02 g59232_u3 ( .a(g59232_p), .o(n_7716) );
oa12f02 g59233_u0 ( .a(n_8480), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309), .c(FE_OFN1651_n_9428), .o(n_8551) );
in01f02 g59234_u0 ( .a(FE_OFN1145_n_15261), .o(g59234_sb) );
na03f01 TIMEBOOST_cell_67974 ( .a(TIMEBOOST_net_15231), .b(FE_OFN1179_n_3476), .c(g60619_sb), .o(n_4835) );
na04f04 TIMEBOOST_cell_24796 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q), .b(g58806_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q), .d(FE_OFN2153_n_16439), .o(n_8635) );
na02m02 TIMEBOOST_cell_68881 ( .a(TIMEBOOST_net_21648), .b(g64795_db), .o(TIMEBOOST_net_17542) );
oa12f02 g59235_u0 ( .a(n_8485), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465), .c(FE_OFN1691_n_9528), .o(n_8550) );
oa12f02 g59236_u0 ( .a(n_8484), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543), .c(FE_OFN1655_n_9502), .o(n_8549) );
oa12f02 g59237_u0 ( .a(n_8482), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582), .c(FE_OFN1667_n_9477), .o(n_8548) );
oa12f02 g59238_u0 ( .a(n_8481), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621), .c(FE_OFN1631_n_9531), .o(n_8547) );
in01m02 g59239_u0 ( .a(FE_OFN999_n_15978), .o(g59239_sb) );
na02f02 TIMEBOOST_cell_71746 ( .a(TIMEBOOST_net_13807), .b(n_13903), .o(TIMEBOOST_net_23081) );
na03s02 TIMEBOOST_cell_41952 ( .a(FE_OFN213_n_9124), .b(g58174_sb), .c(g58174_db), .o(n_9061) );
na03s02 TIMEBOOST_cell_33794 ( .a(n_1573), .b(g61933_sb), .c(g61933_db), .o(n_7957) );
in01f01 g59240_u0 ( .a(FE_OFN1698_n_5751), .o(g59240_sb) );
na02s01 TIMEBOOST_cell_25607 ( .a(TIMEBOOST_net_12), .b(pci_target_unit_wishbone_master_reset_rty_cnt), .o(TIMEBOOST_net_6908) );
na03f02 TIMEBOOST_cell_66065 ( .a(n_3951), .b(g62863_sb), .c(TIMEBOOST_net_7508), .o(n_5240) );
na02f10 TIMEBOOST_cell_47550 ( .a(TIMEBOOST_net_13992), .b(n_1689), .o(TIMEBOOST_net_188) );
in01f02 g59294_u0 ( .a(n_5747), .o(n_7092) );
no02f04 g59296_u0 ( .a(n_8759), .b(pci_target_unit_pcit_if_strd_bc_in_719), .o(g59296_p) );
in01f02 g59296_u1 ( .a(g59296_p), .o(n_8760) );
na02m02 g59297_u0 ( .a(n_8759), .b(wbm_adr_o_0_), .o(n_8880) );
na02m02 g59298_u0 ( .a(n_8759), .b(wbm_adr_o_1_), .o(n_8879) );
no02f02 g59299_u0 ( .a(n_3352), .b(FE_OFN1142_n_15261), .o(n_4207) );
na02f04 g59300_u0 ( .a(n_3202), .b(n_3194), .o(g59300_p) );
in01f04 g59300_u1 ( .a(g59300_p), .o(n_3203) );
in01f06 g59302_u0 ( .a(n_15188), .o(n_7712) );
na02f02 g59309_u0 ( .a(n_3200), .b(wbu_addr_in_271), .o(n_3201) );
in01f01 g59311_u0 ( .a(n_8582), .o(n_8527) );
na02f04 g59312_u0 ( .a(n_7027), .b(n_7624), .o(n_8582) );
na02f01 g59313_u0 ( .a(FE_OFN1691_n_9528), .b(n_8483), .o(n_8485) );
na02f01 g59314_u0 ( .a(FE_OFN1655_n_9502), .b(n_8483), .o(n_8484) );
na03f02 TIMEBOOST_cell_34902 ( .a(TIMEBOOST_net_10009), .b(FE_OFN1422_n_8567), .c(g57482_sb), .o(n_11254) );
na02f01 g59316_u0 ( .a(FE_OFN1667_n_9477), .b(n_8483), .o(n_8482) );
na02f01 g59317_u0 ( .a(FE_OFN1631_n_9531), .b(n_8483), .o(n_8481) );
no02m01 g59318_u0 ( .a(n_2997), .b(FE_OFN778_n_4152), .o(n_3355) );
na02f01 g59319_u0 ( .a(FE_OFN1651_n_9428), .b(n_8483), .o(n_8480) );
no02m08 g59320_u0 ( .a(n_1119), .b(n_3014), .o(n_3015) );
no02f02 g59321_u0 ( .a(n_16738), .b(n_8759), .o(n_14688) );
no02f06 g59322_u0 ( .a(n_1410), .b(n_3014), .o(n_3013) );
no02f04 g59323_u0 ( .a(n_2752), .b(FE_OFN1143_n_15261), .o(n_3199) );
na02f02 g59324_u0 ( .a(n_3197), .b(wbm_adr_o_18_), .o(n_3198) );
na02f02 TIMEBOOST_cell_72283 ( .a(TIMEBOOST_net_23349), .b(g58341_sb), .o(TIMEBOOST_net_9358) );
na02s02 TIMEBOOST_cell_69305 ( .a(TIMEBOOST_net_21860), .b(g65735_sb), .o(n_1608) );
no02f02 g59327_u0 ( .a(n_7322), .b(n_3310), .o(n_8493) );
ao12f04 g59329_u0 ( .a(n_7552), .b(n_7309), .c(n_3036), .o(n_7824) );
in01f02 g59330_u0 ( .a(n_8590), .o(n_8526) );
in01f08 g59331_u1 ( .a(g59331_p), .o(n_8590) );
ao12f02 g59332_u0 ( .a(n_7822), .b(n_7032), .c(n_3033), .o(n_7709) );
na02f04 g59333_u0 ( .a(n_3195), .b(wbm_adr_o_22_), .o(n_3196) );
ao12f02 g59334_u0 ( .a(n_7822), .b(n_7030), .c(n_3055), .o(n_7708) );
ao12f02 g59335_u0 ( .a(n_7822), .b(n_7029), .c(n_3072), .o(n_7707) );
ao12s02 g59336_u0 ( .a(n_2979), .b(n_7047), .c(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_7706) );
na02f02 TIMEBOOST_cell_18291 ( .a(n_1161), .b(n_1162), .o(TIMEBOOST_net_5509) );
na02f02 TIMEBOOST_cell_18224 ( .a(TIMEBOOST_net_5475), .b(n_7538), .o(n_7539) );
in01f08 g59339_u0 ( .a(n_7704), .o(n_7705) );
na02m02 TIMEBOOST_cell_18297 ( .a(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81), .b(n_8757), .o(TIMEBOOST_net_5512) );
ao12f02 g59341_u0 ( .a(n_7822), .b(n_7308), .c(n_2768), .o(n_7823) );
na02f01 TIMEBOOST_cell_26509 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_412), .b(n_13447), .o(TIMEBOOST_net_7359) );
in01f02 g59344_u1 ( .a(g59344_p), .o(n_7551) );
na04f02 TIMEBOOST_cell_36844 ( .a(n_4890), .b(n_8935), .c(TIMEBOOST_net_10018), .d(g52614_sb), .o(n_11857) );
in01f02 g59345_u1 ( .a(g59345_p), .o(n_7550) );
in01s01 TIMEBOOST_cell_73840 ( .a(n_11450), .o(TIMEBOOST_net_23405) );
in01f02 g59346_u1 ( .a(g59346_p), .o(n_7548) );
na04f02 TIMEBOOST_cell_66571 ( .a(n_4889), .b(FE_OFN1698_n_5751), .c(TIMEBOOST_net_684), .d(g52403_db), .o(n_14816) );
in01f02 g59347_u1 ( .a(g59347_p), .o(n_7547) );
ao12f02 g59348_u0 ( .a(n_12595), .b(n_7220), .c(n_3051), .o(n_7702) );
in01f02 g59350_u0 ( .a(FE_OFN1189_n_5742), .o(g59350_sb) );
in01s01 TIMEBOOST_cell_63570 ( .a(TIMEBOOST_net_20750), .o(wbs_adr_i_14_) );
na02f02 TIMEBOOST_cell_69901 ( .a(TIMEBOOST_net_22158), .b(g64187_db), .o(TIMEBOOST_net_16414) );
na02f02 g59351_u0 ( .a(n_7315), .b(n_1105), .o(n_8529) );
na02m02 TIMEBOOST_cell_18295 ( .a(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82), .b(n_8757), .o(TIMEBOOST_net_5511) );
na02f01 TIMEBOOST_cell_72300 ( .a(TIMEBOOST_net_17024), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_23358) );
ao12s01 g59354_u0 ( .a(n_7324), .b(pci_target_unit_del_sync_comp_done_reg_clr), .c(n_2146), .o(n_7699) );
ao12f02 g59355_u0 ( .a(n_7684), .b(n_1069), .c(n_7529), .o(n_7698) );
no02f06 g59356_u0 ( .a(n_1356), .b(n_3197), .o(n_3191) );
na02s02 TIMEBOOST_cell_53374 ( .a(TIMEBOOST_net_16904), .b(FE_OFN1017_n_2053), .o(TIMEBOOST_net_14371) );
oa12f02 g59358_u0 ( .a(n_7079), .b(n_7078), .c(wishbone_slave_unit_pci_initiator_if_read_count_3_), .o(n_7544) );
no02f02 g59359_u0 ( .a(n_7325), .b(n_4188), .o(n_7697) );
ao12f02 g59361_u0 ( .a(n_1536), .b(n_7538), .c(n_3386), .o(n_7543) );
ao12f02 g59362_u0 ( .a(n_7316), .b(n_2999), .c(n_15407), .o(n_7695) );
oa12f02 g59363_u0 ( .a(n_7816), .b(n_6943), .c(FE_OCPN1875_n_14526), .o(n_8525) );
no02m02 g59364_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_14_), .b(n_2478), .o(g59364_p) );
ao12m02 g59364_u1 ( .a(g59364_p), .b(pci_target_unit_del_sync_comp_cycle_count_14_), .c(n_2478), .o(n_3185) );
ao12f02 g59365_u0 ( .a(n_3354), .b(conf_wb_err_addr_in_962), .c(FE_OFN1142_n_15261), .o(n_4206) );
oa12f02 g59366_u0 ( .a(n_5735), .b(FE_OFN1188_n_5742), .c(FE_OFN983_n_2700), .o(n_7542) );
no02m04 g59367_u0 ( .a(n_2474), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q), .o(g59367_p) );
ao12m02 g59367_u1 ( .a(g59367_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q), .c(n_2474), .o(n_3184) );
in01f02 g59368_u0 ( .a(FE_OFN1188_n_5742), .o(g59368_sb) );
na03s02 TIMEBOOST_cell_72968 ( .a(n_1950), .b(g61765_sb), .c(g61765_db), .o(n_8281) );
in01f02 g59369_u0 ( .a(FE_OFN1188_n_5742), .o(g59369_sb) );
na02s01 TIMEBOOST_cell_28947 ( .a(n_1680), .b(wbu_addr_in_253), .o(TIMEBOOST_net_8578) );
na03f02 TIMEBOOST_cell_66450 ( .a(TIMEBOOST_net_17141), .b(FE_OFN1319_n_6436), .c(g62453_sb), .o(n_6691) );
in01f01 g59370_u0 ( .a(FE_OFN1126_g64577_p), .o(g59370_sb) );
na02s01 TIMEBOOST_cell_52408 ( .a(TIMEBOOST_net_16421), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_9492) );
na04f04 TIMEBOOST_cell_73052 ( .a(n_2185), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q), .c(FE_OFN699_n_7845), .d(g61993_sb), .o(n_7909) );
in01m01 g59371_u0 ( .a(FE_OFN1126_g64577_p), .o(g59371_sb) );
na02m02 TIMEBOOST_cell_69880 ( .a(FE_OFN1628_n_4438), .b(n_18), .o(TIMEBOOST_net_22148) );
in01f06 g59372_u0 ( .a(FE_OFN1128_g64577_p), .o(g59372_sb) );
na03f02 TIMEBOOST_cell_66831 ( .a(TIMEBOOST_net_16842), .b(FE_OFN1345_n_8567), .c(g57153_sb), .o(n_10463) );
na03s02 TIMEBOOST_cell_42230 ( .a(g58413_sb), .b(FE_OFN203_n_9228), .c(g58413_db), .o(n_9204) );
na03m06 TIMEBOOST_cell_64553 ( .a(n_3761), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q), .c(FE_OFN1677_n_4655), .o(TIMEBOOST_net_12757) );
in01m01 g59373_u0 ( .a(FE_OFN1126_g64577_p), .o(g59373_sb) );
na03f01 TIMEBOOST_cell_64552 ( .a(n_3741), .b(n_3608), .c(FE_OFN620_n_4490), .o(TIMEBOOST_net_14429) );
na02s02 TIMEBOOST_cell_51315 ( .a(g58186_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q), .o(TIMEBOOST_net_15875) );
no02f04 g59374_u0 ( .a(wbm_adr_o_29_), .b(n_3170), .o(g59374_p) );
ao12f02 g59374_u1 ( .a(g59374_p), .b(wbm_adr_o_29_), .c(n_3170), .o(n_4205) );
ao22f02 g59376_u0 ( .a(n_9175), .b(n_7684), .c(n_7039), .d(n_2763), .o(n_7685) );
no02f01 g59377_u0 ( .a(n_1716), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_), .o(g59377_p) );
ao12f02 g59377_u1 ( .a(g59377_p), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_), .c(n_1716), .o(n_2559) );
in01f01 g59378_u0 ( .a(FE_OFN1126_g64577_p), .o(g59378_sb) );
na02s01 TIMEBOOST_cell_52197 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q), .o(TIMEBOOST_net_16316) );
na03f01 TIMEBOOST_cell_64551 ( .a(n_3752), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q), .c(FE_OFN686_n_4417), .o(TIMEBOOST_net_10494) );
in01m02 g59379_u0 ( .a(FE_OFN1132_g64577_p), .o(g59379_sb) );
na02m02 TIMEBOOST_cell_68577 ( .a(TIMEBOOST_net_21496), .b(n_4473), .o(TIMEBOOST_net_17407) );
na03m02 TIMEBOOST_cell_72700 ( .a(TIMEBOOST_net_21560), .b(FE_OFN649_n_4497), .c(TIMEBOOST_net_22002), .o(TIMEBOOST_net_13250) );
na02m02 TIMEBOOST_cell_68675 ( .a(TIMEBOOST_net_21545), .b(g64998_db), .o(TIMEBOOST_net_17533) );
in01m02 g59380_u0 ( .a(FE_OFN1132_g64577_p), .o(g59380_sb) );
na03f02 TIMEBOOST_cell_65491 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q), .b(FE_OFN712_n_8140), .c(n_1901), .o(TIMEBOOST_net_16468) );
na02f02 TIMEBOOST_cell_70539 ( .a(TIMEBOOST_net_22477), .b(g63122_sb), .o(n_5012) );
na03s02 TIMEBOOST_cell_64550 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q), .b(n_3761), .c(FE_OFN1810_n_4454), .o(TIMEBOOST_net_14682) );
in01f06 g59381_u0 ( .a(FE_OFN1126_g64577_p), .o(g59381_sb) );
na02m02 TIMEBOOST_cell_52910 ( .a(TIMEBOOST_net_16672), .b(g58085_db), .o(TIMEBOOST_net_9546) );
in01f02 g59382_u0 ( .a(FE_OFN1699_n_5751), .o(g59382_sb) );
na02f02 TIMEBOOST_cell_71726 ( .a(TIMEBOOST_net_13795), .b(n_13903), .o(TIMEBOOST_net_23071) );
na02m06 TIMEBOOST_cell_54079 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_123), .o(TIMEBOOST_net_17257) );
na02s01 TIMEBOOST_cell_3975 ( .a(TIMEBOOST_net_547), .b(FE_OCPN1832_n_16949), .o(TIMEBOOST_net_400) );
in01f02 g59383_u0 ( .a(FE_OFN1145_n_15261), .o(g59383_sb) );
na02f01 TIMEBOOST_cell_43512 ( .a(TIMEBOOST_net_12650), .b(g65215_sb), .o(n_2672) );
na02s01 TIMEBOOST_cell_40362 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_), .o(TIMEBOOST_net_11793) );
na04f04 TIMEBOOST_cell_67854 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q), .b(FE_OFN1012_n_4734), .c(TIMEBOOST_net_20831), .d(g60678_sb), .o(TIMEBOOST_net_13052) );
in01f01 g59384_u0 ( .a(n_4936), .o(g59384_sb) );
na02s01 TIMEBOOST_cell_71366 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q), .o(TIMEBOOST_net_22891) );
na03f02 TIMEBOOST_cell_67943 ( .a(TIMEBOOST_net_13086), .b(FE_OFN1126_g64577_p), .c(g59378_sb), .o(n_7683) );
no02f01 g59385_u0 ( .a(wbu_addr_in_259), .b(n_2762), .o(g59385_p) );
ao12f01 g59385_u1 ( .a(g59385_p), .b(wbu_addr_in_259), .c(n_2762), .o(n_3006) );
no02f04 g59386_u0 ( .a(n_2761), .b(wbm_adr_o_10_), .o(g59386_p) );
ao12f02 g59386_u1 ( .a(g59386_p), .b(wbm_adr_o_10_), .c(n_2761), .o(n_3005) );
in01f02 g59387_u0 ( .a(FE_OFN1699_n_5751), .o(g59387_sb) );
na03m04 TIMEBOOST_cell_72492 ( .a(n_3755), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q), .c(TIMEBOOST_net_21555), .o(TIMEBOOST_net_17509) );
na03f02 TIMEBOOST_cell_73555 ( .a(TIMEBOOST_net_17498), .b(FE_OFN1231_n_6391), .c(g62982_sb), .o(n_5918) );
no02f02 g59388_u0 ( .a(n_1406), .b(n_4702), .o(g59388_p) );
ao12f02 g59388_u1 ( .a(g59388_p), .b(n_1406), .c(n_4702), .o(n_4704) );
no02m06 g59389_u0 ( .a(conf_wb_err_addr_in_951), .b(n_2769), .o(g59389_p) );
ao12m02 g59389_u1 ( .a(g59389_p), .b(conf_wb_err_addr_in_951), .c(n_2769), .o(n_2770) );
no02f02 g59588_u0 ( .a(FE_OFN1189_n_5742), .b(n_2933), .o(n_5745) );
oa12f02 g59589_u0 ( .a(n_4859), .b(n_1660), .c(n_5229), .o(n_7333) );
in01f08 g59591_u0 ( .a(n_16437), .o(n_17032) );
in01f04 g59593_u0 ( .a(n_8483), .o(n_8561) );
in01m06 g59594_u0 ( .a(n_8489), .o(n_8483) );
na02f80 g59595_u0 ( .a(n_16435), .b(n_6943), .o(n_8489) );
na02f02 g59596_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1183), .o(n_7673) );
na02f02 g59597_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1184), .o(n_7672) );
na02f02 g59598_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1185), .o(n_7671) );
na02f02 g59599_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1186), .o(n_7669) );
na02m02 g59600_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_5_), .o(n_7535) );
na02f02 g59601_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1168), .o(n_7667) );
na02m02 g59602_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_4_), .o(n_7534) );
na02f02 g59603_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1187), .o(n_7666) );
na02m02 g59604_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_2_), .o(n_7532) );
na02m02 g59605_u0 ( .a(FE_OFN1709_n_4868), .b(pci_ad_o_29_), .o(n_7665) );
na02f02 g59606_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1188), .o(n_7664) );
na02f02 g59607_u0 ( .a(FE_OFN1706_n_4868), .b(parchk_pci_ad_out_in_1189), .o(n_7663) );
na02f02 g59608_u0 ( .a(FE_OFN1706_n_4868), .b(parchk_pci_ad_out_in_1190), .o(n_7661) );
na02f02 g59610_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1192), .o(n_7658) );
na02f02 g59611_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1193), .o(n_7657) );
na02f02 g59612_u0 ( .a(FE_OFN1709_n_4868), .b(parchk_pci_ad_out_in_1194), .o(n_7656) );
na02f02 g59613_u0 ( .a(FE_OFN1709_n_4868), .b(parchk_pci_ad_out_in_1195), .o(n_7655) );
na02f02 g59614_u0 ( .a(FE_OFN1709_n_4868), .b(parchk_pci_ad_out_in_1196), .o(n_7654) );
na02f02 g59615_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1169), .o(n_7653) );
na02f02 g59616_u0 ( .a(FE_OFN1709_n_4868), .b(parchk_pci_ad_out_in_1197), .o(n_7652) );
na02f02 g59617_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in_1170), .o(n_7651) );
na02f02 g59618_u0 ( .a(FE_OFN1705_n_4868), .b(parchk_pci_ad_out_in_1171), .o(n_7650) );
na02f02 g59619_u0 ( .a(FE_OFN1705_n_4868), .b(parchk_pci_ad_out_in_1172), .o(n_7649) );
na02f02 g59620_u0 ( .a(FE_OFN1705_n_4868), .b(parchk_pci_ad_out_in_1173), .o(n_7648) );
na02f02 g59621_u0 ( .a(FE_OFN1705_n_4868), .b(parchk_pci_ad_out_in_1174), .o(n_7647) );
na02f08 g59622_u0 ( .a(n_2762), .b(n_2755), .o(g59622_p) );
in01f08 g59622_u1 ( .a(g59622_p), .o(n_3202) );
na02f04 g59623_u0 ( .a(n_7530), .b(n_7529), .o(g59623_p) );
in01f02 g59623_u1 ( .a(g59623_p), .o(n_7531) );
na02f02 g59624_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1175), .o(n_7528) );
na02f02 g59626_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1176), .o(n_7646) );
na02f10 g59627_u0 ( .a(n_2761), .b(n_2756), .o(g59627_p) );
in01f08 g59627_u1 ( .a(g59627_p), .o(n_3189) );
na02m02 g59628_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_26_), .o(n_7527) );
na02s02 g59629_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_23_), .o(n_7525) );
na02s02 g59630_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_20_), .o(n_7524) );
na02m02 g59632_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_0_), .o(n_7523) );
na02m02 g59633_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_13_), .o(n_7522) );
na02m02 g59634_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_14_), .o(n_7521) );
na02s02 g59635_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_15_), .o(n_7519) );
na02m02 g59636_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_17_), .o(n_7518) );
na02m02 g59637_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_18_), .o(n_7645) );
na02s02 g59638_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_19_), .o(n_7643) );
na02m02 g59639_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_1_), .o(n_7517) );
na02m02 g59640_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_21_), .o(n_7516) );
na02s02 g59641_u0 ( .a(FE_OFN1706_n_4868), .b(pci_ad_o_22_), .o(n_7515) );
na02m02 g59642_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_24_), .o(n_7514) );
na02m02 g59643_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_25_), .o(n_7642) );
na02m02 g59644_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_27_), .o(n_7640) );
na02m02 g59645_u0 ( .a(FE_OFN1709_n_4868), .b(pci_ad_o_28_), .o(n_7639) );
na02m02 g59646_u0 ( .a(FE_OFN1709_n_4868), .b(pci_ad_o_30_), .o(n_7513) );
na02m02 g59647_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_3_), .o(n_7512) );
na02m02 g59648_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_6_), .o(n_7511) );
na02m02 g59649_u0 ( .a(FE_OFN1710_n_4868), .b(pci_ad_o_7_), .o(n_7638) );
na02s02 g59650_u0 ( .a(FE_OFN1708_n_4868), .b(pci_ad_o_8_), .o(n_7510) );
na02s02 g59651_u0 ( .a(FE_OFN1708_n_4868), .b(pci_ad_o_9_), .o(n_7637) );
na02f10 g59652_u0 ( .a(n_1270), .b(n_2769), .o(n_3014) );
no02f02 g59653_u0 ( .a(n_2986), .b(FE_OFN1142_n_15261), .o(n_3354) );
na03f02 TIMEBOOST_cell_66918 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_16494), .c(FE_OFN1513_n_14987), .o(n_12624) );
no02f01 g59655_u0 ( .a(n_2304), .b(FE_OFN778_n_4152), .o(n_2757) );
na02s02 g59656_u0 ( .a(FE_OFN1708_n_4868), .b(pci_ad_o_10_), .o(n_7636) );
na02s02 g59657_u0 ( .a(FE_OFN1708_n_4868), .b(pci_ad_o_11_), .o(n_7509) );
na02f02 g59658_u0 ( .a(FE_OFN1189_n_5742), .b(n_7329), .o(n_7330) );
no02f02 g59659_u0 ( .a(n_16435), .b(n_2134), .o(g59659_p) );
in01f02 g59659_u1 ( .a(g59659_p), .o(n_7508) );
na02m02 TIMEBOOST_cell_68485 ( .a(TIMEBOOST_net_21450), .b(TIMEBOOST_net_16169), .o(TIMEBOOST_net_17491) );
no02f02 g59664_u0 ( .a(FE_OFN1189_n_5742), .b(n_1826), .o(n_5743) );
na02m02 g59665_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_hit_2_), .o(g59665_p) );
in01f02 g59665_u1 ( .a(g59665_p), .o(n_5741) );
na02m02 g59666_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_hit_3_), .o(g59666_p) );
in01f02 g59666_u1 ( .a(g59666_p), .o(n_5740) );
na02f04 g59667_u0 ( .a(TIMEBOOST_net_20763), .b(n_5725), .o(n_7717) );
na02f01 g59668_u0 ( .a(FE_OFN1188_n_5742), .b(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q), .o(n_5739) );
na02f01 g59669_u0 ( .a(FE_OFN1188_n_5742), .b(wishbone_slave_unit_wishbone_slave_pref_en_reg_Q), .o(n_5737) );
na02f02 g59670_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(g59670_p) );
in01f01 g59670_u1 ( .a(g59670_p), .o(n_5736) );
na02f02 g59671_u0 ( .a(FE_OFN1710_n_4868), .b(parchk_pci_ad_out_in), .o(n_7635) );
na02f02 g59672_u0 ( .a(FE_OFN1188_n_5742), .b(wishbone_slave_unit_wishbone_slave_map), .o(n_5735) );
na02m02 TIMEBOOST_cell_49472 ( .a(TIMEBOOST_net_14953), .b(FE_OFN1635_n_9531), .o(TIMEBOOST_net_11183) );
na02m02 g59674_u0 ( .a(FE_OFN1189_n_5742), .b(wishbone_slave_unit_wishbone_slave_img_hit_4_), .o(g59674_p) );
in01f02 g59674_u1 ( .a(g59674_p), .o(n_5733) );
na02f02 g59676_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1177), .o(n_7634) );
na02f02 g59677_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1178), .o(n_7633) );
ao12f02 g59678_u0 ( .a(n_7552), .b(n_4691), .c(n_2906), .o(n_7091) );
na02f02 g59679_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1179), .o(n_7632) );
na02f02 g59681_u0 ( .a(FE_OFN1708_n_4868), .b(parchk_pci_ad_out_in_1180), .o(n_7631) );
na02f02 g59682_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1181), .o(n_7630) );
na02m02 g59683_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_16_), .o(n_7629) );
na02f02 g59684_u0 ( .a(FE_OFN1707_n_4868), .b(parchk_pci_ad_out_in_1182), .o(n_7628) );
na02m02 g59685_u0 ( .a(FE_OFN1707_n_4868), .b(pci_ad_o_12_), .o(n_7505) );
na02m02 TIMEBOOST_cell_68660 ( .a(FE_OFN689_n_4438), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_21538) );
na03f02 TIMEBOOST_cell_73228 ( .a(TIMEBOOST_net_22133), .b(FE_OFN710_n_8232), .c(g61813_sb), .o(n_8166) );
na04f04 TIMEBOOST_cell_36851 ( .a(n_9756), .b(g57163_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q), .d(FE_OFN1417_n_8567), .o(n_11587) );
na02m02 TIMEBOOST_cell_53012 ( .a(TIMEBOOST_net_16723), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_15296) );
na04m08 TIMEBOOST_cell_67172 ( .a(n_3792), .b(FE_OFN672_n_4505), .c(g64754_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q), .o(n_3789) );
na02m02 TIMEBOOST_cell_53853 ( .a(n_4302), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q), .o(TIMEBOOST_net_17144) );
no02f02 g59694_u0 ( .a(FE_OFN1189_n_5742), .b(n_2709), .o(n_5732) );
ao12f02 g59695_u0 ( .a(n_12595), .b(n_4819), .c(n_3066), .o(n_7084) );
ao12f02 g59696_u0 ( .a(n_7552), .b(n_4820), .c(n_3064), .o(n_7083) );
ao12f02 g59697_u0 ( .a(n_7552), .b(n_4823), .c(n_3061), .o(n_7082) );
ao12f02 g59698_u0 ( .a(n_7552), .b(n_4824), .c(n_3045), .o(n_7081) );
ao12f02 g59699_u0 ( .a(n_7552), .b(n_4825), .c(n_3059), .o(n_7080) );
in01f20 g59702_u0 ( .a(n_8759), .o(n_14839) );
in01f20 g59716_u0 ( .a(n_8759), .o(n_8757) );
in01f20 g59717_u0 ( .a(n_14837), .o(n_8759) );
in01f10 g59718_u0 ( .a(n_16475), .o(n_14837) );
na02f02 TIMEBOOST_cell_49398 ( .a(TIMEBOOST_net_14916), .b(g61919_sb), .o(n_7983) );
in01f02 g59721_u1 ( .a(g59721_p), .o(n_7821) );
ao12s01 g59723_u0 ( .a(wbu_pci_drcomp_pending_in), .b(pci_target_unit_del_sync_comp_in), .c(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_7324) );
na04f04 TIMEBOOST_cell_24231 ( .a(n_9544), .b(g57392_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q), .d(FE_OFN1406_n_8567), .o(n_11350) );
ao12f02 g59726_u0 ( .a(n_3157), .b(n_2289), .c(wbm_rty_i), .o(n_2998) );
ao12f02 g59727_u0 ( .a(n_7822), .b(n_4899), .c(n_3043), .o(n_7320) );
na02s02 TIMEBOOST_cell_38437 ( .a(TIMEBOOST_net_10830), .b(g57944_db), .o(n_9869) );
in01f02 g59730_u0 ( .a(n_7715), .o(n_7317) );
oa12f04 g59731_u0 ( .a(n_3402), .b(n_4717), .c(n_2888), .o(n_7715) );
na02m02 TIMEBOOST_cell_18293 ( .a(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83), .b(n_8757), .o(TIMEBOOST_net_5510) );
oa12f02 g59734_u0 ( .a(n_2616), .b(FE_OCPN1836_n_16798), .c(n_1435), .o(n_7316) );
oa12f02 g59735_u0 ( .a(n_7313), .b(n_7818), .c(n_8540), .o(n_7627) );
na03f02 TIMEBOOST_cell_73459 ( .a(TIMEBOOST_net_17363), .b(FE_OFN1288_n_4098), .c(g62714_sb), .o(n_6142) );
na02m02 TIMEBOOST_cell_70173 ( .a(TIMEBOOST_net_22294), .b(g60675_sb), .o(n_7226) );
oa12f02 g59738_u0 ( .a(n_7311), .b(n_1758), .c(n_3123), .o(n_7626) );
oa12f02 g59739_u0 ( .a(n_7074), .b(FE_OFN732_n_7498), .c(n_2075), .o(n_7500) );
oa12f02 g59740_u0 ( .a(n_7073), .b(FE_OFN732_n_7498), .c(n_2067), .o(n_7499) );
oa12f02 g59741_u0 ( .a(n_7071), .b(FE_OFN732_n_7498), .c(n_2077), .o(n_7497) );
oa12f01 g59742_u0 ( .a(n_7475), .b(n_7818), .c(n_8517), .o(n_7820) );
oa12f02 g59743_u0 ( .a(n_7069), .b(FE_OFN732_n_7498), .c(n_2082), .o(n_7496) );
oa12f02 g59744_u0 ( .a(n_7070), .b(FE_OFN732_n_7498), .c(n_2069), .o(n_7495) );
oa12f02 g59745_u0 ( .a(n_7068), .b(n_7498), .c(n_2076), .o(n_7494) );
oa12f01 g59746_u0 ( .a(n_7474), .b(n_7818), .c(n_2464), .o(n_7819) );
oa12s02 g59747_u0 ( .a(n_7067), .b(n_7498), .c(n_2068), .o(n_7493) );
oa12f01 g59748_u0 ( .a(n_7472), .b(n_7818), .c(n_2319), .o(n_7817) );
oa12f02 g59749_u0 ( .a(n_7066), .b(n_7498), .c(n_2083), .o(n_7492) );
oa12f02 g59750_u0 ( .a(n_7064), .b(n_7498), .c(n_2286), .o(n_7491) );
oa12f02 g59751_u0 ( .a(n_7063), .b(n_7498), .c(n_2080), .o(n_7490) );
oa12f02 g59752_u0 ( .a(n_7062), .b(n_7498), .c(n_2079), .o(n_7489) );
oa12f02 g59753_u0 ( .a(n_7061), .b(n_7498), .c(n_2072), .o(n_7488) );
oa12f02 g59754_u0 ( .a(n_7060), .b(n_7498), .c(n_2070), .o(n_7487) );
oa12f02 g59755_u0 ( .a(n_7059), .b(n_7498), .c(n_8540), .o(n_7486) );
oa12f02 g59756_u0 ( .a(n_7057), .b(FE_OFN732_n_7498), .c(n_1737), .o(n_7485) );
oa12f02 g59757_u0 ( .a(n_7058), .b(n_7498), .c(n_3280), .o(n_7484) );
oa12f02 g59758_u0 ( .a(n_7613), .b(n_8476), .c(n_8517), .o(n_8478) );
oa12f02 g59759_u0 ( .a(n_7610), .b(n_8476), .c(n_2319), .o(n_8477) );
oa12f02 g59760_u0 ( .a(n_7612), .b(n_8476), .c(n_2464), .o(n_8474) );
no02f04 g59761_u0 ( .a(conf_wb_err_addr_in_966), .b(n_2983), .o(g59761_p) );
ao12f02 g59761_u1 ( .a(g59761_p), .b(conf_wb_err_addr_in_966), .c(n_2983), .o(n_3352) );
oa12f02 g59762_u0 ( .a(n_2992), .b(n_2991), .c(wbu_addr_in_274), .o(n_3351) );
in01f02 g59763_u0 ( .a(FE_OFN1330_n_13547), .o(g59763_sb) );
in01s01 TIMEBOOST_cell_67782 ( .a(TIMEBOOST_net_21208), .o(TIMEBOOST_net_21209) );
na02s01 TIMEBOOST_cell_3966 ( .a(n_12179), .b(n_657), .o(TIMEBOOST_net_543) );
na03f02 TIMEBOOST_cell_73611 ( .a(TIMEBOOST_net_13366), .b(n_6287), .c(g62964_sb), .o(n_5954) );
oa12f02 g59764_u0 ( .a(n_7815), .b(n_8521), .c(n_2464), .o(n_8523) );
ao12f02 g59765_u0 ( .a(n_4696), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .c(FE_OFN1144_n_15261), .o(n_5731) );
oa12m02 g59766_u0 ( .a(n_7814), .b(n_8521), .c(n_2319), .o(n_8522) );
ao12f02 g59767_u0 ( .a(n_3475), .b(conf_wb_err_addr_in_969), .c(FE_OFN1144_n_15261), .o(n_4700) );
ao12f02 g59768_u0 ( .a(n_3172), .b(conf_wb_err_addr_in_950), .c(FE_OFN1142_n_15261), .o(n_3479) );
oa12f02 g59769_u0 ( .a(n_2990), .b(n_2989), .c(wbm_adr_o_17_), .o(n_3350) );
na02f02 TIMEBOOST_cell_49904 ( .a(TIMEBOOST_net_15169), .b(g63021_sb), .o(n_5205) );
na02s02 TIMEBOOST_cell_38270 ( .a(g57909_sb), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_10747) );
oa12f01 g59771_u0 ( .a(n_3455), .b(n_2034), .c(n_4662), .o(n_4202) );
oa12f02 g59772_u0 ( .a(FE_OCPN1875_n_14526), .b(n_7096), .c(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_7816) );
oa12f02 g59773_u0 ( .a(n_3175), .b(n_3174), .c(wbm_adr_o_25_), .o(n_3478) );
oa12f02 g59774_u0 ( .a(n_7055), .b(FE_OFN732_n_7498), .c(n_1743), .o(n_7483) );
oa12f02 g59775_u0 ( .a(n_7054), .b(FE_OFN732_n_7498), .c(n_2041), .o(n_7482) );
oa12f02 g59776_u0 ( .a(n_7053), .b(FE_OFN732_n_7498), .c(n_2040), .o(n_7481) );
oa12f02 g59777_u0 ( .a(n_7052), .b(FE_OFN732_n_7498), .c(n_1746), .o(n_7480) );
oa12f02 g59778_u0 ( .a(n_7051), .b(FE_OFN732_n_7498), .c(n_2052), .o(n_7479) );
oa12f02 g59779_u0 ( .a(n_7050), .b(FE_OFN732_n_7498), .c(n_1740), .o(n_7478) );
oa12f02 g59780_u0 ( .a(n_7049), .b(FE_OFN732_n_7498), .c(n_2074), .o(n_7477) );
oa12f02 g59781_u0 ( .a(n_7048), .b(FE_OFN732_n_7498), .c(n_2084), .o(n_7476) );
na02m06 TIMEBOOST_cell_70271 ( .a(TIMEBOOST_net_22343), .b(TIMEBOOST_net_13119), .o(TIMEBOOST_net_16840) );
no02m04 g59783_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_11_), .b(n_2421), .o(g59783_p) );
ao12m02 g59783_u1 ( .a(g59783_p), .b(pci_target_unit_del_sync_comp_cycle_count_11_), .c(n_2421), .o(n_2997) );
ao12f02 g59784_u0 ( .a(n_3173), .b(conf_wb_err_addr_in_946), .c(FE_OFN1143_n_15261), .o(n_3477) );
no02f04 g59785_u0 ( .a(n_193), .b(n_2425), .o(g59785_p) );
ao12f02 g59785_u1 ( .a(g59785_p), .b(n_193), .c(n_2425), .o(n_2996) );
ao22m06 g59786_u0 ( .a(n_5642), .b(n_13447), .c(FE_OFN1619_n_1787), .d(conf_wb_err_bc_in_846), .o(n_7315) );
na03m02 TIMEBOOST_cell_69900 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(g64187_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q), .o(TIMEBOOST_net_22158) );
in01m02 g59788_u0 ( .a(n_4883), .o(n_5730) );
ao22f02 g59789_u0 ( .a(n_925), .b(n_72), .c(n_4694), .d(configuration_icr_bit_2967), .o(n_4883) );
no02f01 g59790_u0 ( .a(conf_wb_err_addr_in_947), .b(n_2035), .o(g59790_p) );
ao12f01 g59790_u1 ( .a(g59790_p), .b(conf_wb_err_addr_in_947), .c(n_2035), .o(n_2752) );
no02f01 g59791_u0 ( .a(wbu_addr_in_255), .b(n_2487), .o(g59791_p) );
ao12m01 g59791_u1 ( .a(g59791_p), .b(wbu_addr_in_255), .c(n_2487), .o(n_2488) );
ao22f02 g59792_u0 ( .a(n_2405), .b(n_7078), .c(n_2014), .d(n_5228), .o(n_7079) );
no02m02 g59793_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_4_), .b(n_1693), .o(g59793_p) );
ao12m02 g59793_u1 ( .a(g59793_p), .b(pci_target_unit_del_sync_comp_cycle_count_4_), .c(n_1693), .o(n_2327) );
no02f01 g59794_u0 ( .a(n_2485), .b(wbm_adr_o_6_), .o(g59794_p) );
ao12f01 g59794_u1 ( .a(g59794_p), .b(wbm_adr_o_6_), .c(n_2485), .o(n_2486) );
no02f01 g59795_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_4_), .b(n_1695), .o(g59795_p) );
ao12m01 g59795_u1 ( .a(g59795_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_4_), .c(n_1695), .o(n_2326) );
in01f01 g59796_u0 ( .a(n_13547), .o(g59796_sb) );
na02f01 g59796_u2 ( .a(n_5641), .b(n_13547), .o(g59796_db) );
na02m10 TIMEBOOST_cell_53001 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q), .b(wishbone_slave_unit_pcim_sm_data_in_655), .o(TIMEBOOST_net_16718) );
in01m02 g59797_u0 ( .a(FE_OFN1698_n_5751), .o(g59797_sb) );
in01s01 TIMEBOOST_cell_45867 ( .a(TIMEBOOST_net_13935), .o(TIMEBOOST_net_13828) );
na03f02 TIMEBOOST_cell_68014 ( .a(TIMEBOOST_net_17520), .b(FE_OFN1250_n_4093), .c(g62581_sb), .o(n_6390) );
na02f08 TIMEBOOST_cell_3645 ( .a(TIMEBOOST_net_382), .b(n_7108), .o(n_8468) );
in01m02 g59798_u0 ( .a(FE_OFN1700_n_5751), .o(g59798_sb) );
na02s01 TIMEBOOST_cell_45391 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q), .o(TIMEBOOST_net_13590) );
na02m10 TIMEBOOST_cell_45357 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q), .o(TIMEBOOST_net_13573) );
no02f02 TIMEBOOST_cell_3973 ( .a(TIMEBOOST_net_546), .b(n_3126), .o(g63307_p) );
in01f02 g59799_u0 ( .a(FE_OFN1083_n_13221), .o(g59799_sb) );
na03m02 TIMEBOOST_cell_64547 ( .a(n_3764), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q), .c(FE_OFN689_n_4438), .o(TIMEBOOST_net_16201) );
in01f01 g59800_u0 ( .a(FE_OFN1697_n_5751), .o(g59800_sb) );
na02f02 g59800_u2 ( .a(n_2739), .b(FE_OFN1697_n_5751), .o(g59800_db) );
na02s01 TIMEBOOST_cell_39787 ( .a(TIMEBOOST_net_11505), .b(g58063_db), .o(n_9089) );
in01f02 g59801_u0 ( .a(FE_OFN1697_n_5751), .o(g59801_sb) );
na03m02 TIMEBOOST_cell_66364 ( .a(TIMEBOOST_net_13385), .b(g54182_sb), .c(g54182_db), .o(n_13431) );
no02f04 g59802_u0 ( .a(conf_wb_err_addr_in_958), .b(n_2751), .o(g59802_p) );
ao12f02 g59802_u1 ( .a(g59802_p), .b(conf_wb_err_addr_in_958), .c(n_2751), .o(n_3347) );
no02f08 g59803_u0 ( .a(wbu_addr_in_266), .b(n_2968), .o(g59803_p) );
ao12f04 g59803_u1 ( .a(g59803_p), .b(wbu_addr_in_266), .c(n_2968), .o(n_3346) );
in01f02 g59804_u0 ( .a(n_7618), .o(g59804_sb) );
na02m02 TIMEBOOST_cell_70765 ( .a(TIMEBOOST_net_22590), .b(g52399_sb), .o(TIMEBOOST_net_8849) );
na02m01 TIMEBOOST_cell_71904 ( .a(FE_OFN665_n_4495), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q), .o(TIMEBOOST_net_23160) );
na02f02 TIMEBOOST_cell_69372 ( .a(wbu_latency_tim_val_in_243), .b(n_6986), .o(TIMEBOOST_net_21894) );
in01f02 g59805_u0 ( .a(n_7618), .o(g59805_sb) );
na02s01 TIMEBOOST_cell_37616 ( .a(g58145_sb), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_10420) );
na02f01 TIMEBOOST_cell_44336 ( .a(TIMEBOOST_net_13062), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_11348) );
in01s01 TIMEBOOST_cell_45868 ( .a(TIMEBOOST_net_13828), .o(TIMEBOOST_net_13829) );
in01f02 g59806_u0 ( .a(n_7618), .o(g59806_sb) );
na02f01 TIMEBOOST_cell_26071 ( .a(pci_target_unit_pcit_if_strd_addr_in_699), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7140) );
na04m02 TIMEBOOST_cell_67199 ( .a(TIMEBOOST_net_20182), .b(FE_OFN903_n_4736), .c(g60677_sb), .d(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q), .o(TIMEBOOST_net_13065) );
in01f02 g59807_u0 ( .a(n_7618), .o(g59807_sb) );
na04f04 TIMEBOOST_cell_24653 ( .a(n_9711), .b(g57225_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q), .d(FE_OFN2189_n_8567), .o(n_11531) );
na02f01 TIMEBOOST_cell_48102 ( .a(TIMEBOOST_net_14268), .b(FE_OFN787_n_2678), .o(TIMEBOOST_net_12647) );
na04f04 TIMEBOOST_cell_24651 ( .a(n_9707), .b(g57230_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q), .d(FE_OFN2179_n_8567), .o(n_11524) );
in01f02 g59808_u0 ( .a(n_7618), .o(g59808_sb) );
na03f02 TIMEBOOST_cell_69642 ( .a(TIMEBOOST_net_14164), .b(TIMEBOOST_net_10248), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_22029) );
na02f02 TIMEBOOST_cell_49814 ( .a(TIMEBOOST_net_15124), .b(g62774_sb), .o(n_5446) );
in01f02 g59809_u0 ( .a(n_7618), .o(g59809_sb) );
na02m02 TIMEBOOST_cell_48104 ( .a(TIMEBOOST_net_14269), .b(TIMEBOOST_net_10321), .o(TIMEBOOST_net_9454) );
na02s01 TIMEBOOST_cell_68524 ( .a(g58025_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q), .o(TIMEBOOST_net_21470) );
in01f02 g59_u0 ( .a(n_15538), .o(n_15539) );
na02f01 TIMEBOOST_cell_18205 ( .a(n_2407), .b(n_7078), .o(TIMEBOOST_net_5466) );
na02f01 TIMEBOOST_cell_18208 ( .a(TIMEBOOST_net_5467), .b(FE_OCPN1836_n_16798), .o(TIMEBOOST_net_399) );
na03f02 TIMEBOOST_cell_66856 ( .a(TIMEBOOST_net_20666), .b(n_14971), .c(g58640_sb), .o(n_9238) );
na02f02 TIMEBOOST_cell_18207 ( .a(n_15405), .b(n_13745), .o(TIMEBOOST_net_5467) );
na02f02 g60264_u0 ( .a(n_7072), .b(pciu_bar1_in_389), .o(n_7074) );
na02f02 g60265_u0 ( .a(n_7072), .b(pciu_bar1_in_390), .o(n_7073) );
na02f02 g60266_u0 ( .a(n_7072), .b(pciu_bar1_in_391), .o(n_7071) );
na02f02 g60267_u0 ( .a(n_7072), .b(pciu_bar1_in_392), .o(n_7070) );
na02f02 g60268_u0 ( .a(n_7072), .b(pciu_bar1_in_393), .o(n_7069) );
na02f02 g60269_u0 ( .a(n_7072), .b(pciu_bar1_in_394), .o(n_7068) );
na02f02 g60270_u0 ( .a(n_7473), .b(configuration_icr_bit2_0), .o(n_7475) );
na02f02 g60271_u0 ( .a(n_7065), .b(pciu_bar1_in_395), .o(n_7067) );
na02f02 g60272_u0 ( .a(n_7065), .b(pciu_bar1_in_396), .o(n_7066) );
na02f02 g60273_u0 ( .a(n_7473), .b(configuration_icr_bit_2961), .o(n_7474) );
na02f02 g60274_u0 ( .a(n_7065), .b(pciu_bar1_in_397), .o(n_7064) );
na02f02 g60275_u0 ( .a(n_7473), .b(configuration_icr_bit_2967), .o(n_7472) );
na02f02 g60276_u0 ( .a(n_7065), .b(pciu_bar1_in_398), .o(n_7063) );
na02f02 g60277_u0 ( .a(n_7065), .b(pciu_bar1_in_399), .o(n_7062) );
oa12f01 g60278_u0 ( .a(pci_resi_conf_soft_res_in), .b(n_7818), .c(n_8511), .o(n_7313) );
na02f02 g60279_u0 ( .a(n_7065), .b(pciu_bar1_in_400), .o(n_7061) );
na02f02 g60280_u0 ( .a(n_7065), .b(pciu_bar1_in_401), .o(n_7060) );
na02f02 g60281_u0 ( .a(n_7065), .b(pciu_bar1_in_402), .o(n_7059) );
na02f02 g60282_u0 ( .a(n_7056), .b(pciu_bar1_in), .o(n_7058) );
na02f02 g60283_u0 ( .a(n_7056), .b(pciu_bar1_in_380), .o(n_7057) );
na02f03 g60284_u0 ( .a(n_7611), .b(wbu_mrl_en_in_141), .o(n_7613) );
na02f03 g60285_u0 ( .a(n_7611), .b(wbu_pref_en_in_136), .o(n_7612) );
na02f03 g60286_u0 ( .a(n_7611), .b(n_14907), .o(n_7610) );
na02f02 g60287_u0 ( .a(n_7813), .b(pciu_pref_en_in_320), .o(n_7815) );
na02f01 g60288_u0 ( .a(n_7813), .b(n_14910), .o(n_7814) );
na02f02 g60289_u0 ( .a(n_7056), .b(pciu_bar1_in_381), .o(n_7055) );
na02f02 g60290_u0 ( .a(n_7056), .b(pciu_bar1_in_382), .o(n_7054) );
na02f02 g60291_u0 ( .a(n_7056), .b(pciu_bar1_in_383), .o(n_7053) );
na02f02 g60292_u0 ( .a(n_7056), .b(pciu_bar1_in_384), .o(n_7052) );
na02f02 g60293_u0 ( .a(n_7056), .b(pciu_bar1_in_385), .o(n_7051) );
na02f02 g60294_u0 ( .a(n_7056), .b(pciu_bar1_in_386), .o(n_7050) );
na02f02 g60295_u0 ( .a(n_7072), .b(pciu_bar1_in_387), .o(n_7049) );
na02f02 g60296_u0 ( .a(n_7072), .b(pciu_bar1_in_388), .o(n_7048) );
na02f04 g60297_u0 ( .a(n_3174), .b(wbm_adr_o_25_), .o(n_3175) );
no02f02 g60298_u0 ( .a(pci_target_unit_del_sync_comp_in), .b(n_4177), .o(g60298_p) );
in01f02 g60298_u1 ( .a(g60298_p), .o(n_7047) );
na03f02 TIMEBOOST_cell_72244 ( .a(n_3922), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q), .c(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_23330) );
no02f08 g60303_u0 ( .a(n_2476), .b(n_2750), .o(n_2993) );
na02f08 g60304_u0 ( .a(n_2306), .b(n_2487), .o(g60304_p) );
in01f06 g60304_u1 ( .a(g60304_p), .o(n_2762) );
ao12f02 g60305_u0 ( .a(n_7552), .b(n_4803), .c(n_2853), .o(n_7046) );
ao12f02 g60306_u0 ( .a(n_12595), .b(n_4802), .c(n_2848), .o(n_7045) );
na02f02 g60307_u0 ( .a(FE_OCPN1836_n_16798), .b(n_7044), .o(g60307_p) );
in01f02 g60307_u1 ( .a(g60307_p), .o(n_7529) );
na02f04 g60308_u0 ( .a(n_2991), .b(wbu_addr_in_274), .o(n_2992) );
in01f02 g60309_u0 ( .a(n_7310), .o(n_7311) );
na02f04 g60310_u0 ( .a(FE_OCPN1836_n_16798), .b(n_9175), .o(g60310_p) );
in01f02 g60310_u1 ( .a(g60310_p), .o(n_7310) );
na03m04 TIMEBOOST_cell_72821 ( .a(g65336_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q), .c(TIMEBOOST_net_16626), .o(TIMEBOOST_net_13366) );
na02f02 g60312_u0 ( .a(n_2343), .b(n_16452), .o(n_7043) );
in01f01 g60314_u0 ( .a(n_7040), .o(n_7039) );
na02f02 g60315_u0 ( .a(n_16798), .b(n_15407), .o(n_7040) );
no02f20 g60318_u0 ( .a(n_1972), .b(n_2035), .o(n_2769) );
na02f20 g60319_u0 ( .a(n_2485), .b(n_2305), .o(g60319_p) );
in01f10 g60319_u1 ( .a(g60319_p), .o(n_2761) );
no02f02 g60320_u0 ( .a(n_3344), .b(FE_OFN1144_n_15261), .o(n_3475) );
na02f01 g60321_u0 ( .a(n_1714), .b(n_1715), .o(g60321_p) );
in01f02 g60321_u1 ( .a(g60321_p), .o(n_1716) );
no02f02 g60322_u0 ( .a(n_4162), .b(FE_OFN1144_n_15261), .o(n_4696) );
no02f04 g60323_u0 ( .a(n_2272), .b(FE_OFN1143_n_15261), .o(n_3173) );
no02f04 g60324_u0 ( .a(n_2981), .b(FE_OFN1142_n_15261), .o(n_3172) );
na02f02 g60325_u0 ( .a(n_2989), .b(wbm_adr_o_17_), .o(n_2990) );
no02f01 g60326_u0 ( .a(n_2024), .b(FE_OFN778_n_4152), .o(n_2748) );
na03m06 TIMEBOOST_cell_64546 ( .a(n_3747), .b(FE_OFN686_n_4417), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q), .o(TIMEBOOST_net_14288) );
in01f04 g60328_u0 ( .a(n_15446), .o(n_7038) );
na02f02 g60330_u0 ( .a(FE_OCPN1836_n_16798), .b(pci_target_unit_pci_target_sm_cnf_progress), .o(g60330_p) );
in01f02 g60330_u1 ( .a(g60330_p), .o(n_7684) );
no02f04 g60331_u0 ( .a(n_5728), .b(n_7031), .o(n_7309) );
no02m01 g60333_u0 ( .a(n_2964), .b(FE_OFN778_n_4152), .o(n_3171) );
in01f02 g60335_u0 ( .a(FE_OFN1188_n_5742), .o(n_5725) );
na02m02 TIMEBOOST_cell_68579 ( .a(TIMEBOOST_net_21497), .b(TIMEBOOST_net_10397), .o(TIMEBOOST_net_20578) );
na03f02 TIMEBOOST_cell_73229 ( .a(g64100_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q), .c(TIMEBOOST_net_14874), .o(TIMEBOOST_net_15103) );
in01f02 g60339_u1 ( .a(g60339_p), .o(n_7307) );
ao12f02 g60340_u0 ( .a(n_5643), .b(n_16000), .c(n_2856), .o(n_7033) );
in01s01 TIMEBOOST_cell_73975 ( .a(TIMEBOOST_net_23539), .o(TIMEBOOST_net_23540) );
na04f04 TIMEBOOST_cell_25012 ( .a(n_9332), .b(n_11008), .c(n_9331), .d(n_10235), .o(n_12165) );
oa12f01 g60343_u0 ( .a(n_4591), .b(n_3437), .c(n_4869), .o(n_4870) );
na02m10 TIMEBOOST_cell_45773 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q), .o(TIMEBOOST_net_13781) );
no02f01 g60345_u0 ( .a(n_1191), .b(n_4694), .o(g60345_p) );
in01f01 g60345_u1 ( .a(g60345_p), .o(n_4695) );
oa12f02 g60346_u0 ( .a(n_4080), .b(n_3289), .c(n_15856), .o(n_4693) );
no02f08 g60347_u0 ( .a(n_1353), .b(n_2874), .o(n_3170) );
no02f02 g60348_u0 ( .a(n_4856), .b(n_7031), .o(n_7032) );
no02f02 g60349_u0 ( .a(n_4857), .b(n_7031), .o(n_7030) );
no02f02 g60350_u0 ( .a(n_4858), .b(n_7031), .o(n_7029) );
ao12f02 g60353_u0 ( .a(n_3157), .b(n_2451), .c(wbm_rty_i), .o(n_2988) );
oa12f02 g60354_u0 ( .a(FE_OFN1083_n_13221), .b(n_4719), .c(FE_OCPN1839_n_1238), .o(n_7028) );
oa12f02 g60355_u0 ( .a(n_8451), .b(n_8450), .c(n_8540), .o(n_8520) );
oa12m02 g60356_u0 ( .a(n_8447), .b(n_8446), .c(n_8517), .o(n_8519) );
oa12f02 g60357_u0 ( .a(n_7789), .b(n_8468), .c(n_8517), .o(n_8470) );
oa12f02 g60358_u0 ( .a(n_8515), .b(n_8514), .c(n_8540), .o(n_8542) );
oa12f02 g60359_u0 ( .a(n_8513), .b(n_8512), .c(n_8540), .o(n_8541) );
oa12f02 g60360_u0 ( .a(n_7790), .b(n_8468), .c(n_8540), .o(n_8469) );
oa12f02 g60361_u0 ( .a(n_7788), .b(n_8465), .c(n_8517), .o(n_8467) );
oa12f02 g60362_u0 ( .a(n_7787), .b(n_8465), .c(n_8540), .o(n_8466) );
oa12f02 g60363_u0 ( .a(n_7786), .b(n_7785), .c(n_3280), .o(n_8464) );
oa12f02 g60364_u0 ( .a(n_8445), .b(n_8444), .c(n_8517), .o(n_8518) );
oa12f02 g60365_u0 ( .a(n_2135), .b(n_4816), .c(n_4853), .o(n_7027) );
ao12f10 g60398_u0 ( .a(n_2951), .b(n_3408), .c(FE_OFN191_n_1193), .o(n_4868) );
oa12f02 g60399_u0 ( .a(n_8449), .b(n_8540), .c(FE_OFN2086_n_8448), .o(n_8516) );
oa12f02 g60400_u0 ( .a(n_4211), .b(FE_OFN1183_n_3476), .c(wbm_sel_o_0_), .o(n_4867) );
oa12m02 g60401_u0 ( .a(n_4212), .b(FE_OFN1183_n_3476), .c(wbm_sel_o_1_), .o(n_4866) );
oa12m02 g60402_u0 ( .a(n_4213), .b(FE_OFN1181_n_3476), .c(wbm_sel_o_2_), .o(n_4864) );
oa12f02 g60403_u0 ( .a(n_4216), .b(FE_OFN1181_n_3476), .c(wbm_sel_o_3_), .o(n_4863) );
ao12f02 g60404_u0 ( .a(n_3376), .b(conf_wb_err_addr_in_965), .c(FE_OFN1143_n_15261), .o(n_4201) );
ao12f02 g60405_u0 ( .a(n_4504), .b(conf_wb_err_addr_in_968), .c(FE_OFN1145_n_15261), .o(n_4862) );
oa12f02 g60406_u0 ( .a(n_5758), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q), .c(n_15741), .o(n_7300) );
in01m01 g60407_u0 ( .a(n_7078), .o(g60407_sb) );
in01s01 TIMEBOOST_cell_67770 ( .a(TIMEBOOST_net_21196), .o(TIMEBOOST_net_21197) );
na03f02 TIMEBOOST_cell_47231 ( .a(FE_OFN1579_n_12306), .b(TIMEBOOST_net_13521), .c(FE_OFN1761_n_10780), .o(n_12653) );
na02f02 TIMEBOOST_cell_49708 ( .a(TIMEBOOST_net_15071), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_13185) );
na02m02 TIMEBOOST_cell_54714 ( .a(TIMEBOOST_net_17574), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_15401) );
in01f01 g60409_u0 ( .a(n_7078), .o(g60409_sb) );
na03f02 TIMEBOOST_cell_33292 ( .a(TIMEBOOST_net_582), .b(n_7321), .c(n_4897), .o(n_7322) );
na02f02 TIMEBOOST_cell_63333 ( .a(TIMEBOOST_net_20613), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_15374) );
na03m02 TIMEBOOST_cell_73017 ( .a(wbs_adr_i_0_), .b(g63582_sb), .c(g63582_db), .o(n_4106) );
oa12s02 g60410_u0 ( .a(n_4811), .b(n_4197), .c(FE_OFN1171_n_5592), .o(n_5718) );
oa12f01 g60411_u0 ( .a(n_7339), .b(n_3251), .c(n_7608), .o(n_7609) );
ao12f02 g60412_u0 ( .a(n_4198), .b(FE_OFN1612_n_2122), .c(wishbone_slave_unit_pcim_sm_data_in), .o(n_4692) );
ao12f02 g60413_u0 ( .a(n_3375), .b(conf_wb_err_addr_in_957), .c(FE_OFN1144_n_15261), .o(n_4200) );
no02f04 g60414_u0 ( .a(wbm_adr_o_21_), .b(n_2456), .o(g60414_p) );
ao12f02 g60414_u1 ( .a(g60414_p), .b(wbm_adr_o_21_), .c(n_2456), .o(n_2987) );
no02f06 g60415_u0 ( .a(conf_wb_err_addr_in_962), .b(n_2459), .o(g60415_p) );
ao12f02 g60415_u1 ( .a(g60415_p), .b(conf_wb_err_addr_in_962), .c(n_2459), .o(n_2986) );
in01f02 g60416_u0 ( .a(n_7019), .o(n_7298) );
ao22f02 g60417_u0 ( .a(n_7007), .b(n_14922), .c(FE_OFN1159_n_15325), .d(n_7241), .o(n_7019) );
in01f02 g60418_u0 ( .a(n_7018), .o(n_7297) );
ao22f02 g60419_u0 ( .a(n_7015), .b(n_14932), .c(FE_OFN1158_n_15325), .d(n_7295), .o(n_7018) );
in01m01 g60420_u0 ( .a(n_7812), .o(n_8463) );
ao22f01 g60421_u0 ( .a(n_7810), .b(configuration_interrupt_line), .c(n_7809), .d(n_7806), .o(n_7812) );
in01m02 g60422_u0 ( .a(n_7811), .o(n_8462) );
ao22f02 g60423_u0 ( .a(n_7810), .b(configuration_interrupt_line_37), .c(n_7809), .d(n_7802), .o(n_7811) );
in01m02 g60424_u0 ( .a(n_7808), .o(n_8461) );
ao22f02 g60425_u0 ( .a(n_7810), .b(configuration_interrupt_line_38), .c(n_7809), .d(n_7800), .o(n_7808) );
in01f02 g60426_u0 ( .a(n_7807), .o(n_8460) );
ao22f02 g60427_u0 ( .a(n_7804), .b(wbu_mrl_en_in_142), .c(n_7803), .d(n_7806), .o(n_7807) );
in01f02 g60428_u0 ( .a(n_7805), .o(n_8459) );
ao22f02 g60429_u0 ( .a(n_7804), .b(wbu_pref_en_in_137), .c(n_7803), .d(n_7802), .o(n_7805) );
in01f02 g60430_u0 ( .a(n_7801), .o(n_8458) );
ao22f02 g60431_u0 ( .a(n_7804), .b(n_14906), .c(n_7803), .d(n_7800), .o(n_7801) );
in01m02 g60432_u0 ( .a(n_7799), .o(n_8457) );
ao22f02 g60433_u0 ( .a(n_7810), .b(configuration_interrupt_line_42), .c(n_7792), .d(n_7809), .o(n_7799) );
in01f02 g60434_u0 ( .a(n_7296), .o(n_7470) );
ao22f02 g60435_u0 ( .a(n_7293), .b(pciu_am1_in_538), .c(n_16916), .d(n_7295), .o(n_7296) );
in01f01 g60436_u0 ( .a(n_7469), .o(n_7607) );
ao22f01 g60437_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in), .c(n_7466), .d(n_7289), .o(n_7469) );
in01f02 g60438_u0 ( .a(n_7468), .o(n_7606) );
ao22f02 g60439_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_243), .c(n_7466), .d(n_7231), .o(n_7468) );
in01f02 g60440_u0 ( .a(n_7465), .o(n_7605) );
ao22f02 g60441_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_244), .c(n_7466), .d(n_7282), .o(n_7465) );
in01f02 g60442_u0 ( .a(n_7294), .o(n_7464) );
ao22f02 g60443_u0 ( .a(n_7293), .b(pciu_am1_in_539), .c(n_16916), .d(n_7291), .o(n_7294) );
in01f01 g60444_u0 ( .a(n_7463), .o(n_7604) );
ao22f01 g60445_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_245), .c(n_7466), .d(n_7279), .o(n_7463) );
in01f02 g60446_u0 ( .a(n_7462), .o(n_7603) );
ao22f02 g60447_u0 ( .a(n_7420), .b(pciu_bar0_in_364), .c(n_15931), .d(n_7272), .o(n_7462) );
in01f01 g60448_u0 ( .a(n_7461), .o(n_7602) );
ao22f01 g60449_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_246), .c(n_7466), .d(n_7426), .o(n_7461) );
in01f02 g60450_u0 ( .a(n_7290), .o(n_7460) );
ao22f02 g60451_u0 ( .a(n_7283), .b(pciu_am1_in), .c(n_16916), .d(n_7289), .o(n_7290) );
in01f02 g60452_u0 ( .a(n_7459), .o(n_7601) );
ao22f02 g60453_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_247), .c(n_7466), .d(n_7424), .o(n_7459) );
in01f02 g60454_u0 ( .a(n_7288), .o(n_7458) );
ao22f02 g60455_u0 ( .a(n_7273), .b(pciu_am1_in_531), .c(n_16916), .d(n_7287), .o(n_7288) );
in01f02 g60456_u0 ( .a(n_7457), .o(n_7600) );
ao22f02 g60457_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_248), .c(n_7466), .d(n_7422), .o(n_7457) );
in01f02 g60458_u0 ( .a(n_7286), .o(n_7456) );
ao22f02 g60459_u0 ( .a(n_7293), .b(pciu_am1_in_535), .c(n_16916), .d(n_7285), .o(n_7286) );
in01f02 g60460_u0 ( .a(n_7455), .o(n_7599) );
ao22f02 g60461_u0 ( .a(n_7467), .b(wbu_latency_tim_val_in_249), .c(n_7466), .d(n_7440), .o(n_7455) );
in01f01 g60462_u0 ( .a(n_7454), .o(n_7598) );
ao22m01 g60463_u0 ( .a(n_7437), .b(configuration_cache_line_size_reg), .c(n_7466), .d(n_7806), .o(n_7454) );
in01f02 g60464_u0 ( .a(n_7284), .o(n_7453) );
ao22f02 g60465_u0 ( .a(n_7283), .b(pciu_am1_in_519), .c(n_16916), .d(n_7282), .o(n_7284) );
in01f02 g60466_u0 ( .a(n_7016), .o(n_7281) );
ao22f02 g60467_u0 ( .a(n_7015), .b(n_14930), .c(FE_OFN1158_n_15325), .d(n_7239), .o(n_7016) );
in01f02 g60468_u0 ( .a(n_7280), .o(n_7452) );
ao22f02 g60469_u0 ( .a(n_7283), .b(pciu_am1_in_520), .c(n_16916), .d(n_7279), .o(n_7280) );
in01f02 g60470_u0 ( .a(n_7278), .o(n_7451) );
ao22f02 g60471_u0 ( .a(n_7283), .b(pciu_am1_in_521), .c(n_16916), .d(n_7426), .o(n_7278) );
in01f02 g60472_u0 ( .a(n_7277), .o(n_7450) );
ao22f02 g60473_u0 ( .a(n_7283), .b(pciu_am1_in_522), .c(n_16916), .d(n_7424), .o(n_7277) );
in01f02 g60474_u0 ( .a(n_7276), .o(n_7449) );
ao22f02 g60475_u0 ( .a(n_7283), .b(pciu_am1_in_523), .c(n_16916), .d(n_7422), .o(n_7276) );
in01f02 g60476_u0 ( .a(n_7275), .o(n_7448) );
ao22f02 g60477_u0 ( .a(n_7283), .b(pciu_am1_in_524), .c(n_16916), .d(n_7440), .o(n_7275) );
in01f02 g60478_u0 ( .a(n_7274), .o(n_7447) );
ao22f02 g60479_u0 ( .a(n_7273), .b(pciu_am1_in_525), .c(n_16916), .d(n_7272), .o(n_7274) );
in01f02 g60480_u0 ( .a(n_7014), .o(n_7271) );
ao22f02 g60481_u0 ( .a(n_7012), .b(n_14913), .c(FE_OFN1159_n_15325), .d(n_7282), .o(n_7014) );
in01f02 g60482_u0 ( .a(n_7270), .o(n_7446) );
ao22f02 g60483_u0 ( .a(n_7273), .b(pciu_am1_in_526), .c(n_16916), .d(n_7269), .o(n_7270) );
in01f02 g60484_u0 ( .a(n_7268), .o(n_7445) );
ao22f02 g60485_u0 ( .a(n_7273), .b(pciu_am1_in_527), .c(n_16916), .d(n_7267), .o(n_7268) );
in01f02 g60486_u0 ( .a(n_7266), .o(n_7444) );
ao22f02 g60487_u0 ( .a(n_7273), .b(pciu_am1_in_529), .c(n_16916), .d(n_7265), .o(n_7266) );
in01f02 g60488_u0 ( .a(n_7013), .o(n_7264) );
ao22f02 g60489_u0 ( .a(n_7012), .b(n_14914), .c(FE_OFN1159_n_15325), .d(n_7279), .o(n_7013) );
in01f02 g60490_u0 ( .a(n_7011), .o(n_7263) );
ao22f02 g60491_u0 ( .a(n_7012), .b(n_14915), .c(FE_OFN1159_n_15325), .d(n_7426), .o(n_7011) );
in01f02 g60492_u0 ( .a(n_7010), .o(n_7262) );
ao22f02 g60493_u0 ( .a(n_7012), .b(n_14916), .c(FE_OFN1159_n_15325), .d(n_7424), .o(n_7010) );
in01f02 g60494_u0 ( .a(n_7009), .o(n_7261) );
ao22f02 g60495_u0 ( .a(n_7012), .b(n_14917), .c(FE_OFN1159_n_15325), .d(n_7422), .o(n_7009) );
in01f02 g60496_u0 ( .a(n_7260), .o(n_7443) );
ao22f02 g60497_u0 ( .a(n_7273), .b(pciu_am1_in_530), .c(n_16916), .d(n_7259), .o(n_7260) );
in01f02 g60498_u0 ( .a(n_7442), .o(n_7597) );
ao22f02 g60499_u0 ( .a(n_7427), .b(pciu_bar0_in_363), .c(n_15931), .d(n_7440), .o(n_7442) );
in01f02 g60500_u0 ( .a(n_7008), .o(n_7258) );
ao22f02 g60501_u0 ( .a(n_7007), .b(n_14919), .c(FE_OFN1159_n_15325), .d(n_7272), .o(n_7008) );
in01f02 g60502_u0 ( .a(n_7006), .o(n_7257) );
ao22f02 g60503_u0 ( .a(n_7007), .b(n_14920), .c(FE_OFN1159_n_15325), .d(n_7269), .o(n_7006) );
in01f02 g60504_u0 ( .a(n_7005), .o(n_7256) );
ao22f02 g60505_u0 ( .a(n_7007), .b(n_14921), .c(FE_OFN1159_n_15325), .d(n_7267), .o(n_7005) );
in01f02 g60506_u0 ( .a(n_7255), .o(n_7439) );
ao22f02 g60507_u0 ( .a(n_7273), .b(pciu_am1_in_532), .c(n_16916), .d(n_7254), .o(n_7255) );
in01f02 g60508_u0 ( .a(n_7004), .o(n_7253) );
ao22f02 g60509_u0 ( .a(n_7007), .b(n_14923), .c(FE_OFN1159_n_15325), .d(n_7265), .o(n_7004) );
in01f02 g60510_u0 ( .a(n_7003), .o(n_7252) );
ao22f02 g60511_u0 ( .a(n_7007), .b(n_14924), .c(FE_OFN1159_n_15325), .d(n_7259), .o(n_7003) );
in01f02 g60512_u0 ( .a(n_7002), .o(n_7251) );
ao22f02 g60513_u0 ( .a(n_7007), .b(n_14925), .c(FE_OFN1158_n_15325), .d(n_7287), .o(n_7002) );
in01f01 g60514_u0 ( .a(n_7438), .o(n_7596) );
ao22f01 g60515_u0 ( .a(n_7437), .b(configuration_cache_line_size_reg_2996), .c(n_7466), .d(n_7802), .o(n_7438) );
in01f02 g60516_u0 ( .a(n_7250), .o(n_7436) );
ao22f02 g60517_u0 ( .a(n_7293), .b(pciu_am1_in_533), .c(n_16916), .d(n_7249), .o(n_7250) );
in01f02 g60518_u0 ( .a(n_7001), .o(n_7248) );
ao22f02 g60519_u0 ( .a(n_7007), .b(n_14926), .c(FE_OFN1158_n_15325), .d(n_7254), .o(n_7001) );
in01f02 g60520_u0 ( .a(n_7000), .o(n_7247) );
ao22f02 g60521_u0 ( .a(n_7015), .b(n_14927), .c(FE_OFN1158_n_15325), .d(n_7249), .o(n_7000) );
in01f01 g60522_u0 ( .a(n_6999), .o(n_7246) );
ao22f01 g60523_u0 ( .a(n_7015), .b(n_14928), .c(FE_OFN1158_n_15325), .d(n_7244), .o(n_6999) );
in01f02 g60524_u0 ( .a(n_7245), .o(n_7435) );
ao22f02 g60525_u0 ( .a(n_7293), .b(pciu_am1_in_534), .c(n_16916), .d(n_7244), .o(n_7245) );
in01f02 g60526_u0 ( .a(n_6998), .o(n_7243) );
ao22f02 g60527_u0 ( .a(n_7015), .b(n_14929), .c(FE_OFN1158_n_15325), .d(n_7285), .o(n_6998) );
in01f01 g60528_u0 ( .a(n_7434), .o(n_7595) );
ao22f01 g60529_u0 ( .a(n_7437), .b(wbu_cache_line_size_in_206), .c(n_7466), .d(n_7800), .o(n_7434) );
in01f02 g60530_u0 ( .a(n_7242), .o(n_7433) );
ao22f02 g60531_u0 ( .a(n_7273), .b(pciu_am1_in_528), .c(n_16916), .d(n_7241), .o(n_7242) );
in01f02 g60532_u0 ( .a(n_7240), .o(n_7432) );
ao22f02 g60533_u0 ( .a(n_7293), .b(pciu_am1_in_536), .c(n_16916), .d(n_7239), .o(n_7240) );
in01f02 g60534_u0 ( .a(n_6997), .o(n_7238) );
ao22f02 g60535_u0 ( .a(n_7015), .b(n_14934), .c(FE_OFN1158_n_15325), .d(n_6996), .o(n_6997) );
in01f02 g60536_u0 ( .a(n_6995), .o(n_7237) );
ao22f02 g60537_u0 ( .a(n_7012), .b(n_14911), .c(FE_OFN1159_n_15325), .d(n_7289), .o(n_6995) );
in01f02 g60538_u0 ( .a(n_6994), .o(n_7236) );
ao22f02 g60539_u0 ( .a(n_7012), .b(n_14912), .c(FE_OFN1159_n_15325), .d(n_7231), .o(n_6994) );
in01f02 g60540_u0 ( .a(n_7235), .o(n_7431) );
ao22f02 g60541_u0 ( .a(n_7293), .b(pciu_am1_in_537), .c(n_16916), .d(n_7234), .o(n_7235) );
in01s01 TIMEBOOST_cell_63605 ( .a(TIMEBOOST_net_20785), .o(TIMEBOOST_net_20784) );
in01f02 g60543_u0 ( .a(n_7233), .o(n_7430) );
ao22f02 g60544_u0 ( .a(n_7293), .b(pciu_am1_in_540), .c(n_16916), .d(n_6996), .o(n_7233) );
in01f02 g60545_u0 ( .a(n_7232), .o(n_7429) );
ao22f02 g60546_u0 ( .a(n_7283), .b(pciu_am1_in_518), .c(n_16916), .d(n_7231), .o(n_7232) );
in01f02 g60547_u0 ( .a(n_7428), .o(n_7594) );
ao22f02 g60548_u0 ( .a(n_7427), .b(pciu_bar0_in), .c(n_15931), .d(n_7426), .o(n_7428) );
in01f02 g60549_u0 ( .a(n_7425), .o(n_7593) );
ao22f02 g60550_u0 ( .a(n_7427), .b(pciu_bar0_in_361), .c(n_15931), .d(n_7424), .o(n_7425) );
in01f02 g60551_u0 ( .a(n_7423), .o(n_7592) );
ao22f02 g60552_u0 ( .a(n_7427), .b(pciu_bar0_in_362), .c(n_15931), .d(n_7422), .o(n_7423) );
in01f02 g60553_u0 ( .a(n_7421), .o(n_7591) );
ao22f02 g60554_u0 ( .a(n_7420), .b(pciu_bar0_in_366), .c(n_15931), .d(n_7267), .o(n_7421) );
in01f01 g60555_u0 ( .a(n_7419), .o(n_7590) );
ao22f01 g60556_u0 ( .a(n_7437), .b(wbu_cache_line_size_in_210), .c(n_7792), .d(n_7466), .o(n_7419) );
no02s02 g60557_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_7_), .b(n_2295), .o(g60557_p) );
ao12s02 g60557_u1 ( .a(g60557_p), .b(pci_target_unit_del_sync_comp_cycle_count_7_), .c(n_2295), .o(n_2304) );
in01f02 g60558_u0 ( .a(n_7418), .o(n_7589) );
ao22f02 g60559_u0 ( .a(n_7420), .b(pciu_bar0_in_365), .c(n_15931), .d(n_7269), .o(n_7418) );
in01f02 g60560_u0 ( .a(n_7417), .o(n_7588) );
ao22f02 g60561_u0 ( .a(n_7420), .b(pciu_bar0_in_367), .c(n_15931), .d(n_7241), .o(n_7417) );
in01f02 g60562_u0 ( .a(n_7416), .o(n_7587) );
ao22f02 g60563_u0 ( .a(n_7420), .b(pciu_bar0_in_368), .c(n_15931), .d(n_7265), .o(n_7416) );
in01f02 g60564_u0 ( .a(n_7415), .o(n_7586) );
ao22f02 g60565_u0 ( .a(n_7420), .b(pciu_bar0_in_369), .c(n_15931), .d(n_7259), .o(n_7415) );
in01f02 g60566_u0 ( .a(n_7414), .o(n_7585) );
ao22f02 g60567_u0 ( .a(n_7420), .b(pciu_bar0_in_370), .c(n_15931), .d(n_7287), .o(n_7414) );
in01f02 g60568_u0 ( .a(n_7413), .o(n_7584) );
ao22f02 g60569_u0 ( .a(n_7420), .b(pciu_bar0_in_371), .c(n_15931), .d(n_7254), .o(n_7413) );
in01f02 g60570_u0 ( .a(n_7412), .o(n_7583) );
ao22f02 g60571_u0 ( .a(n_7410), .b(pciu_bar0_in_372), .c(n_15931), .d(n_7249), .o(n_7412) );
in01f02 g60572_u0 ( .a(n_7411), .o(n_7582) );
ao22f02 g60573_u0 ( .a(n_7410), .b(pciu_bar0_in_373), .c(n_15931), .d(n_7244), .o(n_7411) );
in01f02 g60574_u0 ( .a(n_7798), .o(n_8456) );
ao22f06 g60575_u0 ( .a(n_7796), .b(configuration_sync_command_bit0), .c(n_7795), .d(n_7806), .o(n_7798) );
in01f02 g60576_u0 ( .a(n_7409), .o(n_7581) );
ao22f02 g60577_u0 ( .a(n_7410), .b(pciu_bar0_in_374), .c(n_15931), .d(n_7285), .o(n_7409) );
in01f02 g60578_u0 ( .a(n_7408), .o(n_7580) );
ao22f02 g60579_u0 ( .a(n_7410), .b(pciu_bar0_in_375), .c(n_15931), .d(n_7239), .o(n_7408) );
in01f02 g60580_u0 ( .a(n_7407), .o(n_7579) );
ao22f02 g60581_u0 ( .a(n_7410), .b(pciu_bar0_in_376), .c(n_15931), .d(n_7234), .o(n_7407) );
in01f02 g60582_u0 ( .a(n_7406), .o(n_7578) );
ao22f02 g60583_u0 ( .a(n_7410), .b(pciu_bar0_in_377), .c(n_15931), .d(n_7295), .o(n_7406) );
in01f02 g60584_u0 ( .a(n_7405), .o(n_7577) );
ao22f02 g60585_u0 ( .a(n_7410), .b(pciu_bar0_in_378), .c(n_15931), .d(n_7291), .o(n_7405) );
na02f08 TIMEBOOST_cell_18464 ( .a(TIMEBOOST_net_5595), .b(n_16967), .o(n_13807) );
in01f02 g60587_u0 ( .a(n_7797), .o(n_8455) );
ao22f02 g60588_u0 ( .a(n_7796), .b(configuration_sync_command_bit1), .c(n_7795), .d(n_7802), .o(n_7797) );
in01f02 g60589_u0 ( .a(n_7404), .o(n_7576) );
ao22f02 g60590_u0 ( .a(n_7410), .b(pciu_bar0_in_379), .c(n_15931), .d(n_6996), .o(n_7404) );
no02m02 g60591_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .b(n_2275), .o(g60591_p) );
ao12m01 g60591_u1 ( .a(g60591_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .c(n_2275), .o(n_2302) );
in01f01 g60592_u0 ( .a(n_7794), .o(n_8454) );
ao22f01 g60593_u0 ( .a(n_7796), .b(configuration_command_bit), .c(n_7795), .d(n_7800), .o(n_7794) );
in01f02 g60595_u0 ( .a(n_7793), .o(n_8453) );
ao22f02 g60596_u0 ( .a(n_7796), .b(configuration_sync_command_bit6), .c(n_7795), .d(n_7792), .o(n_7793) );
in01f02 g60597_u0 ( .a(n_6993), .o(n_7229) );
ao22f02 g60598_u0 ( .a(n_7015), .b(n_14931), .c(FE_OFN1158_n_15325), .d(n_7234), .o(n_6993) );
in01f02 g60599_u0 ( .a(n_6992), .o(n_7228) );
ao22f02 g60600_u0 ( .a(n_7012), .b(n_14918), .c(FE_OFN1159_n_15325), .d(n_7440), .o(n_6992) );
in01f02 g60601_u0 ( .a(n_6991), .o(n_7227) );
ao22f02 g60602_u0 ( .a(n_7015), .b(n_14933), .c(FE_OFN1158_n_15325), .d(n_7291), .o(n_6991) );
in01f01 g60603_u0 ( .a(n_6986), .o(g60603_sb) );
na02f02 g60603_u1 ( .a(wbu_latency_tim_val_in_248), .b(g60603_sb), .o(g60603_da) );
in01f01 g60604_u0 ( .a(FE_OFN1183_n_3476), .o(g60604_sb) );
na02f08 TIMEBOOST_cell_3251 ( .a(TIMEBOOST_net_185), .b(n_2993), .o(n_3353) );
na02m10 TIMEBOOST_cell_53003 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q), .b(wishbone_slave_unit_pcim_sm_data_in_662), .o(TIMEBOOST_net_16719) );
na02s01 TIMEBOOST_cell_3252 ( .a(n_2648), .b(n_8511), .o(TIMEBOOST_net_186) );
in01f01 g60605_u0 ( .a(FE_OFN1179_n_3476), .o(g60605_sb) );
na02s06 TIMEBOOST_cell_52181 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q), .o(TIMEBOOST_net_16308) );
na02m02 TIMEBOOST_cell_69488 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q), .o(TIMEBOOST_net_21952) );
na02s01 TIMEBOOST_cell_54179 ( .a(configuration_wb_err_addr_561), .b(conf_wb_err_addr_in_970), .o(TIMEBOOST_net_17307) );
in01m01 g60606_u0 ( .a(FE_OFN1185_n_3476), .o(g60606_sb) );
na02m04 TIMEBOOST_cell_37182 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q), .o(TIMEBOOST_net_10203) );
na02f02 TIMEBOOST_cell_53085 ( .a(n_3978), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q), .o(TIMEBOOST_net_16760) );
na03m02 TIMEBOOST_cell_73574 ( .a(TIMEBOOST_net_17388), .b(FE_OFN1219_n_6886), .c(g62466_sb), .o(n_6662) );
in01f01 g60607_u0 ( .a(FE_OFN1185_n_3476), .o(g60607_sb) );
na04m02 TIMEBOOST_cell_64951 ( .a(n_3741), .b(n_65), .c(g64949_sb), .d(FE_OFN647_n_4497), .o(n_3667) );
na03f02 TIMEBOOST_cell_66449 ( .a(TIMEBOOST_net_17113), .b(FE_OFN1310_n_6624), .c(g62439_sb), .o(n_6718) );
in01f02 g60608_u0 ( .a(FE_OFN1185_n_3476), .o(g60608_sb) );
na03m02 TIMEBOOST_cell_72701 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q), .b(g63570_sb), .c(g63570_db), .o(n_4592) );
in01f02 g60609_u0 ( .a(FE_OFN1179_n_3476), .o(g60609_sb) );
na02m04 TIMEBOOST_cell_69610 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_22013) );
na02m01 TIMEBOOST_cell_37184 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q), .o(TIMEBOOST_net_10204) );
na02m01 TIMEBOOST_cell_37185 ( .a(TIMEBOOST_net_10204), .b(n_4730), .o(TIMEBOOST_net_176) );
in01f02 g60610_u0 ( .a(FE_OFN1185_n_3476), .o(g60610_sb) );
na02m10 TIMEBOOST_cell_28015 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_8112) );
na02s01 TIMEBOOST_cell_47525 ( .a(pci_target_unit_del_sync_comp_rty_exp_clr), .b(pci_target_unit_wbm_sm_pci_tar_read_request), .o(TIMEBOOST_net_13980) );
na02f10 TIMEBOOST_cell_47549 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_4_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .o(TIMEBOOST_net_13992) );
in01m01 g60611_u0 ( .a(FE_OFN1185_n_3476), .o(g60611_sb) );
na03s02 TIMEBOOST_cell_46227 ( .a(TIMEBOOST_net_12417), .b(FE_OFN250_n_9789), .c(TIMEBOOST_net_10562), .o(TIMEBOOST_net_9487) );
na02s08 TIMEBOOST_cell_47551 ( .a(wbs_dat_i_7_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q), .o(TIMEBOOST_net_13993) );
in01f02 g60612_u0 ( .a(FE_OFN1185_n_3476), .o(g60612_sb) );
na03f02 TIMEBOOST_cell_73379 ( .a(TIMEBOOST_net_16697), .b(FE_OFN1301_n_5763), .c(g62049_sb), .o(n_7761) );
na02s02 TIMEBOOST_cell_54104 ( .a(TIMEBOOST_net_17269), .b(g57969_sb), .o(TIMEBOOST_net_14639) );
na02f02 TIMEBOOST_cell_39555 ( .a(TIMEBOOST_net_11389), .b(g62847_sb), .o(n_5277) );
in01f02 g60613_u0 ( .a(FE_OFN1185_n_3476), .o(g60613_sb) );
na03f02 TIMEBOOST_cell_71158 ( .a(TIMEBOOST_net_15573), .b(wishbone_slave_unit_del_sync_addr_out_reg_6__Q), .c(n_13221), .o(TIMEBOOST_net_22787) );
in01f02 g60614_u0 ( .a(FE_OFN1179_n_3476), .o(g60614_sb) );
in01f01 g60615_u0 ( .a(FE_OFN1183_n_3476), .o(g60615_sb) );
na02s01 TIMEBOOST_cell_3253 ( .a(TIMEBOOST_net_186), .b(n_3021), .o(n_3377) );
na02s02 TIMEBOOST_cell_68193 ( .a(TIMEBOOST_net_21304), .b(g65907_sb), .o(n_2174) );
in01f02 g60616_u0 ( .a(FE_OFN1185_n_3476), .o(g60616_sb) );
na02f08 TIMEBOOST_cell_37111 ( .a(TIMEBOOST_net_10167), .b(n_15981), .o(n_15982) );
in01f02 g60617_u0 ( .a(FE_OFN1184_n_3476), .o(g60617_sb) );
na02m02 TIMEBOOST_cell_25845 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q), .b(g64290_sb), .o(TIMEBOOST_net_7027) );
na03f02 TIMEBOOST_cell_66069 ( .a(n_3524), .b(g63553_sb), .c(TIMEBOOST_net_7660), .o(n_4924) );
na04f04 TIMEBOOST_cell_24647 ( .a(n_9081), .b(g57239_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q), .d(FE_OFN2167_n_8567), .o(n_10428) );
in01f01 g60618_u0 ( .a(FE_OFN1179_n_3476), .o(g60618_sb) );
na02s06 TIMEBOOST_cell_47571 ( .a(wbs_dat_i_2_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q), .o(TIMEBOOST_net_14003) );
na02m10 TIMEBOOST_cell_49541 ( .a(g53892_sb), .b(wishbone_slave_unit_pcim_if_wbw_cbe_in_416), .o(TIMEBOOST_net_14988) );
in01f01 g60619_u0 ( .a(FE_OFN1179_n_3476), .o(g60619_sb) );
in01m01 g60620_u0 ( .a(FE_OFN1180_n_3476), .o(g60620_sb) );
in01f02 g60621_u0 ( .a(FE_OFN1181_n_3476), .o(g60621_sb) );
na02m08 TIMEBOOST_cell_37186 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q), .b(pci_target_unit_fifos_pciw_control_in_157), .o(TIMEBOOST_net_10205) );
na02f02 TIMEBOOST_cell_71079 ( .a(TIMEBOOST_net_22747), .b(g62935_sb), .o(n_6011) );
na03m02 TIMEBOOST_cell_72597 ( .a(TIMEBOOST_net_23152), .b(FE_OFN1642_n_4671), .c(TIMEBOOST_net_21689), .o(TIMEBOOST_net_17033) );
in01f02 g60622_u0 ( .a(FE_OFN1180_n_3476), .o(g60622_sb) );
na02s01 TIMEBOOST_cell_40364 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_), .o(TIMEBOOST_net_11794) );
na02s02 TIMEBOOST_cell_49280 ( .a(TIMEBOOST_net_14857), .b(TIMEBOOST_net_10856), .o(TIMEBOOST_net_9543) );
na02s02 TIMEBOOST_cell_48259 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q), .o(TIMEBOOST_net_14347) );
in01m01 g60623_u0 ( .a(FE_OFN1180_n_3476), .o(g60623_sb) );
na03f02 TIMEBOOST_cell_73505 ( .a(TIMEBOOST_net_22586), .b(g52447_sb), .c(TIMEBOOST_net_22854), .o(n_14845) );
na03f02 TIMEBOOST_cell_73380 ( .a(TIMEBOOST_net_16692), .b(FE_OFN1299_n_5763), .c(g62036_sb), .o(n_7780) );
in01f02 g60624_u0 ( .a(FE_OFN1181_n_3476), .o(g60624_sb) );
na02m08 TIMEBOOST_cell_52199 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_127), .o(TIMEBOOST_net_16317) );
na02f06 TIMEBOOST_cell_52467 ( .a(g58375_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q), .o(TIMEBOOST_net_16451) );
in01f02 g60625_u0 ( .a(FE_OFN1181_n_3476), .o(g60625_sb) );
in01m08 TIMEBOOST_cell_35518 ( .a(conf_wb_err_addr_in_950), .o(TIMEBOOST_net_10109) );
na03f02 TIMEBOOST_cell_25014 ( .a(FE_RN_137_0), .b(n_10907), .c(n_12570), .o(n_12832) );
na02f01 g63091_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q), .b(FE_OFN1104_g64577_p), .o(g63091_db) );
in01m01 g60626_u0 ( .a(FE_OFN1182_n_3476), .o(g60626_sb) );
na02m01 g63089_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q), .b(FE_OFN1104_g64577_p), .o(g63089_db) );
in01s01 TIMEBOOST_cell_64266 ( .a(pci_target_unit_fifos_pcir_data_in_171), .o(TIMEBOOST_net_21122) );
in01m01 g60627_u0 ( .a(FE_OFN1181_n_3476), .o(g60627_sb) );
na03f02 TIMEBOOST_cell_34855 ( .a(TIMEBOOST_net_9321), .b(FE_OFN1368_n_8567), .c(g57289_sb), .o(n_11463) );
na02s01 TIMEBOOST_cell_45441 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q), .o(TIMEBOOST_net_13615) );
na02m01 g63056_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q), .b(FE_OFN1104_g64577_p), .o(g63056_db) );
in01f02 g60628_u0 ( .a(FE_OFN1181_n_3476), .o(g60628_sb) );
na02f02 TIMEBOOST_cell_30467 ( .a(n_9456), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q), .o(TIMEBOOST_net_9338) );
na02m01 g63052_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q), .b(FE_OFN1104_g64577_p), .o(g63052_db) );
na03f02 TIMEBOOST_cell_25016 ( .a(FE_RN_227_0), .b(n_11730), .c(n_12568), .o(n_12830) );
in01f02 g60629_u0 ( .a(FE_OFN1182_n_3476), .o(g60629_sb) );
na03m06 TIMEBOOST_cell_69074 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q), .b(FE_OFN1012_n_4734), .c(TIMEBOOST_net_17235), .o(TIMEBOOST_net_21745) );
na02m02 TIMEBOOST_cell_69013 ( .a(TIMEBOOST_net_21714), .b(g65378_sb), .o(TIMEBOOST_net_12548) );
in01m01 g60630_u0 ( .a(FE_OFN1180_n_3476), .o(g60630_sb) );
in01m06 TIMEBOOST_cell_35519 ( .a(TIMEBOOST_net_10109), .o(TIMEBOOST_net_10110) );
na03f02 TIMEBOOST_cell_25018 ( .a(n_10974), .b(FE_RN_35_0), .c(n_12584), .o(n_12846) );
na02m01 g63013_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q), .b(FE_OFN1104_g64577_p), .o(g63013_db) );
in01f02 g60631_u0 ( .a(FE_OFN1180_n_3476), .o(g60631_sb) );
na04s02 TIMEBOOST_cell_67969 ( .a(TIMEBOOST_net_12469), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q), .c(FE_OFN560_n_9895), .d(g57931_sb), .o(TIMEBOOST_net_9408) );
na03f02 TIMEBOOST_cell_25020 ( .a(FE_RN_185_0), .b(n_10895), .c(n_12567), .o(n_12829) );
na02f01 g62852_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q), .b(FE_OFN1104_g64577_p), .o(g62852_db) );
in01f01 g60632_u0 ( .a(FE_OFN1186_n_3476), .o(g60632_sb) );
na03f02 TIMEBOOST_cell_72952 ( .a(pci_target_unit_del_sync_addr_in_218), .b(g65214_sb), .c(TIMEBOOST_net_7159), .o(n_2673) );
na02f01 g62843_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q), .b(FE_OFN1104_g64577_p), .o(g62843_db) );
na02m02 g62833_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q), .b(FE_OFN1104_g64577_p), .o(g62833_db) );
in01f01 g60633_u0 ( .a(FE_OFN1179_n_3476), .o(g60633_sb) );
in01s01 TIMEBOOST_cell_35520 ( .a(TIMEBOOST_net_10111), .o(TIMEBOOST_net_10076) );
na02f01 g62811_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q), .b(FE_OFN1104_g64577_p), .o(g62811_db) );
na03f02 TIMEBOOST_cell_25022 ( .a(n_11717), .b(FE_RN_101_0), .c(n_12561), .o(n_12823) );
in01m01 g60634_u0 ( .a(FE_OFN1179_n_3476), .o(g60634_sb) );
in01s01 TIMEBOOST_cell_35521 ( .a(TIMEBOOST_net_10112), .o(TIMEBOOST_net_10111) );
na02f01 g62803_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN1104_g64577_p), .o(g62803_db) );
na03f02 TIMEBOOST_cell_25024 ( .a(n_10918), .b(FE_RN_197_0), .c(n_12572), .o(n_12834) );
in01m01 g60635_u0 ( .a(FE_OFN1179_n_3476), .o(g60635_sb) );
na02s01 TIMEBOOST_cell_53043 ( .a(wbm_adr_o_24_), .b(configuration_pci_err_addr_494), .o(TIMEBOOST_net_16739) );
na02m02 TIMEBOOST_cell_47672 ( .a(TIMEBOOST_net_14053), .b(g65957_db), .o(n_2165) );
in01f01 g60636_u0 ( .a(FE_OFN1183_n_3476), .o(g60636_sb) );
na02f08 TIMEBOOST_cell_3255 ( .a(n_1692), .b(TIMEBOOST_net_187), .o(n_2179) );
na02s02 TIMEBOOST_cell_48844 ( .a(TIMEBOOST_net_14639), .b(TIMEBOOST_net_12907), .o(TIMEBOOST_net_9367) );
na03m02 TIMEBOOST_cell_70368 ( .a(FE_OFN2021_n_4778), .b(TIMEBOOST_net_16654), .c(TIMEBOOST_net_632), .o(TIMEBOOST_net_22392) );
in01f02 g60637_u0 ( .a(FE_OFN1183_n_3476), .o(g60637_sb) );
na02m02 TIMEBOOST_cell_31745 ( .a(n_826), .b(TIMEBOOST_net_683), .o(TIMEBOOST_net_9977) );
na02s02 TIMEBOOST_cell_43144 ( .a(TIMEBOOST_net_12466), .b(g58103_sb), .o(n_9693) );
in01m01 g60638_u0 ( .a(FE_OFN1183_n_3476), .o(g60638_sb) );
na03f10 TIMEBOOST_cell_20892 ( .a(n_16504), .b(n_168), .c(n_16474), .o(n_15117) );
na02f02 TIMEBOOST_cell_28951 ( .a(n_14674), .b(n_14839), .o(TIMEBOOST_net_8580) );
na04f04 TIMEBOOST_cell_67918 ( .a(TIMEBOOST_net_11033), .b(FE_OFN1150_n_13249), .c(TIMEBOOST_net_20885), .d(g54146_sb), .o(n_13663) );
in01m01 g60639_u0 ( .a(FE_OFN1183_n_3476), .o(g60639_sb) );
na02f02 TIMEBOOST_cell_54490 ( .a(TIMEBOOST_net_17462), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_15410) );
in01m01 g60640_u0 ( .a(FE_OFN1182_n_3476), .o(g60640_sb) );
na02f01 g61958_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q), .b(FE_OFN1094_g64577_p), .o(g61958_db) );
in01f02 g60641_u0 ( .a(FE_OFN1179_n_3476), .o(g60641_sb) );
na02m01 TIMEBOOST_cell_37188 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q), .o(TIMEBOOST_net_10206) );
na04f04 TIMEBOOST_cell_24844 ( .a(wbs_dat_o_30_), .b(g52526_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_129), .d(FE_OFN2243_g52675_p), .o(n_13794) );
na02f02 TIMEBOOST_cell_71169 ( .a(TIMEBOOST_net_22792), .b(g54201_sb), .o(n_13418) );
in01f02 g60642_u0 ( .a(FE_OFN1185_n_3476), .o(g60642_sb) );
na02s01 TIMEBOOST_cell_48398 ( .a(TIMEBOOST_net_14416), .b(FE_OFN1794_n_9904), .o(TIMEBOOST_net_12694) );
na02m02 TIMEBOOST_cell_68448 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q), .b(FE_OFN671_n_4505), .o(TIMEBOOST_net_21432) );
na02s02 TIMEBOOST_cell_48209 ( .a(FE_OFN223_n_9844), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q), .o(TIMEBOOST_net_14322) );
in01f02 g60643_u0 ( .a(FE_OFN1185_n_3476), .o(g60643_sb) );
na03s01 TIMEBOOST_cell_46713 ( .a(TIMEBOOST_net_12816), .b(g58030_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q), .o(TIMEBOOST_net_9395) );
in01s01 TIMEBOOST_cell_67786 ( .a(TIMEBOOST_net_21213), .o(TIMEBOOST_net_21212) );
in01f02 g60644_u0 ( .a(FE_OFN1185_n_3476), .o(g60644_sb) );
no04f08 TIMEBOOST_cell_20893 ( .a(FE_RN_338_0), .b(FE_RN_348_0), .c(FE_RN_353_0), .d(FE_RN_343_0), .o(FE_RN_354_0) );
na02f02 g64253_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q), .b(g64253_sb), .o(g64253_da) );
in01f02 g60645_u0 ( .a(FE_OFN1185_n_3476), .o(g60645_sb) );
in01s01 TIMEBOOST_cell_35522 ( .a(TIMEBOOST_net_10113), .o(TIMEBOOST_net_10078) );
in01s01 TIMEBOOST_cell_67758 ( .a(TIMEBOOST_net_21184), .o(TIMEBOOST_net_21185) );
in01f02 g60646_u0 ( .a(FE_OFN1179_n_3476), .o(g60646_sb) );
in01s01 TIMEBOOST_cell_35523 ( .a(TIMEBOOST_net_10114), .o(TIMEBOOST_net_10113) );
na02m02 TIMEBOOST_cell_69487 ( .a(TIMEBOOST_net_21951), .b(g65732_sb), .o(n_1935) );
na04f04 TIMEBOOST_cell_73053 ( .a(n_2059), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q), .c(FE_OFN717_n_8176), .d(g62001_sb), .o(n_7893) );
in01f02 g60647_u0 ( .a(FE_OFN1185_n_3476), .o(g60647_sb) );
na03f02 TIMEBOOST_cell_70750 ( .a(n_2580), .b(n_2172), .c(n_2377), .o(TIMEBOOST_net_22583) );
na02f01 g61840_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN1094_g64577_p), .o(g61840_db) );
na02s01 TIMEBOOST_cell_48441 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_14438) );
in01f02 g60648_u0 ( .a(FE_OFN1184_n_3476), .o(g60648_sb) );
na04m02 TIMEBOOST_cell_67385 ( .a(n_3744), .b(g64944_sb), .c(g64944_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q), .o(TIMEBOOST_net_17574) );
na02s02 TIMEBOOST_cell_48521 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q), .b(g65910_sb), .o(TIMEBOOST_net_14478) );
na02f01 g63569_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q), .b(g63569_sb), .o(g63569_da) );
in01f02 g60649_u0 ( .a(FE_OFN1185_n_3476), .o(g60649_sb) );
na03m02 TIMEBOOST_cell_71846 ( .a(g65069_sb), .b(g65069_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q), .o(TIMEBOOST_net_23131) );
na03m02 TIMEBOOST_cell_64721 ( .a(FE_OFN662_n_4392), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q), .c(n_3761), .o(TIMEBOOST_net_14282) );
na02s02 TIMEBOOST_cell_50000 ( .a(TIMEBOOST_net_15217), .b(g58104_sb), .o(TIMEBOOST_net_9441) );
in01m01 g60650_u0 ( .a(FE_OFN1185_n_3476), .o(g60650_sb) );
na02m10 TIMEBOOST_cell_45241 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q), .o(TIMEBOOST_net_13515) );
na03f02 TIMEBOOST_cell_73777 ( .a(TIMEBOOST_net_8110), .b(n_13987), .c(FE_OFN1589_n_13736), .o(n_16259) );
no02f04 TIMEBOOST_cell_63424 ( .a(TIMEBOOST_net_7528), .b(FE_RN_371_0), .o(TIMEBOOST_net_20659) );
in01f01 g60651_u0 ( .a(FE_OFN1183_n_3476), .o(g60651_sb) );
na02f10 TIMEBOOST_cell_3257 ( .a(TIMEBOOST_net_188), .b(n_1694), .o(n_2175) );
in01s01 TIMEBOOST_cell_35524 ( .a(TIMEBOOST_net_10115), .o(TIMEBOOST_net_10082) );
no02f10 TIMEBOOST_cell_3258 ( .a(wishbone_slave_unit_pcim_if_del_req_in), .b(wishbone_slave_unit_pci_initiator_if_err_recovery), .o(TIMEBOOST_net_189) );
in01f02 g60652_u0 ( .a(FE_OFN1185_n_3476), .o(g60652_sb) );
na02s01 TIMEBOOST_cell_48851 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q), .o(TIMEBOOST_net_14643) );
na03f02 TIMEBOOST_cell_66451 ( .a(TIMEBOOST_net_17058), .b(n_6645), .c(g62472_sb), .o(n_6647) );
na03f02 TIMEBOOST_cell_66074 ( .a(TIMEBOOST_net_20910), .b(n_2559), .c(TIMEBOOST_net_668), .o(n_4892) );
in01f02 g60653_u0 ( .a(FE_OFN1184_n_3476), .o(g60653_sb) );
in01s01 TIMEBOOST_cell_35525 ( .a(TIMEBOOST_net_10116), .o(TIMEBOOST_net_10115) );
na02s01 TIMEBOOST_cell_48741 ( .a(g61810_sb), .b(g61810_db), .o(TIMEBOOST_net_14588) );
in01m01 g60654_u0 ( .a(FE_OFN1180_n_3476), .o(g60654_sb) );
na03f02 TIMEBOOST_cell_73054 ( .a(TIMEBOOST_net_22029), .b(FE_OFN2084_n_8407), .c(g61720_sb), .o(n_8384) );
na03f02 TIMEBOOST_cell_25086 ( .a(n_11823), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q), .c(n_12068), .o(n_12489) );
na02m04 TIMEBOOST_cell_62444 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_142), .o(TIMEBOOST_net_20169) );
in01m01 g60655_u0 ( .a(FE_OFN1185_n_3476), .o(g60655_sb) );
na02m02 TIMEBOOST_cell_63391 ( .a(TIMEBOOST_net_20642), .b(TIMEBOOST_net_13350), .o(TIMEBOOST_net_9350) );
na03f02 TIMEBOOST_cell_65168 ( .a(TIMEBOOST_net_20318), .b(g64180_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q), .o(TIMEBOOST_net_15065) );
na02s02 TIMEBOOST_cell_38414 ( .a(FE_OFN215_n_9856), .b(g57952_sb), .o(TIMEBOOST_net_10819) );
in01m01 g60656_u0 ( .a(FE_OFN1181_n_3476), .o(g60656_sb) );
na02s02 TIMEBOOST_cell_68276 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q), .b(g65891_sb), .o(TIMEBOOST_net_21346) );
in01s01 TIMEBOOST_cell_67767 ( .a(pci_target_unit_fifos_pcir_data_in_181), .o(TIMEBOOST_net_21194) );
na04f04 TIMEBOOST_cell_24662 ( .a(n_9748), .b(g57175_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q), .d(FE_OFN2180_n_8567), .o(n_11580) );
in01m01 g60657_u0 ( .a(FE_OFN1180_n_3476), .o(g60657_sb) );
na03f02 TIMEBOOST_cell_73815 ( .a(TIMEBOOST_net_13779), .b(FE_OFN1775_n_13800), .c(FE_OFN1768_n_14054), .o(n_16208) );
na04f04 TIMEBOOST_cell_24664 ( .a(n_9752), .b(g57172_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q), .d(FE_OFN2173_n_8567), .o(n_11584) );
na04f04 TIMEBOOST_cell_24666 ( .a(n_9473), .b(g57487_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q), .d(FE_OFN2178_n_8567), .o(n_11250) );
in01f02 g60658_u0 ( .a(FE_OFN1179_n_3476), .o(g60658_sb) );
in01s02 TIMEBOOST_cell_63536 ( .a(pci_target_unit_fifos_pcir_data_in_185), .o(TIMEBOOST_net_20716) );
in01m01 g60659_u0 ( .a(FE_OFN1181_n_3476), .o(g60659_sb) );
na02s02 TIMEBOOST_cell_48632 ( .a(TIMEBOOST_net_14533), .b(TIMEBOOST_net_12427), .o(TIMEBOOST_net_9470) );
na02s02 TIMEBOOST_cell_39717 ( .a(TIMEBOOST_net_11470), .b(g58412_db), .o(n_9205) );
in01m01 g60660_u0 ( .a(FE_OFN1182_n_3476), .o(g60660_sb) );
na02s02 TIMEBOOST_cell_48582 ( .a(TIMEBOOST_net_14508), .b(FE_OFN1668_n_9477), .o(TIMEBOOST_net_11084) );
na03s01 TIMEBOOST_cell_72726 ( .a(g58194_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q), .c(TIMEBOOST_net_12906), .o(TIMEBOOST_net_14657) );
in01m01 g60661_u0 ( .a(FE_OFN1182_n_3476), .o(g60661_sb) );
na02f02 TIMEBOOST_cell_69675 ( .a(TIMEBOOST_net_22045), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_14797) );
na03f02 TIMEBOOST_cell_34899 ( .a(TIMEBOOST_net_9512), .b(FE_OFN1388_n_8567), .c(g57526_sb), .o(n_11215) );
na02f02 TIMEBOOST_cell_49934 ( .a(TIMEBOOST_net_15184), .b(g62862_sb), .o(n_5242) );
in01m01 g60662_u0 ( .a(FE_OFN1182_n_3476), .o(g60662_sb) );
na03f01 TIMEBOOST_cell_64542 ( .a(n_3741), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q), .c(FE_OFN631_n_4454), .o(TIMEBOOST_net_10390) );
in01m01 g60663_u0 ( .a(FE_OFN1180_n_3476), .o(g60663_sb) );
na02f02 TIMEBOOST_cell_40839 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_12031), .o(n_12761) );
in01f01 g60664_u0 ( .a(FE_OFN1183_n_3476), .o(g60664_sb) );
no02f10 TIMEBOOST_cell_3259 ( .a(TIMEBOOST_net_189), .b(FE_OCPN1841_n_16089), .o(n_3160) );
na02s01 TIMEBOOST_cell_31839 ( .a(wbu_sel_in_312), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__Q), .o(TIMEBOOST_net_10024) );
na02f01 TIMEBOOST_cell_3260 ( .a(n_16151), .b(pci_target_unit_wishbone_master_first_wb_data_access), .o(TIMEBOOST_net_190) );
in01m01 g60665_u0 ( .a(FE_OFN1180_n_3476), .o(g60665_sb) );
na02f02 TIMEBOOST_cell_70979 ( .a(TIMEBOOST_net_22697), .b(g62942_sb), .o(n_5997) );
na02m02 TIMEBOOST_cell_68602 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q), .b(g65024_sb), .o(TIMEBOOST_net_21509) );
na02m02 TIMEBOOST_cell_50306 ( .a(TIMEBOOST_net_15370), .b(g62496_sb), .o(n_6592) );
in01m01 g60666_u0 ( .a(FE_OFN1181_n_3476), .o(g60666_sb) );
in01s01 TIMEBOOST_cell_35526 ( .a(TIMEBOOST_net_10117), .o(TIMEBOOST_net_10092) );
na03f02 TIMEBOOST_cell_73778 ( .a(n_13993), .b(TIMEBOOST_net_13717), .c(FE_OFN1586_n_13736), .o(n_14430) );
in01m01 g60667_u0 ( .a(FE_OFN1180_n_3476), .o(g60667_sb) );
in01s01 TIMEBOOST_cell_35527 ( .a(TIMEBOOST_net_10118), .o(TIMEBOOST_net_10117) );
na02f02 TIMEBOOST_cell_70689 ( .a(TIMEBOOST_net_22552), .b(g62794_sb), .o(n_5399) );
na02s02 TIMEBOOST_cell_50002 ( .a(TIMEBOOST_net_15218), .b(g57972_sb), .o(TIMEBOOST_net_9549) );
in01f02 g60668_u0 ( .a(FE_OFN1180_n_3476), .o(g60668_sb) );
na03m02 TIMEBOOST_cell_65089 ( .a(TIMEBOOST_net_12569), .b(g65417_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q), .o(TIMEBOOST_net_17367) );
na02s01 TIMEBOOST_cell_52647 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_16541) );
in01f02 g60669_u0 ( .a(FE_OFN1179_n_3476), .o(g60669_sb) );
na02m02 TIMEBOOST_cell_68583 ( .a(TIMEBOOST_net_21499), .b(g65889_sb), .o(n_1860) );
in01f01 g60670_u0 ( .a(FE_OFN1183_n_3476), .o(g60670_sb) );
na02f04 TIMEBOOST_cell_3261 ( .a(TIMEBOOST_net_190), .b(n_4874), .o(n_3267) );
na02m02 TIMEBOOST_cell_54653 ( .a(n_7373), .b(n_4907), .o(TIMEBOOST_net_17544) );
na02f01 TIMEBOOST_cell_18041 ( .a(n_2306), .b(n_2755), .o(TIMEBOOST_net_5384) );
in01m01 g60671_u0 ( .a(n_6986), .o(g60671_sb) );
na02m02 TIMEBOOST_cell_50644 ( .a(TIMEBOOST_net_15539), .b(g62997_sb), .o(n_5888) );
na02s01 TIMEBOOST_cell_42785 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q), .o(TIMEBOOST_net_12287) );
in01m01 g60672_u0 ( .a(n_6986), .o(g60672_sb) );
in01s01 TIMEBOOST_cell_73962 ( .a(wbm_dat_i_30_), .o(TIMEBOOST_net_23527) );
na04f04 TIMEBOOST_cell_36848 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q), .b(FE_OFN2168_n_8567), .c(n_9729), .d(g57198_sb), .o(n_11555) );
na02m01 TIMEBOOST_cell_49331 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q), .o(TIMEBOOST_net_14883) );
in01f02 g60673_u0 ( .a(FE_OFN1183_n_3476), .o(g60673_sb) );
in01s01 TIMEBOOST_cell_35528 ( .a(TIMEBOOST_net_10119), .o(TIMEBOOST_net_10094) );
na03m04 TIMEBOOST_cell_72785 ( .a(n_4465), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q), .c(TIMEBOOST_net_12547), .o(TIMEBOOST_net_17082) );
in01f01 g60674_u0 ( .a(n_6986), .o(g60674_sb) );
na03f02 TIMEBOOST_cell_66181 ( .a(TIMEBOOST_net_15234), .b(FE_OFN1179_n_3476), .c(g60609_sb), .o(n_4845) );
na03m10 TIMEBOOST_cell_65334 ( .a(g64131_sb), .b(TIMEBOOST_net_12710), .c(FE_OFN1046_n_16657), .o(n_4031) );
in01m01 g60675_u0 ( .a(FE_OFN923_n_4740), .o(g60675_sb) );
na02m01 TIMEBOOST_cell_53367 ( .a(TIMEBOOST_net_12414), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q), .o(TIMEBOOST_net_16901) );
in01m02 g60676_u0 ( .a(FE_OFN1046_n_16657), .o(g60676_sb) );
no03f04 TIMEBOOST_cell_67021 ( .a(FE_RN_810_0), .b(FE_RN_811_0), .c(FE_RN_812_0), .o(n_14261) );
in01m02 g60677_u0 ( .a(FE_OFN903_n_4736), .o(g60677_sb) );
na02m06 TIMEBOOST_cell_54113 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q), .o(TIMEBOOST_net_17274) );
na03m01 TIMEBOOST_cell_68056 ( .a(TIMEBOOST_net_13985), .b(FE_OFN2114_wishbone_slave_unit_pci_initiator_if_data_source), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q), .o(TIMEBOOST_net_21236) );
in01m02 TIMEBOOST_cell_67746 ( .a(TIMEBOOST_net_21172), .o(TIMEBOOST_net_21173) );
in01f02 g60678_u0 ( .a(FE_OFN1012_n_4734), .o(g60678_sb) );
na04f04 TIMEBOOST_cell_73612 ( .a(n_1855), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q), .c(FE_OFN716_n_8176), .d(g61872_sb), .o(n_8089) );
na03f02 TIMEBOOST_cell_72519 ( .a(TIMEBOOST_net_20177), .b(g65903_sb), .c(FE_OFN959_n_2299), .o(n_2178) );
na03m02 TIMEBOOST_cell_51925 ( .a(n_3761), .b(FE_OFN624_n_4409), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q), .o(TIMEBOOST_net_16180) );
in01m01 g60679_u0 ( .a(FE_OFN1700_n_5751), .o(g60679_sb) );
in01s01 TIMEBOOST_cell_45869 ( .a(pci_target_unit_fifos_pcir_data_in_169), .o(TIMEBOOST_net_13830) );
na02s02 TIMEBOOST_cell_48716 ( .a(TIMEBOOST_net_14575), .b(TIMEBOOST_net_10500), .o(TIMEBOOST_net_9357) );
na02f08 TIMEBOOST_cell_3607 ( .a(TIMEBOOST_net_363), .b(n_3130), .o(n_3141) );
oa12f01 g60680_u0 ( .a(n_7369), .b(n_3316), .c(n_7608), .o(n_7791) );
in01m02 g60681_u0 ( .a(FE_OFN1697_n_5751), .o(g60681_sb) );
in01s01 TIMEBOOST_cell_45870 ( .a(TIMEBOOST_net_13830), .o(TIMEBOOST_net_13831) );
na02f01 g60681_u2 ( .a(n_3331), .b(FE_OFN1697_n_5751), .o(g60681_db) );
na02f20 TIMEBOOST_cell_3449 ( .a(TIMEBOOST_net_284), .b(n_2777), .o(n_3278) );
in01f01 g60682_u0 ( .a(n_6986), .o(g60682_sb) );
na03f02 TIMEBOOST_cell_70584 ( .a(n_3879), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q), .c(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_22500) );
na04f02 TIMEBOOST_cell_36835 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q), .b(FE_OFN1394_n_8567), .c(n_9906), .d(g57181_sb), .o(n_11573) );
na03f02 TIMEBOOST_cell_72944 ( .a(pci_target_unit_del_sync_addr_in_219), .b(g65210_sb), .c(TIMEBOOST_net_7150), .o(n_2679) );
ao12f02 g60684_u0 ( .a(n_4855), .b(FE_OFN1006_n_16288), .c(configuration_pci_err_addr_479), .o(n_7220) );
ao12f02 g60685_u0 ( .a(n_4799), .b(configuration_wb_err_data), .c(FE_OFN1071_n_15729), .o(n_6983) );
in01m01 g60686_u0 ( .a(FE_OFN1036_n_4732), .o(g60686_sb) );
na02m02 TIMEBOOST_cell_69604 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q), .o(TIMEBOOST_net_22010) );
na02m02 TIMEBOOST_cell_68754 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q), .b(FE_OFN661_n_4392), .o(TIMEBOOST_net_21585) );
in01m02 g60687_u0 ( .a(FE_OFN1059_n_4727), .o(g60687_sb) );
na04f04 TIMEBOOST_cell_24668 ( .a(n_9506), .b(g57442_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q), .d(FE_OFN2173_n_8567), .o(n_11293) );
na02s01 TIMEBOOST_cell_63722 ( .a(g61990_sb), .b(g61990_db), .o(TIMEBOOST_net_20847) );
no03f06 TIMEBOOST_cell_67023 ( .a(FE_RN_767_0), .b(FE_RN_768_0), .c(FE_RN_769_0), .o(n_14251) );
in01m02 g60688_u0 ( .a(n_4730), .o(g60688_sb) );
na03f02 TIMEBOOST_cell_73506 ( .a(TIMEBOOST_net_22588), .b(g52452_sb), .c(TIMEBOOST_net_22957), .o(n_14807) );
in01s01 TIMEBOOST_cell_67720 ( .a(TIMEBOOST_net_21146), .o(TIMEBOOST_net_21147) );
in01m10 g60689_u0 ( .a(n_4725), .o(g60689_sb) );
na02f02 TIMEBOOST_cell_70981 ( .a(TIMEBOOST_net_22698), .b(g62641_sb), .o(n_6266) );
na02s01 TIMEBOOST_cell_43831 ( .a(FE_OFN239_n_9832), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q), .o(TIMEBOOST_net_12810) );
na04m02 TIMEBOOST_cell_72549 ( .a(TIMEBOOST_net_21189), .b(g65675_sb), .c(TIMEBOOST_net_12507), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q), .o(TIMEBOOST_net_22314) );
in01m01 g60690_u0 ( .a(n_6986), .o(g60690_sb) );
in01s01 TIMEBOOST_cell_73969 ( .a(TIMEBOOST_net_23533), .o(TIMEBOOST_net_23534) );
in01f01 g60691_u0 ( .a(FE_OFN1699_n_5751), .o(g60691_sb) );
in01s01 TIMEBOOST_cell_45871 ( .a(TIMEBOOST_net_13832), .o(configuration_sync_isr_2_sync_bckp_bit) );
in01m01 g60692_u0 ( .a(n_7608), .o(g60692_sb) );
na02m02 TIMEBOOST_cell_43473 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q), .b(g64276_sb), .o(TIMEBOOST_net_12631) );
na04m01 TIMEBOOST_cell_46765 ( .a(g58139_sb), .b(FE_OFN258_n_9862), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q), .d(g58139_db), .o(TIMEBOOST_net_9363) );
na03f02 TIMEBOOST_cell_73381 ( .a(TIMEBOOST_net_15224), .b(FE_OFN1300_n_5763), .c(g62054_sb), .o(n_7755) );
no02f01 g60693_u0 ( .a(wbu_addr_in_262), .b(n_2970), .o(g60693_p) );
ao12f01 g60693_u1 ( .a(g60693_p), .b(wbu_addr_in_262), .c(n_2970), .o(n_3169) );
no02f01 g60694_u0 ( .a(wbm_adr_o_13_), .b(n_2873), .o(g60694_p) );
ao12f01 g60694_u1 ( .a(g60694_p), .b(wbm_adr_o_13_), .c(n_2873), .o(n_3168) );
no02f08 g60695_u0 ( .a(wbu_addr_in_270), .b(n_2462), .o(g60695_p) );
ao12f04 g60695_u1 ( .a(g60695_p), .b(wbu_addr_in_270), .c(n_2462), .o(n_3167) );
no02m06 g60696_u0 ( .a(n_2460), .b(conf_wb_err_addr_in_954), .o(g60696_p) );
ao12m02 g60696_u1 ( .a(g60696_p), .b(conf_wb_err_addr_in_954), .c(n_2460), .o(n_3345) );
na03f02 TIMEBOOST_cell_66046 ( .a(TIMEBOOST_net_17346), .b(n_7618), .c(g59805_sb), .o(n_7619) );
na03m02 TIMEBOOST_cell_72867 ( .a(TIMEBOOST_net_21727), .b(g65322_sb), .c(TIMEBOOST_net_21957), .o(TIMEBOOST_net_20523) );
na03f02 TIMEBOOST_cell_65940 ( .a(TIMEBOOST_net_20440), .b(FE_OFN1166_n_5615), .c(g62117_sb), .o(n_5579) );
na02f01 TIMEBOOST_cell_18203 ( .a(n_2418), .b(n_7078), .o(TIMEBOOST_net_5465) );
no02f02 g61546_u0 ( .a(n_4167), .b(n_3227), .o(n_4691) );
in01s01 TIMEBOOST_cell_64265 ( .a(TIMEBOOST_net_21120), .o(TIMEBOOST_net_21121) );
na04f04 TIMEBOOST_cell_24847 ( .a(wbs_dat_o_26_), .b(g52521_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_125), .d(FE_OFN2242_g52675_p), .o(n_13698) );
na04f04 TIMEBOOST_cell_24846 ( .a(wbs_dat_o_27_), .b(g52522_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_126), .d(FE_OFN2243_g52675_p), .o(n_13735) );
oa12f02 g61555_u0 ( .a(n_14909), .b(n_8450), .c(n_8511), .o(n_8451) );
oa12f02 g61556_u0 ( .a(n_14908), .b(FE_OFN2086_n_8448), .c(n_8511), .o(n_8449) );
oa12f01 g61557_u0 ( .a(configuration_pci_err_cs_bit0), .b(n_8446), .c(n_3030), .o(n_8447) );
oa12f04 g61558_u0 ( .a(wbu_bar1_in), .b(n_8468), .c(n_8511), .o(n_7790) );
no02f06 g61559_u0 ( .a(n_2750), .b(n_2735), .o(n_2751) );
oa12f04 g61560_u0 ( .a(wbu_am1_in), .b(n_8514), .c(n_8511), .o(n_8515) );
oa12f02 g61561_u0 ( .a(wbu_map_in_131), .b(n_8468), .c(n_3030), .o(n_7789) );
oa12f02 g61562_u0 ( .a(wbu_map_in_132), .b(n_8465), .c(n_3030), .o(n_7788) );
oa12f02 g61563_u0 ( .a(wbu_bar2_in), .b(n_8465), .c(n_8511), .o(n_7787) );
na04f04 TIMEBOOST_cell_24648 ( .a(n_9220), .b(g57235_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q), .d(FE_OFN2174_n_8567), .o(n_10832) );
oa12f04 g61565_u0 ( .a(wbu_am2_in), .b(n_8512), .c(n_8511), .o(n_8513) );
oa12s02 g61566_u0 ( .a(configuration_sync_command_bit8), .b(n_7785), .c(n_2651), .o(n_7786) );
oa12f02 g61567_u0 ( .a(configuration_wb_err_cs_bit0), .b(n_8444), .c(n_3030), .o(n_8445) );
na02f08 g61569_u0 ( .a(n_2967), .b(n_2970), .o(g61569_p) );
in01f06 g61569_u1 ( .a(g61569_p), .o(n_2968) );
na02f02 g61570_u0 ( .a(n_1971), .b(n_2970), .o(g61570_p) );
in01f02 g61570_u1 ( .a(g61570_p), .o(n_2971) );
na02f01 g61571_u0 ( .a(n_4666), .b(n_7608), .o(n_7369) );
no02m02 g61572_u0 ( .a(n_7818), .b(n_3030), .o(g61572_p) );
in01m02 g61572_u1 ( .a(g61572_p), .o(n_7473) );
no02f02 g61573_u0 ( .a(n_4172), .b(n_7031), .o(n_4819) );
no02f02 g61574_u0 ( .a(n_4171), .b(n_7031), .o(n_4820) );
no02f10 g61575_u0 ( .a(n_7498), .b(n_8511), .o(g61575_p) );
in01f08 g61575_u1 ( .a(g61575_p), .o(n_7065) );
no02f02 g61576_u0 ( .a(n_5549), .b(n_4146), .o(n_7213) );
no02f04 g61577_u0 ( .a(n_4170), .b(n_7031), .o(n_4823) );
no02f02 g61578_u0 ( .a(n_7031), .b(n_4169), .o(n_4824) );
no02f02 g61579_u0 ( .a(FE_OFN1180_n_3476), .b(n_200), .o(n_4694) );
no02f02 g61580_u0 ( .a(n_4168), .b(n_7031), .o(n_4825) );
no02f06 g61581_u0 ( .a(n_8476), .b(n_3030), .o(g61581_p) );
in01f04 g61581_u1 ( .a(g61581_p), .o(n_7611) );
na02f02 g61582_u0 ( .a(n_4155), .b(n_2768), .o(g61582_p) );
in01f02 g61582_u1 ( .a(g61582_p), .o(n_4826) );
in01f04 g61583_u0 ( .a(n_15377), .o(n_7567) );
in01f03 g61586_u0 ( .a(n_7216), .o(n_13814) );
in01f08 g61587_u0 ( .a(n_6989), .o(n_7216) );
in01f08 g61589_u0 ( .a(n_15467), .o(n_6989) );
no02f02 g61593_u0 ( .a(n_4786), .b(n_4812), .o(n_5717) );
na02f02 g61594_u0 ( .a(n_7738), .b(n_1759), .o(n_8472) );
ao12f02 g61595_u0 ( .a(n_7552), .b(n_4780), .c(n_3393), .o(n_7075) );
na02s01 TIMEBOOST_cell_48435 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_14435) );
no02f02 g61597_u0 ( .a(FE_OFN1183_n_3476), .b(n_3342), .o(g61597_p) );
in01f02 g61597_u1 ( .a(g61597_p), .o(n_4871) );
in01s01 TIMEBOOST_cell_35529 ( .a(TIMEBOOST_net_10120), .o(TIMEBOOST_net_10119) );
na02f03 g61599_u0 ( .a(FE_OFN1183_n_3476), .b(configuration_pci_err_cs_bit_467), .o(n_4211) );
na02f02 g61600_u0 ( .a(FE_OFN1183_n_3476), .b(configuration_pci_err_cs_bit_468), .o(n_4212) );
na02f02 g61601_u0 ( .a(FE_OFN1181_n_3476), .b(configuration_pci_err_cs_bit_469), .o(n_4213) );
na02f03 g61602_u0 ( .a(FE_OFN1181_n_3476), .b(configuration_pci_err_cs_bit_470), .o(n_4216) );
na02f01 TIMEBOOST_cell_71048 ( .a(TIMEBOOST_net_17361), .b(FE_OFN1273_n_4096), .o(TIMEBOOST_net_22732) );
na02m04 TIMEBOOST_cell_51647 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q), .o(TIMEBOOST_net_16041) );
no02f04 g61606_u0 ( .a(n_8521), .b(n_3030), .o(g61606_p) );
in01f02 g61606_u1 ( .a(g61606_p), .o(n_7813) );
no02f02 g61608_u0 ( .a(n_3153), .b(FE_OFN1144_n_15261), .o(n_3375) );
no02f02 g61609_u0 ( .a(n_3154), .b(FE_OFN1143_n_15261), .o(n_3376) );
no02f02 g61610_u0 ( .a(n_3467), .b(FE_OFN1145_n_15261), .o(n_4504) );
na02f10 g61611_u0 ( .a(n_2460), .b(n_2475), .o(n_2476) );
in01s01 TIMEBOOST_cell_45872 ( .a(TIMEBOOST_net_13833), .o(TIMEBOOST_net_13832) );
ao12f02 g61614_u0 ( .a(n_7608), .b(n_2807), .c(n_3166), .o(n_7401) );
in01f02 g61616_u0 ( .a(n_5228), .o(n_5229) );
na02f02 g61617_u0 ( .a(n_7078), .b(n_692), .o(g61617_p) );
in01f02 g61617_u1 ( .a(g61617_p), .o(n_5228) );
in01s01 TIMEBOOST_cell_45873 ( .a(TIMEBOOST_net_13834), .o(configuration_sync_pci_err_cs_8_sync_bckp_bit) );
in01f02 g61618_u3 ( .a(g61618_p), .o(n_7115) );
in01s01 TIMEBOOST_cell_63569 ( .a(TIMEBOOST_net_20749), .o(TIMEBOOST_net_20748) );
na02f01 g61620_u0 ( .a(n_7608), .b(n_16512), .o(n_7339) );
no02f04 g61621_u0 ( .a(n_4197), .b(n_1258), .o(n_4198) );
na02f02 g61622_u0 ( .a(n_15689), .b(n_7622), .o(g61622_p) );
in01f02 g61622_u1 ( .a(g61622_p), .o(n_4822) );
no02f10 g61636_u0 ( .a(n_7498), .b(n_2651), .o(g61636_p) );
in01f08 g61636_u1 ( .a(g61636_p), .o(n_7056) );
no02f10 g61637_u0 ( .a(n_7498), .b(n_2648), .o(g61637_p) );
in01f08 g61637_u1 ( .a(g61637_p), .o(n_7072) );
in01f02 g61641_u0 ( .a(n_16452), .o(n_7096) );
na03m02 TIMEBOOST_cell_73018 ( .a(TIMEBOOST_net_17255), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .c(g52636_sb), .o(n_14755) );
na02f01 TIMEBOOST_cell_26274 ( .a(TIMEBOOST_net_7241), .b(TIMEBOOST_net_557), .o(n_4105) );
no02s01 g61647_u0 ( .a(n_2284), .b(n_1551), .o(n_2285) );
oa12f02 g61649_u0 ( .a(n_7743), .b(FE_OFN1169_n_5592), .c(n_24), .o(n_8510) );
in01s01 TIMEBOOST_cell_45874 ( .a(TIMEBOOST_net_13835), .o(TIMEBOOST_net_13834) );
na02f02 g61651_u0 ( .a(n_7734), .b(conf_target_abort_recv_in), .o(n_8509) );
ao12f02 g61652_u0 ( .a(n_4808), .b(n_14928), .c(FE_OCPN1900_n_16810), .o(n_6978) );
na02m02 TIMEBOOST_cell_44702 ( .a(TIMEBOOST_net_13245), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_11630) );
no02f02 g61654_u0 ( .a(n_6944), .b(n_7398), .o(g61654_p) );
in01f02 g61654_u1 ( .a(g61654_p), .o(n_7399) );
na02m20 TIMEBOOST_cell_52691 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q), .o(TIMEBOOST_net_16563) );
oa12s02 g61656_u0 ( .a(n_7742), .b(n_369), .c(FE_OFN1169_n_5592), .o(n_8508) );
na02f02 g61657_u0 ( .a(n_2352), .b(n_3498), .o(n_3499) );
na03s01 TIMEBOOST_cell_48817 ( .a(g58051_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q), .c(g58064_db), .o(TIMEBOOST_net_14626) );
in01m04 g61660_u0 ( .a(n_2420), .o(n_2421) );
no02f04 g61661_u0 ( .a(n_1389), .b(n_2295), .o(n_2420) );
na02f02 g61662_u0 ( .a(n_2369), .b(n_3363), .o(n_3364) );
na02f02 g61663_u0 ( .a(n_2359), .b(n_4894), .o(n_4895) );
na02f01 g61664_u0 ( .a(n_7737), .b(n_2494), .o(n_8506) );
in01s01 TIMEBOOST_cell_45945 ( .a(TIMEBOOST_net_13937), .o(TIMEBOOST_net_13906) );
in01f02 g61666_u0 ( .a(n_3392), .o(n_3832) );
ao12f04 g61667_u0 ( .a(n_3391), .b(n_3160), .c(n_4078), .o(n_3392) );
na02m10 TIMEBOOST_cell_45823 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q), .o(TIMEBOOST_net_13806) );
ao12f02 g61670_u0 ( .a(n_3157), .b(n_1662), .c(wbm_rty_i), .o(n_3076) );
ao12f02 g61671_u0 ( .a(n_4896), .b(n_1200), .c(pci_target_unit_wishbone_master_c_state_2_), .o(n_4897) );
ao12f02 g61672_u0 ( .a(n_4683), .b(FE_OFN1006_n_16288), .c(configuration_pci_err_addr_480), .o(n_4899) );
in01m02 g61673_u0 ( .a(n_2424), .o(n_2425) );
no02f08 g61674_u0 ( .a(n_1392), .b(n_2275), .o(n_2424) );
na02f01 g61675_u0 ( .a(n_2371), .b(n_4894), .o(n_5640) );
in01f01 g61676_u0 ( .a(FE_OFN1166_n_5615), .o(g61676_sb) );
na03m02 TIMEBOOST_cell_68582 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(FE_OFN634_n_4454), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q), .o(TIMEBOOST_net_21499) );
na03f02 TIMEBOOST_cell_66306 ( .a(TIMEBOOST_net_20572), .b(n_6431), .c(g62396_sb), .o(n_7388) );
na02s02 TIMEBOOST_cell_48868 ( .a(TIMEBOOST_net_14651), .b(FE_OFN247_n_9112), .o(n_9071) );
oa12f02 g61677_u0 ( .a(n_4718), .b(n_4680), .c(n_3480), .o(n_4717) );
oa12f02 g61678_u0 ( .a(n_7565), .b(n_8440), .c(n_4784), .o(n_8442) );
oa12m02 g61679_u0 ( .a(n_7564), .b(n_8440), .c(n_4785), .o(n_8441) );
oa12m02 g61680_u0 ( .a(n_7562), .b(n_8440), .c(n_4782), .o(n_8439) );
oa12m02 g61681_u0 ( .a(n_7561), .b(n_8440), .c(n_4781), .o(n_8438) );
oa12f02 g61684_u0 ( .a(n_7559), .b(n_8440), .c(n_4629), .o(n_8437) );
oa12f01 g61685_u0 ( .a(n_7560), .b(n_8440), .c(n_4631), .o(n_8436) );
oa12f02 g61686_u0 ( .a(n_7558), .b(n_8440), .c(n_4633), .o(n_8434) );
ao12f02 g61687_u0 ( .a(n_3339), .b(conf_wb_err_addr_in_960), .c(FE_OFN1142_n_15261), .o(n_4161) );
ao12f02 g61688_u0 ( .a(n_3468), .b(conf_wb_err_addr_in_964), .c(FE_OFN1145_n_15261), .o(n_4668) );
no02f04 g61689_u0 ( .a(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .b(n_3141), .o(g61689_p) );
ao12f02 g61689_u1 ( .a(g61689_p), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .c(n_3141), .o(n_4162) );
oa12f02 g61690_u0 ( .a(n_7731), .b(n_1755), .c(FE_OFN2079_n_8069), .o(n_8502) );
ao12f02 g61691_u0 ( .a(n_3338), .b(conf_wb_err_addr_in_961), .c(FE_OFN1144_n_15261), .o(n_3474) );
oa12f01 g61692_u0 ( .a(n_7557), .b(n_8440), .c(n_4628), .o(n_8433) );
no02f06 g61693_u0 ( .a(n_2939), .b(n_1461), .o(g61693_p) );
ao12f06 g61693_u1 ( .a(g61693_p), .b(n_1461), .c(n_2939), .o(n_3466) );
oa12s02 g61694_u0 ( .a(n_4813), .b(FE_OFN1169_n_5592), .c(n_2494), .o(n_6218) );
ao12s01 g61695_u0 ( .a(n_7571), .b(configuration_sync_isr_2_delayed_bckp_bit), .c(configuration_sync_isr_2_sync_bckp_bit), .o(n_8432) );
ao12s01 g61696_u0 ( .a(n_7574), .b(configuration_sync_pci_err_cs_8_delayed_bckp_bit), .c(configuration_sync_pci_err_cs_8_sync_bckp_bit), .o(n_8431) );
in01f01 g61697_u0 ( .a(FE_OFN1095_g64577_p), .o(g61697_sb) );
na02s02 TIMEBOOST_cell_28193 ( .a(g65780_sb), .b(TIMEBOOST_net_21181), .o(TIMEBOOST_net_8201) );
na04m02 TIMEBOOST_cell_65130 ( .a(g65092_sb), .b(FE_OFN618_n_4490), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q), .d(n_4482), .o(TIMEBOOST_net_7595) );
in01s01 g61698_u0 ( .a(FE_OFN1097_g64577_p), .o(g61698_sb) );
na03f02 TIMEBOOST_cell_73310 ( .a(TIMEBOOST_net_8797), .b(FE_OFN2105_g64577_p), .c(g62809_sb), .o(n_5361) );
na02m01 g61698_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q), .b(FE_OFN1097_g64577_p), .o(g61698_db) );
na02f02 TIMEBOOST_cell_50314 ( .a(TIMEBOOST_net_15374), .b(g62405_sb), .o(n_6789) );
in01m02 g61699_u0 ( .a(FE_OFN720_n_8060), .o(g61699_sb) );
na02s02 TIMEBOOST_cell_38272 ( .a(g58062_sb), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_10748) );
na03m02 TIMEBOOST_cell_73104 ( .a(TIMEBOOST_net_11076), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q), .c(TIMEBOOST_net_7259), .o(TIMEBOOST_net_17394) );
in01f02 g61700_u0 ( .a(FE_OFN2081_n_8176), .o(g61700_sb) );
na02f40 TIMEBOOST_cell_29059 ( .a(pciu_pciif_idsel_reg_in), .b(n_343), .o(TIMEBOOST_net_8634) );
na02m01 TIMEBOOST_cell_53369 ( .a(FE_OFN625_n_4409), .b(n_0), .o(TIMEBOOST_net_16902) );
na02f02 TIMEBOOST_cell_53297 ( .a(wbu_addr_in_272), .b(n_3138), .o(TIMEBOOST_net_16866) );
in01m02 g61701_u0 ( .a(FE_OFN720_n_8060), .o(g61701_sb) );
na02m10 TIMEBOOST_cell_28991 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q), .o(TIMEBOOST_net_8600) );
in01s01 g61702_u0 ( .a(n_8176), .o(g61702_sb) );
in01s01 TIMEBOOST_cell_73841 ( .a(TIMEBOOST_net_23405), .o(TIMEBOOST_net_23406) );
na02s01 g61702_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q), .b(n_8176), .o(g61702_db) );
na03m02 TIMEBOOST_cell_72703 ( .a(g64887_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q), .c(TIMEBOOST_net_16597), .o(TIMEBOOST_net_13244) );
in01s01 g61703_u0 ( .a(n_8407), .o(g61703_sb) );
na03f02 TIMEBOOST_cell_73613 ( .a(TIMEBOOST_net_17561), .b(FE_OFN1253_n_4143), .c(g62417_sb), .o(n_6763) );
na02s01 g61703_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q), .b(n_8407), .o(g61703_db) );
na03f02 TIMEBOOST_cell_66280 ( .a(wbm_dat_o_3_), .b(g60664_sb), .c(g60664_db), .o(n_5655) );
in01m01 g61704_u0 ( .a(FE_OFN716_n_8176), .o(g61704_sb) );
na03f02 TIMEBOOST_cell_67025 ( .a(FE_OFN1602_n_13995), .b(TIMEBOOST_net_13747), .c(FE_OCPN2219_n_13997), .o(n_14443) );
na02m10 TIMEBOOST_cell_45765 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q), .o(TIMEBOOST_net_13777) );
in01s01 g61705_u0 ( .a(n_7102), .o(g61705_sb) );
na03f02 TIMEBOOST_cell_66598 ( .a(TIMEBOOST_net_17549), .b(FE_OFN1193_n_6935), .c(g62916_sb), .o(n_6047) );
na02s01 g61705_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q), .b(n_7102), .o(g61705_db) );
no02f04 TIMEBOOST_cell_68064 ( .a(FE_OCPN1849_n_15998), .b(FE_OCPN1868_n_16289), .o(TIMEBOOST_net_21240) );
in01f02 g61706_u0 ( .a(FE_OFN714_n_8140), .o(g61706_sb) );
na04m04 TIMEBOOST_cell_72885 ( .a(TIMEBOOST_net_10319), .b(g65935_sb), .c(g62012_db), .d(g62012_sb), .o(n_7871) );
na02f02 TIMEBOOST_cell_70201 ( .a(TIMEBOOST_net_22308), .b(g54235_sb), .o(n_13653) );
na02f02 TIMEBOOST_cell_37301 ( .a(TIMEBOOST_net_10262), .b(n_14070), .o(TIMEBOOST_net_501) );
in01s01 g61707_u0 ( .a(n_8272), .o(g61707_sb) );
na03f02 TIMEBOOST_cell_67028 ( .a(FE_OFN1606_n_13997), .b(TIMEBOOST_net_13745), .c(FE_OFN1599_n_13995), .o(n_14461) );
na02f04 TIMEBOOST_cell_52468 ( .a(TIMEBOOST_net_16451), .b(g58375_db), .o(n_9454) );
na03m02 TIMEBOOST_cell_536 ( .a(n_1904), .b(g61858_sb), .c(g61858_db), .o(n_8123) );
in01s01 g61708_u0 ( .a(n_8069), .o(g61708_sb) );
na02s01 g61708_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q), .b(n_8069), .o(g61708_db) );
in01s01 g61709_u0 ( .a(n_8407), .o(g61709_sb) );
na02s01 g61709_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q), .b(n_8407), .o(g61709_db) );
in01s01 g61710_u0 ( .a(n_8140), .o(g61710_sb) );
na02s01 g61710_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q), .b(n_8140), .o(g61710_db) );
na02s02 TIMEBOOST_cell_54256 ( .a(TIMEBOOST_net_17345), .b(g58201_db), .o(TIMEBOOST_net_9450) );
in01m01 g61711_u0 ( .a(FE_OFN702_n_7845), .o(g61711_sb) );
na03s02 TIMEBOOST_cell_21311 ( .a(FE_OFN227_n_9841), .b(g58108_sb), .c(g58122_db), .o(n_9670) );
na02f01 TIMEBOOST_cell_68159 ( .a(TIMEBOOST_net_21287), .b(wbu_addr_in_257), .o(TIMEBOOST_net_12306) );
na03s01 TIMEBOOST_cell_41937 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q), .b(g58370_sb), .c(g58370_db), .o(n_9011) );
in01f01 g61712_u0 ( .a(FE_OFN707_n_8119), .o(g61712_sb) );
na02m10 TIMEBOOST_cell_43649 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_12719) );
na02f01 TIMEBOOST_cell_68327 ( .a(TIMEBOOST_net_21371), .b(FE_OFN611_n_4501), .o(TIMEBOOST_net_237) );
na02m04 TIMEBOOST_cell_69677 ( .a(TIMEBOOST_net_22046), .b(FE_OFN1806_n_4501), .o(TIMEBOOST_net_16378) );
na02s02 TIMEBOOST_cell_48788 ( .a(TIMEBOOST_net_14611), .b(TIMEBOOST_net_11080), .o(TIMEBOOST_net_9442) );
na02s01 g61713_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q), .b(n_7102), .o(g61713_db) );
na02s01 TIMEBOOST_cell_48535 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q), .b(g65814_sb), .o(TIMEBOOST_net_14485) );
in01m01 g61714_u0 ( .a(FE_OFN1812_n_7845), .o(g61714_sb) );
in01m03 TIMEBOOST_cell_31888 ( .a(TIMEBOOST_net_10051), .o(TIMEBOOST_net_10052) );
in01s01 TIMEBOOST_cell_67724 ( .a(TIMEBOOST_net_21150), .o(TIMEBOOST_net_21151) );
na03f02 TIMEBOOST_cell_66120 ( .a(TIMEBOOST_net_16707), .b(FE_OFN1300_n_5763), .c(g62057_sb), .o(n_7752) );
in01s01 g61715_u0 ( .a(n_8232), .o(g61715_sb) );
na02m01 TIMEBOOST_cell_54257 ( .a(n_16860), .b(n_4086), .o(TIMEBOOST_net_17346) );
na02m01 g61715_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q), .b(n_8232), .o(g61715_db) );
na02f02 TIMEBOOST_cell_38979 ( .a(TIMEBOOST_net_11101), .b(FE_OFN1149_n_13249), .o(TIMEBOOST_net_350) );
in01m01 g61716_u0 ( .a(FE_OFN720_n_8060), .o(g61716_sb) );
na02m01 TIMEBOOST_cell_42806 ( .a(TIMEBOOST_net_12297), .b(FE_OFN935_n_2292), .o(TIMEBOOST_net_10236) );
na03m02 TIMEBOOST_cell_72923 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q), .b(g65410_sb), .c(TIMEBOOST_net_22107), .o(TIMEBOOST_net_20953) );
na03f04 TIMEBOOST_cell_65951 ( .a(TIMEBOOST_net_20438), .b(FE_OFN1174_n_5592), .c(g62073_sb), .o(n_5638) );
in01s01 g61717_u0 ( .a(n_8232), .o(g61717_sb) );
na02s01 g61717_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q), .b(n_8232), .o(g61717_db) );
in01f01 g61718_u0 ( .a(FE_OFN2081_n_8176), .o(g61718_sb) );
na02f01 TIMEBOOST_cell_50713 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_386), .b(FE_OFN1001_n_15978), .o(TIMEBOOST_net_15574) );
in01s01 g61719_u0 ( .a(FE_OFN704_n_8069), .o(g61719_sb) );
na03f02 TIMEBOOST_cell_73507 ( .a(TIMEBOOST_net_22638), .b(g62068_db), .c(TIMEBOOST_net_9122), .o(n_14811) );
na03f01 TIMEBOOST_cell_64539 ( .a(FE_OFN679_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q), .c(n_3783), .o(TIMEBOOST_net_14319) );
na03m02 TIMEBOOST_cell_64911 ( .a(TIMEBOOST_net_20269), .b(g64966_sb), .c(g64966_db), .o(TIMEBOOST_net_13231) );
in01f01 g61720_u0 ( .a(FE_OFN2084_n_8407), .o(g61720_sb) );
na02f01 TIMEBOOST_cell_53333 ( .a(n_2675), .b(FE_OFN783_n_2678), .o(TIMEBOOST_net_16884) );
na02m01 TIMEBOOST_cell_53999 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_127), .o(TIMEBOOST_net_17217) );
in01f02 g61721_u0 ( .a(FE_OFN717_n_8176), .o(g61721_sb) );
na02f02 TIMEBOOST_cell_53299 ( .a(wbu_addr_in_268), .b(n_3140), .o(TIMEBOOST_net_16867) );
na03f02 TIMEBOOST_cell_66672 ( .a(TIMEBOOST_net_17537), .b(FE_OFN1212_n_4151), .c(g62458_sb), .o(n_6680) );
in01f02 g61722_u0 ( .a(FE_OFN2081_n_8176), .o(g61722_sb) );
na03f02 TIMEBOOST_cell_66278 ( .a(wbm_adr_o_11_), .b(g60606_sb), .c(TIMEBOOST_net_5516), .o(n_4848) );
na02m02 TIMEBOOST_cell_69904 ( .a(g64255_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q), .o(TIMEBOOST_net_22160) );
in01f02 g61723_u0 ( .a(FE_OFN713_n_8140), .o(g61723_sb) );
na02m20 TIMEBOOST_cell_53463 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_777), .o(TIMEBOOST_net_16949) );
na03f02 TIMEBOOST_cell_66811 ( .a(TIMEBOOST_net_17172), .b(FE_OFN1345_n_8567), .c(g57078_sb), .o(n_11665) );
in01m02 g61724_u0 ( .a(FE_OFN717_n_8176), .o(g61724_sb) );
na03m02 TIMEBOOST_cell_65521 ( .a(g58273_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q), .c(TIMEBOOST_net_12976), .o(TIMEBOOST_net_9503) );
na03m02 TIMEBOOST_cell_72788 ( .a(TIMEBOOST_net_21570), .b(g64892_sb), .c(TIMEBOOST_net_21840), .o(TIMEBOOST_net_17386) );
na02s01 TIMEBOOST_cell_63720 ( .a(g61726_sb), .b(g61726_db), .o(TIMEBOOST_net_20846) );
in01m01 g61725_u0 ( .a(FE_OFN1812_n_7845), .o(g61725_sb) );
na03f02 TIMEBOOST_cell_73072 ( .a(TIMEBOOST_net_8733), .b(FE_OFN2079_n_8069), .c(g62058_sb), .o(n_7836) );
in01s01 g61726_u0 ( .a(n_8069), .o(g61726_sb) );
na02m02 TIMEBOOST_cell_68269 ( .a(TIMEBOOST_net_21342), .b(g65701_db), .o(n_2201) );
na02s01 g61726_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q), .b(n_8069), .o(g61726_db) );
na02s02 TIMEBOOST_cell_49456 ( .a(TIMEBOOST_net_14945), .b(g58239_sb), .o(TIMEBOOST_net_11217) );
in01s01 g61727_u0 ( .a(FE_OFN2257_n_8060), .o(g61727_sb) );
na03f02 TIMEBOOST_cell_73200 ( .a(TIMEBOOST_net_20876), .b(FE_OFN1092_g64577_p), .c(g63561_sb), .o(n_4113) );
na02f02 TIMEBOOST_cell_69775 ( .a(TIMEBOOST_net_22095), .b(g65946_db), .o(n_2575) );
in01f02 g61728_u0 ( .a(FE_OFN713_n_8140), .o(g61728_sb) );
in01f02 g61729_u0 ( .a(FE_OFN713_n_8140), .o(g61729_sb) );
no03f04 TIMEBOOST_cell_73696 ( .a(n_4644), .b(n_7552), .c(n_4878), .o(g59346_p) );
na02f02 TIMEBOOST_cell_70649 ( .a(TIMEBOOST_net_22532), .b(g62740_sb), .o(n_5499) );
in01m01 g61730_u0 ( .a(FE_OFN2256_n_8060), .o(g61730_sb) );
in01s01 TIMEBOOST_cell_67769 ( .a(pci_target_unit_fifos_pcir_data_in_182), .o(TIMEBOOST_net_21196) );
na02m02 TIMEBOOST_cell_52697 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q), .b(TIMEBOOST_net_12329), .o(TIMEBOOST_net_16566) );
in01s02 g61731_u0 ( .a(FE_OFN701_n_7845), .o(g61731_sb) );
in01m01 g61732_u0 ( .a(n_8119), .o(g61732_sb) );
na02s01 TIMEBOOST_cell_25617 ( .a(g61705_sb), .b(g61705_db), .o(TIMEBOOST_net_6913) );
na02m01 g61732_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q), .b(n_8119), .o(g61732_db) );
na02m02 TIMEBOOST_cell_69924 ( .a(n_4498), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_22170) );
in01f02 g61733_u0 ( .a(FE_OFN2212_n_8407), .o(g61733_sb) );
na04m02 TIMEBOOST_cell_67895 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q), .b(n_8272), .c(g61939_sb), .d(n_1567), .o(n_7945) );
in01s01 g61734_u0 ( .a(n_8069), .o(g61734_sb) );
na02s01 g61734_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q), .b(n_8069), .o(g61734_db) );
in01s01 g61735_u0 ( .a(n_8232), .o(g61735_sb) );
na02s01 g61735_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q), .b(n_8232), .o(g61735_db) );
na02m01 TIMEBOOST_cell_69042 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q), .b(FE_OFN653_n_4508), .o(TIMEBOOST_net_21729) );
in01s01 g61736_u0 ( .a(n_8069), .o(g61736_sb) );
na02m02 TIMEBOOST_cell_52411 ( .a(TIMEBOOST_net_13053), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_16423) );
na02s01 g61736_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q), .b(n_8069), .o(g61736_db) );
in01s01 TIMEBOOST_cell_45924 ( .a(TIMEBOOST_net_13884), .o(TIMEBOOST_net_13885) );
in01m01 g61737_u0 ( .a(FE_OFN719_n_8060), .o(g61737_sb) );
in01s01 g61738_u0 ( .a(n_8272), .o(g61738_sb) );
in01s01 TIMEBOOST_cell_45925 ( .a(pci_target_unit_fifos_pcir_data_in_175), .o(TIMEBOOST_net_13886) );
na03f02 TIMEBOOST_cell_73508 ( .a(TIMEBOOST_net_13365), .b(n_6232), .c(g62921_sb), .o(n_6039) );
in01f01 g61739_u0 ( .a(FE_OFN714_n_8140), .o(g61739_sb) );
in01s01 TIMEBOOST_cell_63555 ( .a(TIMEBOOST_net_20735), .o(TIMEBOOST_net_20734) );
in01s01 g61740_u0 ( .a(n_8069), .o(g61740_sb) );
na02s01 TIMEBOOST_cell_31007 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_30__Q), .b(FE_OFN239_n_9832), .o(TIMEBOOST_net_9608) );
na02s01 g61740_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q), .b(n_8069), .o(g61740_db) );
na04f04 TIMEBOOST_cell_24153 ( .a(n_9478), .b(g57481_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q), .d(FE_OFN1419_n_8567), .o(n_11255) );
in01s01 g61741_u0 ( .a(n_8232), .o(g61741_sb) );
na04f04 TIMEBOOST_cell_24154 ( .a(n_9115), .b(g57098_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q), .d(FE_OFN1405_n_8567), .o(n_10483) );
na02s01 g61741_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q), .b(n_8232), .o(g61741_db) );
na02m02 TIMEBOOST_cell_69903 ( .a(TIMEBOOST_net_22159), .b(g64173_sb), .o(TIMEBOOST_net_17328) );
in01s01 g61742_u0 ( .a(n_8119), .o(g61742_sb) );
na03f02 TIMEBOOST_cell_73614 ( .a(TIMEBOOST_net_17093), .b(FE_OFN1284_n_4097), .c(g62567_sb), .o(n_6423) );
na02s01 g61742_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q), .b(n_8119), .o(g61742_db) );
in01m01 g61743_u0 ( .a(n_8407), .o(g61743_sb) );
na03f02 TIMEBOOST_cell_66458 ( .a(TIMEBOOST_net_17137), .b(FE_OFN1317_n_6624), .c(g62486_sb), .o(n_6615) );
na02m01 g61743_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q), .b(n_8407), .o(g61743_db) );
na03f02 TIMEBOOST_cell_72961 ( .a(TIMEBOOST_net_21821), .b(g65275_sb), .c(TIMEBOOST_net_22109), .o(TIMEBOOST_net_20528) );
in01m01 g61744_u0 ( .a(FE_OFN720_n_8060), .o(g61744_sb) );
na04s02 TIMEBOOST_cell_72911 ( .a(TIMEBOOST_net_10531), .b(g65762_sb), .c(g61779_sb), .d(g61779_db), .o(n_8248) );
na02m01 TIMEBOOST_cell_52507 ( .a(FE_OFN576_n_9902), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q), .o(TIMEBOOST_net_16471) );
in01f02 g61745_u0 ( .a(FE_OFN716_n_8176), .o(g61745_sb) );
na02m02 TIMEBOOST_cell_48670 ( .a(TIMEBOOST_net_14552), .b(FE_OFN1057_n_4727), .o(TIMEBOOST_net_12840) );
na04m08 TIMEBOOST_cell_67838 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q), .b(FE_OFN1624_n_4438), .c(g64993_sb), .d(n_4442), .o(n_4357) );
na03f06 TIMEBOOST_cell_73311 ( .a(TIMEBOOST_net_9916), .b(FE_OFN1133_g64577_p), .c(g62750_sb), .o(n_5481) );
in01m01 g61746_u0 ( .a(n_8232), .o(g61746_sb) );
na02m02 TIMEBOOST_cell_52412 ( .a(TIMEBOOST_net_16423), .b(g63125_sb), .o(n_5003) );
na02m01 g61746_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q), .b(n_8232), .o(g61746_db) );
no03f04 TIMEBOOST_cell_47136 ( .a(FE_RN_48_0), .b(FE_OFN1709_n_4868), .c(FE_RN_49_0), .o(TIMEBOOST_net_477) );
in01f01 g61747_u0 ( .a(FE_OFN712_n_8140), .o(g61747_sb) );
na02s02 TIMEBOOST_cell_38562 ( .a(g58191_sb), .b(FE_OFN241_n_9830), .o(TIMEBOOST_net_10893) );
na02m02 TIMEBOOST_cell_47999 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q), .o(TIMEBOOST_net_14217) );
in01s01 g61748_u0 ( .a(n_8232), .o(g61748_sb) );
no02f02 TIMEBOOST_cell_51520 ( .a(TIMEBOOST_net_15977), .b(n_7708), .o(n_13565) );
na02m01 g61748_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q), .b(n_8232), .o(g61748_db) );
na02s01 TIMEBOOST_cell_52649 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q), .o(TIMEBOOST_net_16542) );
in01s01 g61749_u0 ( .a(n_8069), .o(g61749_sb) );
na02s01 g61749_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q), .b(n_8069), .o(g61749_db) );
na02f02 TIMEBOOST_cell_52413 ( .a(TIMEBOOST_net_13081), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_16424) );
in01f02 g61750_u0 ( .a(FE_OFN717_n_8176), .o(g61750_sb) );
na03f02 TIMEBOOST_cell_66454 ( .a(TIMEBOOST_net_17392), .b(FE_OFN1241_n_4092), .c(g62492_sb), .o(n_6601) );
na03f40 TIMEBOOST_cell_41296 ( .a(n_2308), .b(n_3503), .c(n_15927), .o(TIMEBOOST_net_10377) );
na03f02 TIMEBOOST_cell_66774 ( .a(n_3890), .b(g63095_sb), .c(g63095_db), .o(n_5064) );
in01f01 g61751_u0 ( .a(FE_OFN2081_n_8176), .o(g61751_sb) );
na04f06 TIMEBOOST_cell_64350 ( .a(n_1252), .b(n_1340), .c(n_1354), .d(n_1342), .o(n_2402) );
na02m04 TIMEBOOST_cell_68758 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q), .b(FE_OFN660_n_4392), .o(TIMEBOOST_net_21587) );
na02m08 TIMEBOOST_cell_52875 ( .a(wbs_dat_i_18_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q), .o(TIMEBOOST_net_16655) );
in01s02 g61752_u0 ( .a(n_8272), .o(g61752_sb) );
na02f02 TIMEBOOST_cell_71110 ( .a(TIMEBOOST_net_17401), .b(FE_OFN1264_n_4095), .o(TIMEBOOST_net_22763) );
na02m01 TIMEBOOST_cell_68057 ( .a(TIMEBOOST_net_21236), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_389), .o(TIMEBOOST_net_16809) );
na02m02 TIMEBOOST_cell_70161 ( .a(TIMEBOOST_net_22288), .b(g64218_sb), .o(n_3951) );
in01m01 g61753_u0 ( .a(FE_OFN2257_n_8060), .o(g61753_sb) );
na02m02 TIMEBOOST_cell_69435 ( .a(TIMEBOOST_net_21925), .b(TIMEBOOST_net_16259), .o(TIMEBOOST_net_17150) );
na03f01 TIMEBOOST_cell_65072 ( .a(n_3774), .b(FE_OFN643_n_4677), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q), .o(TIMEBOOST_net_14512) );
in01s02 g61754_u0 ( .a(FE_OFN704_n_8069), .o(g61754_sb) );
na02s02 TIMEBOOST_cell_28179 ( .a(TIMEBOOST_net_21179), .b(g65697_sb), .o(TIMEBOOST_net_8194) );
na02f02 TIMEBOOST_cell_28253 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q), .b(g64354_sb), .o(TIMEBOOST_net_8231) );
na03f02 TIMEBOOST_cell_66815 ( .a(TIMEBOOST_net_16846), .b(FE_OFN1345_n_8567), .c(g57148_sb), .o(n_11602) );
in01s02 g61755_u0 ( .a(FE_OFN704_n_8069), .o(g61755_sb) );
na03f01 TIMEBOOST_cell_66775 ( .a(n_14967), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in_84), .c(n_14482), .o(TIMEBOOST_net_11920) );
in01m03 TIMEBOOST_cell_67728 ( .a(TIMEBOOST_net_21155), .o(TIMEBOOST_net_21154) );
in01m01 g61756_u0 ( .a(FE_OFN719_n_8060), .o(g61756_sb) );
na02m02 TIMEBOOST_cell_37970 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q), .b(g58388_sb), .o(TIMEBOOST_net_10597) );
na03m03 TIMEBOOST_cell_66264 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .b(n_4658), .c(n_7136), .o(n_7393) );
na02m02 TIMEBOOST_cell_62804 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_139), .o(TIMEBOOST_net_20349) );
in01m01 g61757_u0 ( .a(FE_OFN2257_n_8060), .o(g61757_sb) );
na02f02 TIMEBOOST_cell_42984 ( .a(TIMEBOOST_net_12386), .b(g58792_sb), .o(n_9828) );
in01f01 g61758_u0 ( .a(FE_OFN2084_n_8407), .o(g61758_sb) );
na03m04 TIMEBOOST_cell_72599 ( .a(TIMEBOOST_net_23153), .b(FE_OFN1660_n_4490), .c(TIMEBOOST_net_21728), .o(TIMEBOOST_net_13378) );
na02s01 TIMEBOOST_cell_43454 ( .a(TIMEBOOST_net_12621), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_10784) );
in01f02 g61759_u0 ( .a(FE_OFN717_n_8176), .o(g61759_sb) );
na02m01 TIMEBOOST_cell_48672 ( .a(TIMEBOOST_net_14553), .b(FE_OFN912_n_4727), .o(TIMEBOOST_net_12841) );
na02s01 TIMEBOOST_cell_43456 ( .a(TIMEBOOST_net_12622), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_10785) );
na02s01 TIMEBOOST_cell_43458 ( .a(TIMEBOOST_net_12623), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_10786) );
in01f01 g61760_u0 ( .a(FE_OFN2084_n_8407), .o(g61760_sb) );
na03f02 TIMEBOOST_cell_66453 ( .a(TIMEBOOST_net_17380), .b(FE_OFN1283_n_4097), .c(g62437_sb), .o(n_6722) );
na03m02 TIMEBOOST_cell_68924 ( .a(n_4493), .b(g65072_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q), .o(TIMEBOOST_net_21670) );
in01f01 g61761_u0 ( .a(FE_OFN714_n_8140), .o(g61761_sb) );
na02m02 TIMEBOOST_cell_69017 ( .a(TIMEBOOST_net_21716), .b(FE_OFN667_n_4495), .o(TIMEBOOST_net_16269) );
na03m02 TIMEBOOST_cell_68584 ( .a(TIMEBOOST_net_10280), .b(FE_OFN623_n_4409), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q), .o(TIMEBOOST_net_21500) );
in01s02 g61762_u0 ( .a(FE_OFN719_n_8060), .o(g61762_sb) );
na03f01 TIMEBOOST_cell_67972 ( .a(TIMEBOOST_net_15238), .b(FE_OFN1179_n_3476), .c(g60633_sb), .o(n_5703) );
na02m02 TIMEBOOST_cell_62498 ( .a(n_4677), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q), .o(TIMEBOOST_net_20196) );
in01s01 g61763_u0 ( .a(FE_OFN2256_n_8060), .o(g61763_sb) );
na02f01 TIMEBOOST_cell_47763 ( .a(pci_idsel_i), .b(FE_OFN989_n_574), .o(TIMEBOOST_net_14099) );
na03f02 TIMEBOOST_cell_66777 ( .a(TIMEBOOST_net_17060), .b(n_6319), .c(g62996_sb), .o(n_5890) );
na02f02 TIMEBOOST_cell_70081 ( .a(TIMEBOOST_net_22248), .b(g64864_db), .o(TIMEBOOST_net_8843) );
in01s01 g61764_u0 ( .a(n_8140), .o(g61764_sb) );
na02s01 g61764_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q), .b(n_8140), .o(g61764_db) );
in01s01 g61765_u0 ( .a(n_8119), .o(g61765_sb) );
in01s01 TIMEBOOST_cell_67712 ( .a(TIMEBOOST_net_21138), .o(TIMEBOOST_net_21139) );
na02s01 g61765_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q), .b(n_8119), .o(g61765_db) );
na03f02 TIMEBOOST_cell_73716 ( .a(TIMEBOOST_net_13550), .b(n_11977), .c(FE_OFN1746_n_12004), .o(n_12640) );
in01m01 g61766_u0 ( .a(FE_OFN2257_n_8060), .o(g61766_sb) );
na02s01 TIMEBOOST_cell_43462 ( .a(TIMEBOOST_net_12625), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_10788) );
in01s01 g61767_u0 ( .a(n_8119), .o(g61767_sb) );
na02m02 TIMEBOOST_cell_39593 ( .a(TIMEBOOST_net_11408), .b(g63431_sb), .o(n_4934) );
na02s01 g61767_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q), .b(n_8119), .o(g61767_db) );
in01s01 g61768_u0 ( .a(n_8272), .o(g61768_sb) );
na02m02 TIMEBOOST_cell_38752 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q), .b(g65856_sb), .o(TIMEBOOST_net_10988) );
in01f02 TIMEBOOST_cell_42692 ( .a(TIMEBOOST_net_12240), .o(TIMEBOOST_net_12239) );
in01f01 g61769_u0 ( .a(FE_OFN714_n_8140), .o(g61769_sb) );
no03f04 TIMEBOOST_cell_73684 ( .a(n_4647), .b(n_7552), .c(n_4881), .o(g59344_p) );
na03m06 TIMEBOOST_cell_70136 ( .a(FE_OFN1676_n_4655), .b(n_4444), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q), .o(TIMEBOOST_net_22276) );
na02s01 TIMEBOOST_cell_18060 ( .a(TIMEBOOST_net_5393), .b(g66398_sb), .o(n_2504) );
in01f01 g61770_u0 ( .a(FE_OFN707_n_8119), .o(g61770_sb) );
na03f04 TIMEBOOST_cell_73164 ( .a(TIMEBOOST_net_17281), .b(FE_OFN2128_n_16497), .c(g54332_sb), .o(n_12984) );
na02m08 TIMEBOOST_cell_52867 ( .a(wbs_dat_i_29_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q), .o(TIMEBOOST_net_16651) );
in01s01 g61771_u0 ( .a(n_8119), .o(g61771_sb) );
na02s01 TIMEBOOST_cell_47919 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q), .o(TIMEBOOST_net_14177) );
na02s01 g61771_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q), .b(n_8119), .o(g61771_db) );
na03f02 TIMEBOOST_cell_47305 ( .a(FE_OFN1554_n_12104), .b(FE_OCP_RBN1979_n_10273), .c(TIMEBOOST_net_13590), .o(n_12597) );
in01s01 g61772_u0 ( .a(n_8232), .o(g61772_sb) );
na02m02 TIMEBOOST_cell_38754 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q), .b(g65920_sb), .o(TIMEBOOST_net_10989) );
na02m01 g61772_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q), .b(n_8232), .o(g61772_db) );
na03m08 TIMEBOOST_cell_72196 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q), .b(FE_OFN1076_n_4740), .c(pci_target_unit_fifos_pciw_addr_data_in_135), .o(TIMEBOOST_net_23306) );
in01m01 g61773_u0 ( .a(FE_OFN699_n_7845), .o(g61773_sb) );
na03s02 TIMEBOOST_cell_72887 ( .a(g61870_sb), .b(g61870_db), .c(n_1854), .o(n_8094) );
na02f02 TIMEBOOST_cell_44568 ( .a(TIMEBOOST_net_13178), .b(g63075_sb), .o(n_5100) );
na03f02 TIMEBOOST_cell_66634 ( .a(TIMEBOOST_net_8543), .b(FE_OCPN1847_n_14981), .c(g59098_sb), .o(n_8695) );
in01s01 g61774_u0 ( .a(FE_OFN702_n_7845), .o(g61774_sb) );
na03f02 TIMEBOOST_cell_66540 ( .a(TIMEBOOST_net_17567), .b(FE_OFN1332_n_13547), .c(g53920_sb), .o(n_13524) );
na03m02 TIMEBOOST_cell_72787 ( .a(n_4672), .b(FE_OFN1640_n_4671), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q), .o(TIMEBOOST_net_23234) );
in01s01 g61775_u0 ( .a(n_8407), .o(g61775_sb) );
na03s01 TIMEBOOST_cell_72460 ( .a(n_2499), .b(FE_OFN2094_n_2520), .c(g66426_db), .o(n_2500) );
na02s01 g61775_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q), .b(n_8407), .o(g61775_db) );
na02f02 TIMEBOOST_cell_50436 ( .a(TIMEBOOST_net_15435), .b(g62934_sb), .o(n_6013) );
na02s01 g61776_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q), .b(n_7102), .o(g61776_db) );
na02f02 TIMEBOOST_cell_50434 ( .a(TIMEBOOST_net_15434), .b(g63173_sb), .o(n_5798) );
in01s01 g61777_u0 ( .a(n_8232), .o(g61777_sb) );
na02m02 TIMEBOOST_cell_72248 ( .a(n_3678), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q), .o(TIMEBOOST_net_23332) );
na02m01 g61777_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q), .b(n_8232), .o(g61777_db) );
in01m01 g61778_u0 ( .a(FE_OFN719_n_8060), .o(g61778_sb) );
in01s01 TIMEBOOST_cell_73885 ( .a(TIMEBOOST_net_23449), .o(TIMEBOOST_net_23450) );
no03f08 TIMEBOOST_cell_64318 ( .a(FE_RN_315_0), .b(FE_RN_317_0), .c(FE_RN_322_0), .o(FE_RN_323_0) );
in01s01 g61779_u0 ( .a(n_8119), .o(g61779_sb) );
na03m02 TIMEBOOST_cell_65118 ( .a(n_3774), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q), .c(FE_OFN1642_n_4671), .o(TIMEBOOST_net_14373) );
na02s01 g61779_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q), .b(n_8119), .o(g61779_db) );
na02m02 TIMEBOOST_cell_70693 ( .a(TIMEBOOST_net_22554), .b(g62800_sb), .o(n_5383) );
in01f01 g61780_u0 ( .a(FE_OFN2084_n_8407), .o(g61780_sb) );
na03f02 TIMEBOOST_cell_71436 ( .a(TIMEBOOST_net_11637), .b(n_7685), .c(TIMEBOOST_net_501), .o(TIMEBOOST_net_22926) );
na02f01 TIMEBOOST_cell_18042 ( .a(TIMEBOOST_net_5384), .b(n_2487), .o(TIMEBOOST_net_183) );
in01s01 g61781_u0 ( .a(n_8272), .o(g61781_sb) );
na04s01 TIMEBOOST_cell_67827 ( .a(g58058_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q), .c(g58058_db), .d(FE_OFN237_n_9118), .o(TIMEBOOST_net_9500) );
in01m01 g61782_u0 ( .a(FE_OFN720_n_8060), .o(g61782_sb) );
na02f02 TIMEBOOST_cell_63197 ( .a(TIMEBOOST_net_20545), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_15693) );
na02f02 TIMEBOOST_cell_70203 ( .a(TIMEBOOST_net_22309), .b(g54336_sb), .o(n_13098) );
na02s02 TIMEBOOST_cell_54546 ( .a(TIMEBOOST_net_17490), .b(TIMEBOOST_net_10889), .o(TIMEBOOST_net_9334) );
in01s01 g61783_u0 ( .a(n_8232), .o(g61783_sb) );
na02f01 TIMEBOOST_cell_38758 ( .a(conf_wb_err_addr_in_944), .b(g53939_sb), .o(TIMEBOOST_net_10991) );
na02s01 g61783_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q), .b(n_8232), .o(g61783_db) );
in01s01 TIMEBOOST_cell_73977 ( .a(TIMEBOOST_net_23541), .o(TIMEBOOST_net_23542) );
in01f01 g61784_u0 ( .a(FE_OFN713_n_8140), .o(g61784_sb) );
na02f01 TIMEBOOST_cell_69603 ( .a(TIMEBOOST_net_22009), .b(FE_OFN1033_n_4732), .o(TIMEBOOST_net_11166) );
na02m02 TIMEBOOST_cell_49132 ( .a(TIMEBOOST_net_14783), .b(g61799_sb), .o(n_8198) );
na03f02 TIMEBOOST_cell_73816 ( .a(TIMEBOOST_net_13780), .b(FE_OFN1773_n_13800), .c(FE_OFN1769_n_14054), .o(n_14462) );
in01m01 g61785_u0 ( .a(FE_OFN709_n_8232), .o(g61785_sb) );
na03f02 TIMEBOOST_cell_35044 ( .a(TIMEBOOST_net_9588), .b(FE_OFN1441_n_9372), .c(g58465_sb), .o(n_9385) );
na03f02 TIMEBOOST_cell_67027 ( .a(FE_OFN1606_n_13997), .b(TIMEBOOST_net_13755), .c(FE_OFN1599_n_13995), .o(n_14474) );
in01f01 g61786_u0 ( .a(FE_OFN2081_n_8176), .o(g61786_sb) );
na04s04 TIMEBOOST_cell_73337 ( .a(FE_OFN600_n_9687), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q), .c(FE_OFN219_n_9853), .d(g58114_sb), .o(n_9680) );
na02s01 TIMEBOOST_cell_38413 ( .a(TIMEBOOST_net_10818), .b(g57958_db), .o(n_9847) );
in01f01 g61787_u0 ( .a(FE_OFN706_n_8119), .o(g61787_sb) );
na03f02 TIMEBOOST_cell_35046 ( .a(TIMEBOOST_net_9596), .b(FE_OFN1441_n_9372), .c(g58458_sb), .o(n_8989) );
na02f02 TIMEBOOST_cell_70985 ( .a(TIMEBOOST_net_22700), .b(g62657_sb), .o(n_6230) );
in01f01 g61788_u0 ( .a(FE_OFN2084_n_8407), .o(g61788_sb) );
na03f02 TIMEBOOST_cell_34862 ( .a(TIMEBOOST_net_9413), .b(FE_OFN1392_n_8567), .c(g57057_sb), .o(n_11680) );
na02s01 TIMEBOOST_cell_52415 ( .a(g57900_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q), .o(TIMEBOOST_net_16425) );
in01f01 g61789_u0 ( .a(FE_OFN707_n_8119), .o(g61789_sb) );
na03m02 TIMEBOOST_cell_72855 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q), .b(g65432_sb), .c(TIMEBOOST_net_23234), .o(TIMEBOOST_net_15339) );
na03m08 TIMEBOOST_cell_69076 ( .a(FE_OFN653_n_4508), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q), .c(n_4493), .o(TIMEBOOST_net_21746) );
na02f02 TIMEBOOST_cell_54225 ( .a(n_4057), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q), .o(TIMEBOOST_net_17330) );
in01f01 g61790_u0 ( .a(FE_OFN706_n_8119), .o(g61790_sb) );
na02f01 TIMEBOOST_cell_54226 ( .a(TIMEBOOST_net_17330), .b(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_15163) );
na04f04 TIMEBOOST_cell_67698 ( .a(TIMEBOOST_net_16855), .b(FE_OFN2198_n_10256), .c(g52620_sb), .d(TIMEBOOST_net_699), .o(n_11850) );
in01s01 g61791_u0 ( .a(FE_OFN2257_n_8060), .o(g61791_sb) );
na03m04 TIMEBOOST_cell_73135 ( .a(FE_OFN1076_n_4740), .b(TIMEBOOST_net_16351), .c(g64103_sb), .o(n_4053) );
in01f01 g61792_u0 ( .a(FE_OFN717_n_8176), .o(g61792_sb) );
na03m02 TIMEBOOST_cell_49171 ( .a(n_1920), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q), .c(FE_OFN702_n_7845), .o(TIMEBOOST_net_14803) );
na03f02 TIMEBOOST_cell_66892 ( .a(FE_OFN1746_n_12004), .b(TIMEBOOST_net_16001), .c(n_11977), .o(n_12646) );
na04f04 TIMEBOOST_cell_73439 ( .a(n_3655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q), .c(FE_OFN1249_n_4093), .d(g62531_sb), .o(n_6512) );
in01f01 g61793_u0 ( .a(FE_OFN2081_n_8176), .o(g61793_sb) );
na02m01 TIMEBOOST_cell_43027 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_12408) );
na02s01 TIMEBOOST_cell_48163 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q), .o(TIMEBOOST_net_14299) );
in01f01 g61794_u0 ( .a(FE_OFN716_n_8176), .o(g61794_sb) );
na03f02 TIMEBOOST_cell_66890 ( .a(FE_OFN1749_n_12004), .b(n_12010), .c(TIMEBOOST_net_13557), .o(n_12765) );
na03m01 TIMEBOOST_cell_64422 ( .a(TIMEBOOST_net_20795), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_405), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q), .o(TIMEBOOST_net_16797) );
na03m02 TIMEBOOST_cell_48121 ( .a(n_3761), .b(FE_OFN667_n_4495), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q), .o(TIMEBOOST_net_14278) );
in01f02 g61795_u0 ( .a(FE_OFN710_n_8232), .o(g61795_sb) );
na03f02 TIMEBOOST_cell_34926 ( .a(TIMEBOOST_net_9564), .b(FE_OFN1401_n_8567), .c(g57398_sb), .o(n_10372) );
na02m02 TIMEBOOST_cell_69052 ( .a(g65311_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q), .o(TIMEBOOST_net_21734) );
in01s01 g61796_u0 ( .a(n_8176), .o(g61796_sb) );
na03f02 TIMEBOOST_cell_67029 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_16533), .c(FE_OFN1601_n_13995), .o(n_16210) );
na02s01 g61796_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q), .b(n_8176), .o(g61796_db) );
na03f02 TIMEBOOST_cell_73779 ( .a(n_13993), .b(TIMEBOOST_net_13719), .c(FE_OFN1588_n_13736), .o(n_14293) );
in01s01 g61797_u0 ( .a(n_8140), .o(g61797_sb) );
na02f02 TIMEBOOST_cell_72255 ( .a(TIMEBOOST_net_23335), .b(g60659_sb), .o(n_5662) );
na02s01 g61797_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q), .b(n_8140), .o(g61797_db) );
in01s01 TIMEBOOST_cell_73842 ( .a(n_13757), .o(TIMEBOOST_net_23407) );
in01s01 g61798_u0 ( .a(n_8232), .o(g61798_sb) );
na02s01 TIMEBOOST_cell_45393 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q), .o(TIMEBOOST_net_13591) );
na02s01 g61798_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q), .b(n_8232), .o(g61798_db) );
na02m04 TIMEBOOST_cell_62472 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_136), .o(TIMEBOOST_net_20183) );
in01s01 g61799_u0 ( .a(FE_OFN701_n_7845), .o(g61799_sb) );
na02f01 TIMEBOOST_cell_62990 ( .a(conf_wb_err_addr_in_959), .b(g62119_sb), .o(TIMEBOOST_net_20442) );
na02m02 TIMEBOOST_cell_50695 ( .a(n_4900), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q), .o(TIMEBOOST_net_15565) );
na03m02 TIMEBOOST_cell_68590 ( .a(FE_OFN624_n_4409), .b(g64899_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q), .o(TIMEBOOST_net_21503) );
in01s01 g61800_u0 ( .a(FE_OFN699_n_7845), .o(g61800_sb) );
in01s01 g61801_u0 ( .a(n_8069), .o(g61801_sb) );
na02s04 TIMEBOOST_cell_64080 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_21026) );
na02s01 g61801_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q), .b(n_8069), .o(g61801_db) );
na03f02 TIMEBOOST_cell_47289 ( .a(FE_OFN1736_n_16317), .b(TIMEBOOST_net_13585), .c(FE_OFN1742_n_11019), .o(n_12701) );
in01m01 g61802_u0 ( .a(FE_OFN716_n_8176), .o(g61802_sb) );
na03f02 TIMEBOOST_cell_35048 ( .a(TIMEBOOST_net_9598), .b(FE_OFN1440_n_9372), .c(g58484_sb), .o(n_9353) );
na02s01 TIMEBOOST_cell_68184 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q), .o(TIMEBOOST_net_21300) );
na02f01 TIMEBOOST_cell_69110 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(g64160_sb), .o(TIMEBOOST_net_21763) );
in01f01 g61803_u0 ( .a(FE_OFN714_n_8140), .o(g61803_sb) );
na02s02 TIMEBOOST_cell_38566 ( .a(g57912_sb), .b(FE_OFN252_n_9868), .o(TIMEBOOST_net_10895) );
na02f02 TIMEBOOST_cell_28010 ( .a(n_13901), .b(TIMEBOOST_net_8109), .o(TIMEBOOST_net_760) );
in01s01 g61804_u0 ( .a(n_8140), .o(g61804_sb) );
na02s01 g61804_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q), .b(n_8140), .o(g61804_db) );
na03f01 TIMEBOOST_cell_624 ( .a(n_4014), .b(g62808_sb), .c(g62808_db), .o(n_5363) );
in01f01 g61805_u0 ( .a(FE_OFN714_n_8140), .o(g61805_sb) );
na02s01 TIMEBOOST_cell_38568 ( .a(FE_OFN215_n_9856), .b(g58112_sb), .o(TIMEBOOST_net_10896) );
na02f02 TIMEBOOST_cell_38981 ( .a(TIMEBOOST_net_11102), .b(FE_OFN1151_n_13249), .o(TIMEBOOST_net_360) );
na03f02 TIMEBOOST_cell_65682 ( .a(pci_target_unit_pcit_if_strd_addr_in_710), .b(g52639_sb), .c(TIMEBOOST_net_14913), .o(n_14751) );
in01f01 g61806_u0 ( .a(FE_OFN714_n_8140), .o(g61806_sb) );
na02s01 TIMEBOOST_cell_38570 ( .a(g58044_sb), .b(FE_OFN213_n_9124), .o(TIMEBOOST_net_10897) );
na02s01 TIMEBOOST_cell_39127 ( .a(TIMEBOOST_net_11175), .b(g58420_sb), .o(n_9427) );
in01s01 g61807_u0 ( .a(n_8272), .o(g61807_sb) );
na02m10 TIMEBOOST_cell_52803 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_136), .o(TIMEBOOST_net_16619) );
na02s02 TIMEBOOST_cell_49463 ( .a(FE_OFN260_n_9860), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q), .o(TIMEBOOST_net_14949) );
na02s06 TIMEBOOST_cell_18002 ( .a(TIMEBOOST_net_5364), .b(g58798_db), .o(n_9825) );
in01s01 g61808_u0 ( .a(n_8176), .o(g61808_sb) );
na02m04 TIMEBOOST_cell_68540 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q), .o(TIMEBOOST_net_21478) );
na02s01 g61808_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q), .b(n_8176), .o(g61808_db) );
na02m02 TIMEBOOST_cell_68887 ( .a(TIMEBOOST_net_21651), .b(TIMEBOOST_net_14245), .o(TIMEBOOST_net_17447) );
in01m01 g61809_u0 ( .a(FE_OFN2258_n_8060), .o(g61809_sb) );
na03f02 TIMEBOOST_cell_73146 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q), .b(FE_OFN1075_n_4740), .c(TIMEBOOST_net_22295), .o(TIMEBOOST_net_8807) );
na02m02 TIMEBOOST_cell_49230 ( .a(g65882_db), .b(TIMEBOOST_net_14832), .o(n_1864) );
na04f04 TIMEBOOST_cell_24159 ( .a(n_8548), .b(g58608_sb), .c(n_317), .d(FE_OFN1403_n_8567), .o(n_8899) );
in01s01 g61810_u0 ( .a(n_8069), .o(g61810_sb) );
na02s02 TIMEBOOST_cell_18001 ( .a(g58798_sb), .b(wbu_addr_in_258), .o(TIMEBOOST_net_5364) );
na02s01 g61810_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q), .b(n_8069), .o(g61810_db) );
na02m04 TIMEBOOST_cell_53845 ( .a(n_4232), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q), .o(TIMEBOOST_net_17140) );
in01f01 g61811_u0 ( .a(FE_OFN716_n_8176), .o(g61811_sb) );
na02s01 TIMEBOOST_cell_38572 ( .a(g58010_sb), .b(FE_OFN254_n_9825), .o(TIMEBOOST_net_10898) );
na03f02 TIMEBOOST_cell_65169 ( .a(TIMEBOOST_net_14443), .b(g64198_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q), .o(TIMEBOOST_net_13090) );
in01s01 g61812_u0 ( .a(n_8176), .o(g61812_sb) );
na02s01 TIMEBOOST_cell_31009 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_16__Q), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_9609) );
na02s01 g61812_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q), .b(n_8176), .o(g61812_db) );
in01s01 TIMEBOOST_cell_63594 ( .a(TIMEBOOST_net_20774), .o(TIMEBOOST_net_20751) );
in01f01 g61813_u0 ( .a(FE_OFN710_n_8232), .o(g61813_sb) );
na02s01 TIMEBOOST_cell_38574 ( .a(g58142_sb), .b(FE_OFN211_n_9858), .o(TIMEBOOST_net_10899) );
in01m08 TIMEBOOST_cell_35517 ( .a(TIMEBOOST_net_10107), .o(TIMEBOOST_net_10108) );
no02f02 TIMEBOOST_cell_51373 ( .a(TIMEBOOST_net_5383), .b(FE_RN_619_0), .o(TIMEBOOST_net_15904) );
in01f01 g61814_u0 ( .a(FE_OFN709_n_8232), .o(g61814_sb) );
na02s01 TIMEBOOST_cell_43133 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q), .o(TIMEBOOST_net_12461) );
na03m02 TIMEBOOST_cell_64537 ( .a(n_3749), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q), .c(FE_OFN687_n_4417), .o(TIMEBOOST_net_16597) );
in01m02 g61815_u0 ( .a(FE_OFN720_n_8060), .o(g61815_sb) );
na04m02 TIMEBOOST_cell_65049 ( .a(TIMEBOOST_net_10456), .b(g64846_sb), .c(n_4476), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_17392) );
na02m06 TIMEBOOST_cell_38290 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q), .b(g65285_sb), .o(TIMEBOOST_net_10757) );
in01f01 g61816_u0 ( .a(FE_OFN706_n_8119), .o(g61816_sb) );
na03m06 TIMEBOOST_cell_72002 ( .a(FE_OFN930_n_4730), .b(TIMEBOOST_net_14258), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_23209) );
na02m01 g61816_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q), .b(n_8119), .o(g61816_db) );
na03m02 TIMEBOOST_cell_65066 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q), .b(n_3785), .c(FE_OFN625_n_4409), .o(TIMEBOOST_net_10638) );
in01f01 g61817_u0 ( .a(FE_OFN1812_n_7845), .o(g61817_sb) );
na03m02 TIMEBOOST_cell_64536 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q), .b(n_3755), .c(FE_OFN687_n_4417), .o(TIMEBOOST_net_10445) );
na02m01 TIMEBOOST_cell_71850 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q), .b(n_3764), .o(TIMEBOOST_net_23133) );
in01s01 g61818_u0 ( .a(FE_OFN701_n_7845), .o(g61818_sb) );
na04f04 TIMEBOOST_cell_36821 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q), .b(FE_OFN1379_n_8567), .c(n_9004), .d(g57543_sb), .o(n_10310) );
na03m02 TIMEBOOST_cell_70154 ( .a(FE_OFN1077_n_4740), .b(pci_target_unit_fifos_pciw_addr_data_in_130), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q), .o(TIMEBOOST_net_22285) );
na03f02 TIMEBOOST_cell_35050 ( .a(TIMEBOOST_net_9602), .b(FE_OFN1440_n_9372), .c(g58483_sb), .o(n_8973) );
in01f01 g61819_u0 ( .a(FE_OFN2084_n_8407), .o(g61819_sb) );
na02m01 TIMEBOOST_cell_43031 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_124), .o(TIMEBOOST_net_12410) );
na03m02 TIMEBOOST_cell_68978 ( .a(FE_OFN908_n_4734), .b(pci_target_unit_fifos_pciw_addr_data_in_128), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q), .o(TIMEBOOST_net_21697) );
na03f02 TIMEBOOST_cell_66274 ( .a(wbm_dat_o_5_), .b(g60666_sb), .c(TIMEBOOST_net_7601), .o(n_5652) );
in01s01 g61820_u0 ( .a(n_8140), .o(g61820_sb) );
na02s01 g61820_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q), .b(n_8140), .o(g61820_db) );
na02m02 TIMEBOOST_cell_68585 ( .a(TIMEBOOST_net_21500), .b(g65673_sb), .o(TIMEBOOST_net_17419) );
in01f01 g61821_u0 ( .a(FE_OFN2081_n_8176), .o(g61821_sb) );
na03f02 TIMEBOOST_cell_67973 ( .a(TIMEBOOST_net_8838), .b(FE_OFN1183_n_3476), .c(g60651_sb), .o(n_5673) );
na02m10 TIMEBOOST_cell_48081 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_141), .o(TIMEBOOST_net_14258) );
na02f02 TIMEBOOST_cell_50944 ( .a(TIMEBOOST_net_15689), .b(g62340_sb), .o(n_6919) );
in01f01 g61822_u0 ( .a(FE_OFN2212_n_8407), .o(g61822_sb) );
na04m02 TIMEBOOST_cell_67897 ( .a(n_3752), .b(FE_OFN1677_n_4655), .c(g65353_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q), .o(TIMEBOOST_net_7592) );
na02m01 TIMEBOOST_cell_68207 ( .a(TIMEBOOST_net_21311), .b(g57795_sb), .o(TIMEBOOST_net_17588) );
na03m02 TIMEBOOST_cell_71992 ( .a(g64979_sb), .b(n_4476), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q), .o(TIMEBOOST_net_23204) );
in01f01 g61823_u0 ( .a(FE_OFN712_n_8140), .o(g61823_sb) );
na02m06 TIMEBOOST_cell_52783 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_133), .o(TIMEBOOST_net_16609) );
na03m02 TIMEBOOST_cell_72332 ( .a(TIMEBOOST_net_20606), .b(FE_OFN1689_n_9528), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q), .o(TIMEBOOST_net_23374) );
in01f01 g61824_u0 ( .a(FE_OFN712_n_8140), .o(g61824_sb) );
na04m06 TIMEBOOST_cell_72500 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q), .b(n_3752), .c(FE_OFN670_n_4505), .d(TIMEBOOST_net_21442), .o(TIMEBOOST_net_17503) );
in01s01 TIMEBOOST_cell_73886 ( .a(n_8316), .o(TIMEBOOST_net_23451) );
na04f04 TIMEBOOST_cell_24158 ( .a(n_8558), .b(g58590_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q), .d(FE_OFN1403_n_8567), .o(n_8910) );
in01f01 g61825_u0 ( .a(FE_OFN2212_n_8407), .o(g61825_sb) );
na04f04 TIMEBOOST_cell_67400 ( .a(g61945_sb), .b(FE_OFN2257_n_8060), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q), .d(n_1582), .o(n_7935) );
na03f02 TIMEBOOST_cell_65958 ( .a(TIMEBOOST_net_20896), .b(FE_OFN1174_n_5592), .c(g62074_sb), .o(n_5637) );
in01f01 g61826_u0 ( .a(FE_OFN2084_n_8407), .o(g61826_sb) );
na02m02 TIMEBOOST_cell_44846 ( .a(TIMEBOOST_net_13317), .b(g60630_sb), .o(n_5707) );
na02f01 TIMEBOOST_cell_18303 ( .a(configuration_pci_err_addr_479), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_5515) );
in01m01 g61827_u0 ( .a(FE_OFN719_n_8060), .o(g61827_sb) );
na02f06 FE_RC_885_0 ( .a(FE_RN_579_0), .b(FE_RN_580_0), .o(FE_RN_581_0) );
in01f01 g61828_u0 ( .a(FE_OFN1812_n_7845), .o(g61828_sb) );
na02s01 TIMEBOOST_cell_43457 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q), .o(TIMEBOOST_net_12623) );
in01m01 g61829_u0 ( .a(FE_OFN720_n_8060), .o(g61829_sb) );
na02f02 TIMEBOOST_cell_70760 ( .a(wbm_adr_o_7_), .b(g63577_sb), .o(TIMEBOOST_net_22588) );
na04f04 TIMEBOOST_cell_24160 ( .a(n_1287), .b(g58576_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .d(FE_OFN1369_n_8567), .o(n_9192) );
na03f02 TIMEBOOST_cell_73382 ( .a(TIMEBOOST_net_16720), .b(FE_OFN1301_n_5763), .c(g62056_sb), .o(n_7753) );
in01m01 g61830_u0 ( .a(FE_OFN701_n_7845), .o(g61830_sb) );
na02s01 TIMEBOOST_cell_43099 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_12444) );
na03m02 TIMEBOOST_cell_64535 ( .a(n_3755), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q), .c(FE_OFN634_n_4454), .o(TIMEBOOST_net_10401) );
na02m04 TIMEBOOST_cell_72330 ( .a(g65304_sb), .b(n_15), .o(TIMEBOOST_net_23373) );
na02s02 TIMEBOOST_cell_43759 ( .a(FE_OFN233_n_9876), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q), .o(TIMEBOOST_net_12774) );
na02f02 TIMEBOOST_cell_70695 ( .a(TIMEBOOST_net_22555), .b(g62854_sb), .o(n_5260) );
no02f04 g61832_u0 ( .a(n_2942), .b(wbm_adr_o_28_), .o(g61832_p) );
ao12f02 g61832_u1 ( .a(g61832_p), .b(wbm_adr_o_28_), .c(n_2942), .o(n_3472) );
no02f06 g61833_u0 ( .a(wbu_addr_in_277), .b(n_2947), .o(g61833_p) );
ao12f04 g61833_u1 ( .a(g61833_p), .b(wbu_addr_in_277), .c(n_2947), .o(n_3471) );
no02f01 g61834_u0 ( .a(n_539), .b(n_3142), .o(g61834_p) );
ao12f01 g61834_u1 ( .a(g61834_p), .b(n_539), .c(n_3142), .o(n_4196) );
in01m02 g61835_u0 ( .a(FE_OFN1118_g64577_p), .o(g61835_sb) );
na02f08 TIMEBOOST_cell_71386 ( .a(TIMEBOOST_net_11794), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_22901) );
na03f02 TIMEBOOST_cell_42232 ( .a(TIMEBOOST_net_11487), .b(g58395_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q), .o(TIMEBOOST_net_9579) );
in01f01 g61836_u0 ( .a(FE_OFN1095_g64577_p), .o(g61836_sb) );
na03m02 TIMEBOOST_cell_64534 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q), .b(n_3792), .c(FE_OFN648_n_4497), .o(TIMEBOOST_net_10725) );
na02m02 TIMEBOOST_cell_38296 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q), .b(g65424_sb), .o(TIMEBOOST_net_10760) );
in01s01 g61837_u0 ( .a(FE_OFN1097_g64577_p), .o(g61837_sb) );
na02m01 g61837_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q), .b(FE_OFN1097_g64577_p), .o(g61837_db) );
no02f04 g61838_u0 ( .a(n_3318), .b(wbm_adr_o_31_), .o(g61838_p) );
ao12f02 g61838_u1 ( .a(g61838_p), .b(wbm_adr_o_31_), .c(n_3318), .o(n_4688) );
no02f04 g61839_u0 ( .a(conf_wb_err_addr_in_969), .b(FE_OFN2074_n_2723), .o(g61839_p) );
ao12f02 g61839_u1 ( .a(g61839_p), .b(conf_wb_err_addr_in_969), .c(FE_OFN2074_n_2723), .o(n_3344) );
in01f01 g61840_u0 ( .a(FE_OFN1094_g64577_p), .o(g61840_sb) );
na02f02 TIMEBOOST_cell_70536 ( .a(TIMEBOOST_net_13057), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_22476) );
na03f02 TIMEBOOST_cell_66712 ( .a(TIMEBOOST_net_16776), .b(FE_OFN1317_n_6624), .c(g63004_sb), .o(n_5874) );
in01f01 g61841_u0 ( .a(FE_OFN1094_g64577_p), .o(g61841_sb) );
na02m02 TIMEBOOST_cell_38298 ( .a(FE_RN_720_0), .b(g65435_sb), .o(TIMEBOOST_net_10761) );
na03f02 TIMEBOOST_cell_72078 ( .a(TIMEBOOST_net_12676), .b(FE_OFN1056_n_4727), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_23247) );
in01f01 g61842_u0 ( .a(FE_OFN1095_g64577_p), .o(g61842_sb) );
na03s01 TIMEBOOST_cell_64417 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q), .b(g65861_sb), .c(g65961_db), .o(n_2161) );
na03f02 TIMEBOOST_cell_66344 ( .a(TIMEBOOST_net_17524), .b(FE_OFN1234_n_6391), .c(g62409_sb), .o(n_6781) );
in01s01 TIMEBOOST_cell_63568 ( .a(TIMEBOOST_net_20748), .o(wbs_adr_i_15_) );
in01f02 g61843_u0 ( .a(n_13825), .o(g61843_sb) );
na03f02 TIMEBOOST_cell_73460 ( .a(TIMEBOOST_net_20522), .b(FE_OFN1289_n_4098), .c(g62637_sb), .o(n_6276) );
na02f06 TIMEBOOST_cell_18463 ( .a(n_16205), .b(FE_OCP_RBN2016_n_16970), .o(TIMEBOOST_net_5595) );
na02f02 TIMEBOOST_cell_49192 ( .a(TIMEBOOST_net_14813), .b(g61906_sb), .o(n_8009) );
no02f01 g61846_u0 ( .a(conf_wb_err_addr_in_950), .b(n_2011), .o(g61846_p) );
ao12f01 g61846_u1 ( .a(g61846_p), .b(conf_wb_err_addr_in_950), .c(n_2011), .o(n_2981) );
in01s01 g61847_u0 ( .a(n_7210), .o(n_7211) );
ao22f02 g61849_u0 ( .a(n_3429), .b(n_1041), .c(n_21), .d(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_4818) );
no02f02 g61850_u0 ( .a(wbu_addr_in_258), .b(n_2680), .o(g61850_p) );
ao12f02 g61850_u1 ( .a(g61850_p), .b(wbu_addr_in_258), .c(n_2680), .o(n_2740) );
no02f01 g61851_u0 ( .a(wbm_adr_o_9_), .b(n_2738), .o(g61851_p) );
ao12f01 g61851_u1 ( .a(g61851_p), .b(wbm_adr_o_9_), .c(n_2738), .o(n_2739) );
na02s02 TIMEBOOST_cell_48010 ( .a(TIMEBOOST_net_14222), .b(FE_OFN229_n_9120), .o(TIMEBOOST_net_10775) );
oa12f02 g61853_u0 ( .a(n_7733), .b(FE_OFN2079_n_8069), .c(n_8876), .o(n_8501) );
oa22f06 g61854_u0 ( .a(n_5763), .b(n_16763), .c(wishbone_slave_unit_pci_initiator_if_write_req_int), .d(n_2354), .o(n_13547) );
in01f02 g61855_u0 ( .a(FE_OFN1699_n_5751), .o(g61855_sb) );
in01s01 TIMEBOOST_cell_45875 ( .a(conf_wb_err_addr_in_958), .o(TIMEBOOST_net_13836) );
na02f02 g61855_u2 ( .a(n_3137), .b(FE_OFN1699_n_5751), .o(g61855_db) );
in01s01 TIMEBOOST_cell_67771 ( .a(pci_target_unit_fifos_pcir_data_in_169), .o(TIMEBOOST_net_21198) );
in01f02 g61856_u0 ( .a(FE_OFN1700_n_5751), .o(g61856_sb) );
in01s01 TIMEBOOST_cell_45876 ( .a(TIMEBOOST_net_13836), .o(TIMEBOOST_net_13837) );
na02f02 TIMEBOOST_cell_3453 ( .a(TIMEBOOST_net_286), .b(n_3132), .o(n_3142) );
no02f02 g61857_u0 ( .a(n_1273), .b(pci_target_unit_wishbone_master_rty_counter_4_), .o(g61857_p) );
ao12f02 g61857_u1 ( .a(g61857_p), .b(pci_target_unit_wishbone_master_rty_counter_4_), .c(n_1273), .o(n_2289) );
in01s01 g61858_u0 ( .a(n_8140), .o(g61858_sb) );
na02s01 TIMEBOOST_cell_47757 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q), .o(TIMEBOOST_net_14096) );
na02s01 g61858_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q), .b(n_8140), .o(g61858_db) );
in01s01 TIMEBOOST_cell_45969 ( .a(pci_target_unit_fifos_pcir_data_in_173), .o(TIMEBOOST_net_13930) );
in01s01 g61859_u0 ( .a(n_8119), .o(g61859_sb) );
na03f02 TIMEBOOST_cell_73803 ( .a(FE_OFN1775_n_13800), .b(TIMEBOOST_net_13783), .c(FE_OFN1769_n_14054), .o(n_14495) );
na02m01 g61859_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q), .b(n_8119), .o(g61859_db) );
na03m02 TIMEBOOST_cell_65119 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q), .b(n_3777), .c(FE_OFN1624_n_4438), .o(TIMEBOOST_net_16274) );
in01m01 g61860_u0 ( .a(FE_OFN719_n_8060), .o(g61860_sb) );
in01s01 TIMEBOOST_cell_73843 ( .a(TIMEBOOST_net_23407), .o(TIMEBOOST_net_23408) );
in01s01 g61861_u0 ( .a(FE_OFN702_n_7845), .o(g61861_sb) );
no02s01 TIMEBOOST_cell_28987 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237), .b(FE_RN_246_0), .o(TIMEBOOST_net_8598) );
na03f02 TIMEBOOST_cell_73658 ( .a(TIMEBOOST_net_14892), .b(FE_OFN1094_g64577_p), .c(g61955_sb), .o(n_6963) );
na02m02 TIMEBOOST_cell_18299 ( .a(pci_target_unit_wbm_sm_pciw_fifo_cbe_in), .b(n_8757), .o(TIMEBOOST_net_5513) );
in01s01 g61862_u0 ( .a(FE_OFN699_n_7845), .o(g61862_sb) );
na02m02 TIMEBOOST_cell_29001 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q), .o(TIMEBOOST_net_8605) );
na03f02 TIMEBOOST_cell_73749 ( .a(TIMEBOOST_net_16496), .b(FE_OFN1513_n_14987), .c(FE_OFN1554_n_12104), .o(FE_RN_908_0) );
na02f02 TIMEBOOST_cell_70416 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_22416) );
in01m01 g61863_u0 ( .a(n_8119), .o(g61863_sb) );
na02m01 g61863_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q), .b(n_8119), .o(g61863_db) );
na02m01 TIMEBOOST_cell_69418 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q), .b(FE_OFN647_n_4497), .o(TIMEBOOST_net_21917) );
in01m01 g61864_u0 ( .a(n_8119), .o(g61864_sb) );
na02f02 TIMEBOOST_cell_71655 ( .a(TIMEBOOST_net_23035), .b(FE_OFN1757_n_12681), .o(n_12524) );
na02m01 g61864_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q), .b(n_8119), .o(g61864_db) );
in01s01 g61865_u0 ( .a(n_8272), .o(g61865_sb) );
in01s01 TIMEBOOST_cell_35491 ( .a(TIMEBOOST_net_10082), .o(TIMEBOOST_net_10081) );
na03f02 TIMEBOOST_cell_66374 ( .a(TIMEBOOST_net_17083), .b(FE_OFN2064_n_6391), .c(g62469_sb), .o(n_6654) );
na02m10 TIMEBOOST_cell_45311 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q), .o(TIMEBOOST_net_13550) );
in01m01 g61866_u0 ( .a(n_8407), .o(g61866_sb) );
na02f01 TIMEBOOST_cell_18281 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_5504) );
na02m01 g61866_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q), .b(n_8407), .o(g61866_db) );
na03s01 TIMEBOOST_cell_72459 ( .a(pci_target_unit_del_sync_addr_in_228), .b(g66412_db), .c(g66399_sb), .o(n_2522) );
in01f01 g61867_u0 ( .a(FE_OFN712_n_8140), .o(g61867_sb) );
na02s02 TIMEBOOST_cell_28263 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(g65741_sb), .o(TIMEBOOST_net_8236) );
na03f02 TIMEBOOST_cell_67031 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_16530), .c(FE_OFN1600_n_13995), .o(n_16256) );
in01s01 g61868_u0 ( .a(n_8069), .o(g61868_sb) );
in01s01 TIMEBOOST_cell_73887 ( .a(TIMEBOOST_net_23451), .o(TIMEBOOST_net_23452) );
na04f04 TIMEBOOST_cell_73073 ( .a(n_1865), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q), .c(FE_OFN710_n_8232), .d(g61883_sb), .o(n_8064) );
na03f02 TIMEBOOST_cell_73575 ( .a(TIMEBOOST_net_20537), .b(FE_OFN1200_n_4090), .c(g62617_sb), .o(n_6323) );
in01f01 g61869_u0 ( .a(FE_OFN714_n_8140), .o(g61869_sb) );
na02f02 TIMEBOOST_cell_50348 ( .a(TIMEBOOST_net_15391), .b(g62943_sb), .o(n_5995) );
na03f02 TIMEBOOST_cell_73804 ( .a(TIMEBOOST_net_16552), .b(FE_OFN1773_n_13800), .c(FE_OFN1769_n_14054), .o(g53289_p) );
in01m01 g61870_u0 ( .a(n_8407), .o(g61870_sb) );
na03f02 TIMEBOOST_cell_66456 ( .a(TIMEBOOST_net_17117), .b(FE_OFN1310_n_6624), .c(g62501_sb), .o(n_6580) );
na02m01 g61870_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q), .b(n_8407), .o(g61870_db) );
na02s01 TIMEBOOST_cell_49486 ( .a(TIMEBOOST_net_14960), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9556) );
in01f01 g61871_u0 ( .a(FE_OFN713_n_8140), .o(g61871_sb) );
na02f01 TIMEBOOST_cell_28869 ( .a(n_1678), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .o(TIMEBOOST_net_8539) );
na02s01 TIMEBOOST_cell_47704 ( .a(TIMEBOOST_net_14069), .b(FE_OFN2094_n_2520), .o(n_2516) );
na02m02 TIMEBOOST_cell_63328 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q), .b(n_4906), .o(TIMEBOOST_net_20611) );
in01f01 g61872_u0 ( .a(FE_OFN716_n_8176), .o(g61872_sb) );
na02s01 TIMEBOOST_cell_28871 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_), .b(n_669), .o(TIMEBOOST_net_8540) );
na02f02 TIMEBOOST_cell_72229 ( .a(TIMEBOOST_net_23322), .b(g58351_sb), .o(TIMEBOOST_net_9443) );
na02m02 TIMEBOOST_cell_70149 ( .a(TIMEBOOST_net_22282), .b(g64170_sb), .o(n_3995) );
in01m01 g61873_u0 ( .a(FE_OFN701_n_7845), .o(g61873_sb) );
na02m20 TIMEBOOST_cell_52493 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59), .b(pci_target_unit_pcit_if_strd_addr_in_695), .o(TIMEBOOST_net_16464) );
in01f01 g61874_u0 ( .a(FE_OFN717_n_8176), .o(g61874_sb) );
na02s01 TIMEBOOST_cell_28873 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_), .o(TIMEBOOST_net_8541) );
na02m01 TIMEBOOST_cell_62451 ( .a(TIMEBOOST_net_20172), .b(FE_OFN906_n_4736), .o(TIMEBOOST_net_14136) );
na03f02 TIMEBOOST_cell_66071 ( .a(n_4074), .b(g62825_sb), .c(TIMEBOOST_net_7519), .o(n_5327) );
in01f02 g61875_u0 ( .a(FE_OFN706_n_8119), .o(g61875_sb) );
na03s02 TIMEBOOST_cell_68678 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q), .b(TIMEBOOST_net_14191), .c(FE_OFN953_n_2055), .o(TIMEBOOST_net_21547) );
na03s01 TIMEBOOST_cell_72445 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q), .b(g65870_sb), .c(g65870_db), .o(n_2300) );
na03m02 TIMEBOOST_cell_64804 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q), .b(FE_OFN1663_n_4490), .c(n_3792), .o(TIMEBOOST_net_16273) );
in01f01 g61876_u0 ( .a(FE_OFN709_n_8232), .o(g61876_sb) );
na02s01 TIMEBOOST_cell_28875 ( .a(n_655), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_), .o(TIMEBOOST_net_8542) );
na03m02 TIMEBOOST_cell_72608 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q), .b(FE_OFN614_n_4501), .c(n_4645), .o(TIMEBOOST_net_306) );
na03m02 TIMEBOOST_cell_72789 ( .a(TIMEBOOST_net_21563), .b(g65037_sb), .c(TIMEBOOST_net_21846), .o(TIMEBOOST_net_17093) );
in01s01 g61877_u0 ( .a(n_8272), .o(g61877_sb) );
na03m06 TIMEBOOST_cell_64533 ( .a(n_3761), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q), .c(FE_OFN670_n_4505), .o(TIMEBOOST_net_14195) );
in01m01 g61878_u0 ( .a(FE_OFN1812_n_7845), .o(g61878_sb) );
na02s01 TIMEBOOST_cell_43459 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q), .o(TIMEBOOST_net_12624) );
na02m02 TIMEBOOST_cell_68271 ( .a(TIMEBOOST_net_21343), .b(g65711_sb), .o(n_2199) );
in01s01 g61879_u0 ( .a(n_8069), .o(g61879_sb) );
na02m02 TIMEBOOST_cell_70085 ( .a(TIMEBOOST_net_22250), .b(FE_OFN701_n_7845), .o(TIMEBOOST_net_20447) );
na02s01 g61879_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q), .b(n_8069), .o(g61879_db) );
na03f02 TIMEBOOST_cell_73509 ( .a(n_6554), .b(TIMEBOOST_net_13380), .c(g62763_sb), .o(n_6117) );
in01m02 g61880_u0 ( .a(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61880_sb) );
na02m10 TIMEBOOST_cell_53005 ( .a(wishbone_slave_unit_pcim_sm_data_in_664), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q), .o(TIMEBOOST_net_16720) );
na02f02 TIMEBOOST_cell_72113 ( .a(TIMEBOOST_net_23264), .b(g64107_sb), .o(TIMEBOOST_net_15073) );
na02s01 g58360_u2 ( .a(FE_OFN270_n_9836), .b(FE_OFN1666_n_9477), .o(g58360_db) );
in01f02 g61881_u0 ( .a(FE_OFN706_n_8119), .o(g61881_sb) );
na02s01 TIMEBOOST_cell_28877 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_), .b(n_599), .o(TIMEBOOST_net_8543) );
na03m02 TIMEBOOST_cell_64831 ( .a(n_3792), .b(TIMEBOOST_net_12347), .c(n_12), .o(TIMEBOOST_net_17109) );
in01f01 g61882_u0 ( .a(FE_OFN707_n_8119), .o(g61882_sb) );
na02f02 TIMEBOOST_cell_72252 ( .a(TIMEBOOST_net_5668), .b(n_8757), .o(TIMEBOOST_net_23334) );
in01f01 g61883_u0 ( .a(FE_OFN710_n_8232), .o(g61883_sb) );
na02f01 TIMEBOOST_cell_71040 ( .a(TIMEBOOST_net_17372), .b(FE_OFN1224_n_6391), .o(TIMEBOOST_net_22728) );
na02m02 TIMEBOOST_cell_54273 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q), .b(TIMEBOOST_net_13010), .o(TIMEBOOST_net_17354) );
na02m02 TIMEBOOST_cell_54383 ( .a(n_3523), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q), .o(TIMEBOOST_net_17409) );
in01s02 g61884_u0 ( .a(FE_OFN2256_n_8060), .o(g61884_sb) );
na02f06 TIMEBOOST_cell_18025 ( .a(n_1826), .b(wishbone_slave_unit_pcim_if_del_we_in), .o(TIMEBOOST_net_5376) );
in01s01 TIMEBOOST_cell_73888 ( .a(n_8295), .o(TIMEBOOST_net_23453) );
na03f02 TIMEBOOST_cell_72953 ( .a(pci_target_unit_del_sync_addr_in_233), .b(g65241_sb), .c(TIMEBOOST_net_7139), .o(n_2641) );
in01m02 g61885_u0 ( .a(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61885_sb) );
na02s01 TIMEBOOST_cell_63004 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q), .o(TIMEBOOST_net_20449) );
na02f02 TIMEBOOST_cell_70013 ( .a(TIMEBOOST_net_22214), .b(g61739_sb), .o(n_8339) );
na02s02 TIMEBOOST_cell_48246 ( .a(TIMEBOOST_net_14340), .b(g57893_db), .o(TIMEBOOST_net_9504) );
in01f01 g61886_u0 ( .a(FE_OFN710_n_8232), .o(g61886_sb) );
na02m02 TIMEBOOST_cell_52707 ( .a(TIMEBOOST_net_12320), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q), .o(TIMEBOOST_net_16571) );
na02f02 TIMEBOOST_cell_71004 ( .a(TIMEBOOST_net_17400), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_22710) );
in01s01 g61887_u0 ( .a(n_8407), .o(g61887_sb) );
na02s01 g61887_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q), .b(n_8407), .o(g61887_db) );
na02s01 TIMEBOOST_cell_38304 ( .a(wbs_adr_i_5_), .b(FE_OFN9_n_11877), .o(TIMEBOOST_net_10764) );
in01f01 g61888_u0 ( .a(FE_OFN712_n_8140), .o(g61888_sb) );
na02s01 TIMEBOOST_cell_62860 ( .a(FE_OFN235_n_9834), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q), .o(TIMEBOOST_net_20377) );
na03s01 TIMEBOOST_cell_68496 ( .a(FE_OFN2095_n_2520), .b(pci_target_unit_del_sync_addr_in_215), .c(parchk_pci_ad_reg_in_1216), .o(TIMEBOOST_net_21456) );
in01s01 g61889_u0 ( .a(n_8176), .o(g61889_sb) );
na02s01 g61889_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q), .b(n_8176), .o(g61889_db) );
na03f02 TIMEBOOST_cell_72983 ( .a(wishbone_slave_unit_pcim_sm_last_in), .b(n_4936), .c(g59384_sb), .o(TIMEBOOST_net_5475) );
in01s02 g61890_u0 ( .a(FE_OFN699_n_7845), .o(g61890_sb) );
in01s01 g61891_u0 ( .a(n_8119), .o(g61891_sb) );
na02s02 TIMEBOOST_cell_52519 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q), .o(TIMEBOOST_net_16477) );
na02s01 g61891_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q), .b(n_8119), .o(g61891_db) );
na02s01 TIMEBOOST_cell_38306 ( .a(wbs_adr_i_4_), .b(FE_OFN9_n_11877), .o(TIMEBOOST_net_10765) );
in01f01 g61892_u0 ( .a(FE_OFN710_n_8232), .o(g61892_sb) );
in01s01 g61893_u0 ( .a(n_8272), .o(g61893_sb) );
na02m04 TIMEBOOST_cell_72115 ( .a(TIMEBOOST_net_23265), .b(g64099_sb), .o(n_4056) );
in01s01 g61894_u0 ( .a(n_8407), .o(g61894_sb) );
na03m02 TIMEBOOST_cell_65131 ( .a(TIMEBOOST_net_20302), .b(g64874_sb), .c(g64874_db), .o(TIMEBOOST_net_13233) );
na02s01 g61894_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q), .b(n_8407), .o(g61894_db) );
na02f02 TIMEBOOST_cell_71480 ( .a(n_3317), .b(FE_OFN1699_n_5751), .o(TIMEBOOST_net_22948) );
in01s01 g61895_u0 ( .a(n_8119), .o(g61895_sb) );
na03f02 TIMEBOOST_cell_73035 ( .a(TIMEBOOST_net_21718), .b(TIMEBOOST_net_16270), .c(FE_OFN1231_n_6391), .o(TIMEBOOST_net_22843) );
na02s01 g61895_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q), .b(n_8119), .o(g61895_db) );
na04f02 TIMEBOOST_cell_73615 ( .a(TIMEBOOST_net_22894), .b(n_8747), .c(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q), .d(g58634_sb), .o(n_8846) );
na02m01 g61896_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q), .b(n_8119), .o(g61896_db) );
na02s01 TIMEBOOST_cell_52521 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q), .o(TIMEBOOST_net_16478) );
in01s01 g61897_u0 ( .a(n_8176), .o(g61897_sb) );
na03f02 TIMEBOOST_cell_72520 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(g64139_sb), .c(g64139_db), .o(n_4024) );
na02s01 g61897_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q), .b(n_8176), .o(g61897_db) );
na03f02 TIMEBOOST_cell_73616 ( .a(TIMEBOOST_net_23375), .b(n_8747), .c(g58632_sb), .o(n_8849) );
na02s01 g61898_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q), .b(n_8407), .o(g61898_db) );
no02s01 TIMEBOOST_cell_52523 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249), .b(FE_RN_240_0), .o(TIMEBOOST_net_16479) );
in01m01 g61899_u0 ( .a(n_8407), .o(g61899_sb) );
in01s01 TIMEBOOST_cell_63552 ( .a(wbs_adr_i_2_), .o(TIMEBOOST_net_20732) );
na02s01 g61899_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q), .b(n_8407), .o(g61899_db) );
na03f02 TIMEBOOST_cell_42408 ( .a(n_3738), .b(g62611_sb), .c(g62611_db), .o(n_6334) );
in01s01 g61900_u0 ( .a(FE_OFN702_n_7845), .o(g61900_sb) );
na03m02 TIMEBOOST_cell_68700 ( .a(FE_OFN1625_n_4438), .b(g64847_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q), .o(TIMEBOOST_net_21558) );
na02m02 TIMEBOOST_cell_50670 ( .a(TIMEBOOST_net_15552), .b(TIMEBOOST_net_11524), .o(TIMEBOOST_net_9537) );
in01m01 g61901_u0 ( .a(FE_OFN2256_n_8060), .o(g61901_sb) );
na02s01 TIMEBOOST_cell_38316 ( .a(g58389_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q), .o(TIMEBOOST_net_10770) );
na02s01 TIMEBOOST_cell_62986 ( .a(conf_wb_err_addr_in_957), .b(configuration_wb_err_addr_548), .o(TIMEBOOST_net_20440) );
in01m01 g61902_u0 ( .a(FE_OFN1812_n_7845), .o(g61902_sb) );
na04m02 TIMEBOOST_cell_67316 ( .a(n_4447), .b(g64885_sb), .c(TIMEBOOST_net_17230), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q), .o(TIMEBOOST_net_17103) );
na03f02 TIMEBOOST_cell_66178 ( .a(TIMEBOOST_net_15232), .b(FE_OFN1179_n_3476), .c(g60614_sb), .o(n_4840) );
in01s01 g61903_u0 ( .a(n_8272), .o(g61903_sb) );
na02m01 TIMEBOOST_cell_54081 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_142), .o(TIMEBOOST_net_17258) );
na02m02 TIMEBOOST_cell_72077 ( .a(TIMEBOOST_net_23246), .b(g64252_db), .o(n_3921) );
in01s01 g61904_u0 ( .a(n_8232), .o(g61904_sb) );
na02f02 TIMEBOOST_cell_70540 ( .a(TIMEBOOST_net_13038), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_22478) );
na02m01 g61904_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q), .b(n_8232), .o(g61904_db) );
in01s01 TIMEBOOST_cell_63565 ( .a(TIMEBOOST_net_20745), .o(TIMEBOOST_net_20744) );
in01f01 g61905_u0 ( .a(FE_OFN706_n_8119), .o(g61905_sb) );
na04m06 TIMEBOOST_cell_72721 ( .a(g65093_sb), .b(g65093_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q), .d(n_4450), .o(TIMEBOOST_net_8852) );
na03f02 TIMEBOOST_cell_66455 ( .a(TIMEBOOST_net_21036), .b(FE_OFN1316_n_6624), .c(g62395_sb), .o(n_7390) );
in01f01 g61906_u0 ( .a(FE_OFN707_n_8119), .o(g61906_sb) );
na03m02 TIMEBOOST_cell_64532 ( .a(n_3792), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q), .c(FE_OFN634_n_4454), .o(TIMEBOOST_net_10393) );
na02s01 TIMEBOOST_cell_62561 ( .a(TIMEBOOST_net_20227), .b(FE_OFN952_n_2055), .o(TIMEBOOST_net_16203) );
in01f02 g61907_u0 ( .a(FE_OFN2212_n_8407), .o(g61907_sb) );
na03f02 TIMEBOOST_cell_66355 ( .a(TIMEBOOST_net_21011), .b(FE_OFN1236_n_6391), .c(g62938_sb), .o(n_6005) );
in01f01 g61908_u0 ( .a(FE_OFN709_n_8232), .o(g61908_sb) );
na02f02 TIMEBOOST_cell_49130 ( .a(TIMEBOOST_net_14782), .b(g61814_sb), .o(n_8163) );
na03f02 TIMEBOOST_cell_73805 ( .a(TIMEBOOST_net_16545), .b(FE_OFN1775_n_13800), .c(FE_OFN1768_n_14054), .o(n_14505) );
in01s01 g61909_u0 ( .a(n_8272), .o(g61909_sb) );
na02f01 TIMEBOOST_cell_71032 ( .a(TIMEBOOST_net_13233), .b(FE_OFN1274_n_4096), .o(TIMEBOOST_net_22724) );
na03f02 TIMEBOOST_cell_66900 ( .a(FE_OFN1748_n_12004), .b(n_12010), .c(TIMEBOOST_net_13548), .o(n_12505) );
in01f01 g61910_u0 ( .a(FE_OFN2081_n_8176), .o(g61910_sb) );
na02s01 TIMEBOOST_cell_39132 ( .a(g58177_sb), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_11178) );
na02f04 TIMEBOOST_cell_47679 ( .a(n_2705), .b(n_1480), .o(TIMEBOOST_net_14057) );
in01f01 g61911_u0 ( .a(FE_OFN701_n_7845), .o(g61911_sb) );
na03m10 TIMEBOOST_cell_72387 ( .a(n_504), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_408), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q), .o(TIMEBOOST_net_20485) );
na03f02 TIMEBOOST_cell_67922 ( .a(TIMEBOOST_net_9971), .b(FE_OFN1100_g64577_p), .c(g62799_sb), .o(n_5386) );
in01m01 g61912_u0 ( .a(FE_OFN2257_n_8060), .o(g61912_sb) );
na03f02 TIMEBOOST_cell_73673 ( .a(TIMEBOOST_net_8334), .b(FE_OFN2105_g64577_p), .c(g63105_sb), .o(n_5044) );
in01f01 g61913_u0 ( .a(FE_OFN709_n_8232), .o(g61913_sb) );
na02f02 TIMEBOOST_cell_70759 ( .a(TIMEBOOST_net_22587), .b(g63202_sb), .o(TIMEBOOST_net_20562) );
na02s01 TIMEBOOST_cell_62560 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q), .o(TIMEBOOST_net_20227) );
na02f02 TIMEBOOST_cell_71553 ( .a(TIMEBOOST_net_22984), .b(FE_OFN1748_n_12004), .o(n_12692) );
in01f01 g61914_u0 ( .a(FE_OFN709_n_8232), .o(g61914_sb) );
na02s01 TIMEBOOST_cell_28911 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_769), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q), .o(TIMEBOOST_net_8560) );
na02s02 TIMEBOOST_cell_43076 ( .a(TIMEBOOST_net_12432), .b(g58210_db), .o(n_9575) );
na02m01 TIMEBOOST_cell_52251 ( .a(n_3741), .b(FE_OFN642_n_4677), .o(TIMEBOOST_net_16343) );
in01s02 g61915_u0 ( .a(FE_OFN704_n_8069), .o(g61915_sb) );
na03m02 TIMEBOOST_cell_72028 ( .a(n_3749), .b(g64948_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q), .o(TIMEBOOST_net_23222) );
na02s01 TIMEBOOST_cell_43080 ( .a(TIMEBOOST_net_12434), .b(FE_OFN531_n_9823), .o(TIMEBOOST_net_8677) );
na04f02 TIMEBOOST_cell_67878 ( .a(FE_OFN644_n_4677), .b(n_4482), .c(TIMEBOOST_net_10757), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q), .o(TIMEBOOST_net_17373) );
in01s02 g61916_u0 ( .a(FE_OFN704_n_8069), .o(g61916_sb) );
na02f02 TIMEBOOST_cell_50508 ( .a(TIMEBOOST_net_15471), .b(g62494_sb), .o(n_6596) );
na02f01 TIMEBOOST_cell_62453 ( .a(TIMEBOOST_net_20173), .b(FE_OFN906_n_4736), .o(TIMEBOOST_net_14140) );
in01m01 g61917_u0 ( .a(FE_OFN1812_n_7845), .o(g61917_sb) );
na02s01 TIMEBOOST_cell_43461 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_12625) );
na03s02 TIMEBOOST_cell_42236 ( .a(g58193_sb), .b(FE_OFN245_n_9114), .c(g58193_db), .o(n_9057) );
in01s01 g61918_u0 ( .a(n_8407), .o(g61918_sb) );
na03f01 TIMEBOOST_cell_64531 ( .a(n_3739), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q), .c(FE_OFN648_n_4497), .o(TIMEBOOST_net_14561) );
na02s01 g61918_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q), .b(n_8407), .o(g61918_db) );
in01s01 TIMEBOOST_cell_63564 ( .a(TIMEBOOST_net_20744), .o(wbs_adr_i_11_) );
in01f01 g61919_u0 ( .a(FE_OFN714_n_8140), .o(g61919_sb) );
na02f01 g64323_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(FE_OFN1034_n_4732), .o(g64323_db) );
na03m02 TIMEBOOST_cell_70018 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q), .b(FE_OFN2257_n_8060), .c(n_1952), .o(TIMEBOOST_net_22217) );
na03m02 TIMEBOOST_cell_65592 ( .a(TIMEBOOST_net_12830), .b(n_8272), .c(g61781_sb), .o(n_8244) );
na02s01 g61920_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q), .b(n_8407), .o(g61920_db) );
na04s02 TIMEBOOST_cell_73074 ( .a(TIMEBOOST_net_10809), .b(g65943_sb), .c(g61889_sb), .d(g61889_db), .o(n_8052) );
in01f02 g61921_u0 ( .a(FE_OFN716_n_8176), .o(g61921_sb) );
na02m02 TIMEBOOST_cell_69219 ( .a(TIMEBOOST_net_21817), .b(TIMEBOOST_net_14514), .o(TIMEBOOST_net_17094) );
na02m04 TIMEBOOST_cell_50921 ( .a(FE_OFN2072_n_15978), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_399), .o(TIMEBOOST_net_15678) );
na04f02 TIMEBOOST_cell_67944 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q), .b(FE_OFN1115_g64577_p), .c(n_3905), .d(g63055_sb), .o(n_5140) );
na02m01 g61922_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q), .b(n_8232), .o(g61922_db) );
na02s01 TIMEBOOST_cell_48014 ( .a(TIMEBOOST_net_14224), .b(FE_OFN237_n_9118), .o(TIMEBOOST_net_10583) );
in01m04 g61923_u0 ( .a(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61923_sb) );
na02m01 g58355_u2 ( .a(FE_OFN268_n_9880), .b(FE_OFN1666_n_9477), .o(g58355_db) );
na02m02 TIMEBOOST_cell_4152 ( .a(g61923_sb), .b(g61923_db), .o(TIMEBOOST_net_636) );
in01s01 g61924_u0 ( .a(n_8069), .o(g61924_sb) );
na02m02 TIMEBOOST_cell_44939 ( .a(n_4437), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q), .o(TIMEBOOST_net_13364) );
na02s01 g61924_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q), .b(n_8069), .o(g61924_db) );
na03f02 TIMEBOOST_cell_67901 ( .a(TIMEBOOST_net_12683), .b(FE_OFN1057_n_4727), .c(g64332_sb), .o(n_4728) );
in01s01 g61925_u0 ( .a(n_8119), .o(g61925_sb) );
na02m02 TIMEBOOST_cell_68967 ( .a(TIMEBOOST_net_21691), .b(g65079_db), .o(TIMEBOOST_net_17493) );
na02s01 g61925_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q), .b(n_8119), .o(g61925_db) );
na02s04 TIMEBOOST_cell_52651 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q), .o(TIMEBOOST_net_16543) );
in01f01 g61926_u0 ( .a(FE_OFN707_n_8119), .o(g61926_sb) );
na03f02 TIMEBOOST_cell_34928 ( .a(TIMEBOOST_net_9497), .b(FE_OFN1413_n_8567), .c(g57400_sb), .o(n_10368) );
na02m01 TIMEBOOST_cell_43096 ( .a(TIMEBOOST_net_12442), .b(FE_OFN928_n_4730), .o(TIMEBOOST_net_10684) );
na02f01 TIMEBOOST_cell_70322 ( .a(TIMEBOOST_net_17312), .b(FE_OFN1100_g64577_p), .o(TIMEBOOST_net_22369) );
in01m01 g61927_u0 ( .a(FE_OFN2256_n_8060), .o(g61927_sb) );
na02f02 TIMEBOOST_cell_52308 ( .a(TIMEBOOST_net_16371), .b(g61769_sb), .o(n_8271) );
na02s02 TIMEBOOST_cell_49412 ( .a(TIMEBOOST_net_14923), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9534) );
na03s01 TIMEBOOST_cell_67805 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_97), .b(FE_OFN2119_wishbone_slave_unit_pci_initiator_if_data_source), .c(g54167_sb), .o(TIMEBOOST_net_14021) );
na02s01 g61928_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q), .b(n_8407), .o(g61928_db) );
na02m80 TIMEBOOST_cell_72170 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .o(TIMEBOOST_net_23293) );
in01s01 g61929_u0 ( .a(n_8272), .o(g61929_sb) );
na03m04 TIMEBOOST_cell_72802 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q), .c(TIMEBOOST_net_14426), .o(TIMEBOOST_net_13249) );
in01s01 g61930_u0 ( .a(n_8272), .o(g61930_sb) );
na02s01 TIMEBOOST_cell_52653 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q), .o(TIMEBOOST_net_16544) );
na02m02 TIMEBOOST_cell_49464 ( .a(TIMEBOOST_net_14949), .b(g57916_sb), .o(TIMEBOOST_net_11193) );
na02f02 TIMEBOOST_cell_63423 ( .a(TIMEBOOST_net_20658), .b(n_2902), .o(TIMEBOOST_net_448) );
in01s01 g61931_u0 ( .a(n_8140), .o(g61931_sb) );
na02m02 TIMEBOOST_cell_70327 ( .a(TIMEBOOST_net_22371), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_15099) );
na02s01 g61931_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q), .b(n_8140), .o(g61931_db) );
na02m04 TIMEBOOST_cell_71886 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q), .b(n_3744), .o(TIMEBOOST_net_23151) );
in01s01 g61932_u0 ( .a(n_8176), .o(g61932_sb) );
na02s01 g61932_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q), .b(n_8176), .o(g61932_db) );
na02s01 TIMEBOOST_cell_18020 ( .a(TIMEBOOST_net_5373), .b(n_13820), .o(TIMEBOOST_net_407) );
in01s01 g61933_u0 ( .a(n_8232), .o(g61933_sb) );
na02s01 TIMEBOOST_cell_18019 ( .a(n_2284), .b(n_12179), .o(TIMEBOOST_net_5373) );
na02m01 g61933_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q), .b(n_8232), .o(g61933_db) );
in01s01 g61934_u0 ( .a(n_8119), .o(g61934_sb) );
na02s01 g61934_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q), .b(n_8119), .o(g61934_db) );
na03f02 TIMEBOOST_cell_34838 ( .a(TIMEBOOST_net_9354), .b(FE_OFN1422_n_8567), .c(g57374_sb), .o(n_11373) );
na02f02 TIMEBOOST_cell_63034 ( .a(n_3968), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q), .o(TIMEBOOST_net_20464) );
na02s01 g61935_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q), .b(n_8407), .o(g61935_db) );
na02m02 TIMEBOOST_cell_68587 ( .a(TIMEBOOST_net_21501), .b(TIMEBOOST_net_10282), .o(TIMEBOOST_net_20585) );
in01m02 g61936_u0 ( .a(FE_OFN1812_n_7845), .o(g61936_sb) );
na02s01 TIMEBOOST_cell_52617 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q), .o(TIMEBOOST_net_16526) );
na03m02 TIMEBOOST_cell_72818 ( .a(g65271_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q), .c(TIMEBOOST_net_20844), .o(TIMEBOOST_net_17059) );
in01f01 g61937_u0 ( .a(FE_OFN716_n_8176), .o(g61937_sb) );
na02m10 TIMEBOOST_cell_45815 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q), .o(TIMEBOOST_net_13802) );
na02m01 TIMEBOOST_cell_43100 ( .a(TIMEBOOST_net_12444), .b(FE_OFN1016_n_2053), .o(TIMEBOOST_net_10696) );
na03f02 TIMEBOOST_cell_66734 ( .a(TIMEBOOST_net_16824), .b(FE_OFN1306_n_13124), .c(g54361_sb), .o(n_13081) );
na02m01 g61938_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q), .b(n_8119), .o(g61938_db) );
na02f01 TIMEBOOST_cell_71582 ( .a(FE_OFN1572_n_11027), .b(TIMEBOOST_net_13630), .o(TIMEBOOST_net_22999) );
in01s01 g61939_u0 ( .a(n_8272), .o(g61939_sb) );
na03s02 TIMEBOOST_cell_72663 ( .a(TIMEBOOST_net_12436), .b(FE_OFN1016_n_2053), .c(g65823_sb), .o(n_1893) );
na02f02 TIMEBOOST_cell_50719 ( .a(TIMEBOOST_net_640), .b(n_7698), .o(TIMEBOOST_net_15577) );
na02s03 TIMEBOOST_cell_54019 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_17227) );
in01f02 g61940_u0 ( .a(FE_OFN713_n_8140), .o(g61940_sb) );
in01s01 TIMEBOOST_cell_63586 ( .a(TIMEBOOST_net_20766), .o(TIMEBOOST_net_20721) );
na02m02 TIMEBOOST_cell_48091 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_123), .o(TIMEBOOST_net_14263) );
in01f02 g61941_u0 ( .a(FE_OFN2212_n_8407), .o(g61941_sb) );
na03f02 TIMEBOOST_cell_72580 ( .a(TIMEBOOST_net_21429), .b(g65089_sb), .c(TIMEBOOST_net_21661), .o(TIMEBOOST_net_20541) );
na02f10 TIMEBOOST_cell_17963 ( .a(pci_target_unit_wbm_sm_pci_tar_burst_ok), .b(n_731), .o(TIMEBOOST_net_5345) );
na03s02 TIMEBOOST_cell_72601 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q), .b(FE_OFN523_n_9428), .c(g58441_sb), .o(TIMEBOOST_net_14979) );
in01m02 g61942_u0 ( .a(FE_OFN2257_n_8060), .o(g61942_sb) );
na02f01 TIMEBOOST_cell_38978 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q), .b(n_13447), .o(TIMEBOOST_net_11101) );
na02f02 TIMEBOOST_cell_68227 ( .a(TIMEBOOST_net_21321), .b(g63590_sb), .o(n_2564) );
in01m02 g61943_u0 ( .a(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61943_sb) );
na03f06 TIMEBOOST_cell_64349 ( .a(n_1160), .b(n_1170), .c(n_2136), .o(TIMEBOOST_net_71) );
in01f01 g61944_u0 ( .a(FE_OFN709_n_8232), .o(g61944_sb) );
in01s01 TIMEBOOST_cell_67773 ( .a(pci_target_unit_fifos_pcir_data_in_174), .o(TIMEBOOST_net_21200) );
na02s01 TIMEBOOST_cell_43108 ( .a(TIMEBOOST_net_12448), .b(FE_OFN955_n_1699), .o(TIMEBOOST_net_10712) );
in01m02 g61945_u0 ( .a(FE_OFN2257_n_8060), .o(g61945_sb) );
na02f01 TIMEBOOST_cell_38980 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q), .b(FE_OFN2059_n_13447), .o(TIMEBOOST_net_11102) );
in01f02 g61946_u0 ( .a(FE_OFN710_n_8232), .o(g61946_sb) );
na02s01 TIMEBOOST_cell_53301 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q), .b(FE_OFN587_n_9692), .o(TIMEBOOST_net_16868) );
na03f01 TIMEBOOST_cell_68120 ( .a(TIMEBOOST_net_13994), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q), .o(TIMEBOOST_net_21268) );
in01m01 g61947_u0 ( .a(FE_OFN2257_n_8060), .o(g61947_sb) );
na02s02 TIMEBOOST_cell_53302 ( .a(TIMEBOOST_net_16868), .b(TIMEBOOST_net_12791), .o(TIMEBOOST_net_9451) );
na03f01 TIMEBOOST_cell_67886 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(g64151_sb), .c(g64151_db), .o(n_4014) );
na02m02 TIMEBOOST_cell_69950 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q), .b(g64307_sb), .o(TIMEBOOST_net_22183) );
in01m04 g61948_u0 ( .a(FE_OFN709_n_8232), .o(g61948_sb) );
na02f02 TIMEBOOST_cell_38982 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q), .b(n_504), .o(TIMEBOOST_net_11103) );
in01s01 TIMEBOOST_cell_45949 ( .a(TIMEBOOST_net_13939), .o(TIMEBOOST_net_13910) );
in01s01 g61949_u0 ( .a(n_8272), .o(g61949_sb) );
na02s01 TIMEBOOST_cell_70087 ( .a(TIMEBOOST_net_22251), .b(FE_OFN2093_n_2301), .o(TIMEBOOST_net_689) );
in01f04 g61950_u0 ( .a(FE_OFN2081_n_8176), .o(g61950_sb) );
na02f02 TIMEBOOST_cell_49388 ( .a(TIMEBOOST_net_14911), .b(g61888_sb), .o(n_8054) );
na03m02 TIMEBOOST_cell_69210 ( .a(TIMEBOOST_net_17224), .b(FE_OFN928_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q), .o(TIMEBOOST_net_21813) );
na03f02 TIMEBOOST_cell_66316 ( .a(TIMEBOOST_net_13367), .b(n_6554), .c(g62421_sb), .o(n_6754) );
in01f02 g61951_u0 ( .a(FE_OFN710_n_8232), .o(g61951_sb) );
na02m08 TIMEBOOST_cell_45795 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_13792) );
na02s02 TIMEBOOST_cell_38443 ( .a(TIMEBOOST_net_10833), .b(g57983_db), .o(n_9816) );
na04f02 TIMEBOOST_cell_67611 ( .a(TIMEBOOST_net_5509), .b(n_3305), .c(TIMEBOOST_net_20993), .d(n_5745), .o(n_7723) );
in01m04 g61952_u0 ( .a(FE_OFN707_n_8119), .o(g61952_sb) );
na02m02 TIMEBOOST_cell_70329 ( .a(TIMEBOOST_net_22372), .b(g63052_db), .o(n_5146) );
na02s02 TIMEBOOST_cell_39731 ( .a(TIMEBOOST_net_11477), .b(g57898_db), .o(n_9226) );
na04f02 TIMEBOOST_cell_73487 ( .a(TIMEBOOST_net_22579), .b(n_8757), .c(TIMEBOOST_net_15245), .d(g52394_sb), .o(n_14803) );
na02s01 g61953_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q), .b(n_7102), .o(g61953_db) );
na02m02 TIMEBOOST_cell_52709 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_143), .o(TIMEBOOST_net_16572) );
in01f01 g61954_u0 ( .a(FE_OFN707_n_8119), .o(g61954_sb) );
na02s01 TIMEBOOST_cell_53371 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q), .o(TIMEBOOST_net_16903) );
na03f02 TIMEBOOST_cell_66833 ( .a(TIMEBOOST_net_15659), .b(g59230_db), .c(g52393_db), .o(n_14828) );
in01f01 g61955_u0 ( .a(FE_OFN1094_g64577_p), .o(g61955_sb) );
in01s01 g61956_u0 ( .a(FE_OFN1097_g64577_p), .o(g61956_sb) );
na02s01 g61956_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q), .b(FE_OFN1097_g64577_p), .o(g61956_db) );
in01f01 g61957_u0 ( .a(FE_OFN1095_g64577_p), .o(g61957_sb) );
na03f01 TIMEBOOST_cell_64530 ( .a(n_3783), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q), .c(FE_OFN1659_n_4490), .o(TIMEBOOST_net_20322) );
na03m02 TIMEBOOST_cell_69902 ( .a(TIMEBOOST_net_17253), .b(FE_OFN1050_n_16657), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q), .o(TIMEBOOST_net_22159) );
in01f01 g61958_u0 ( .a(FE_OFN1094_g64577_p), .o(g61958_sb) );
na02s01 TIMEBOOST_cell_42986 ( .a(TIMEBOOST_net_12387), .b(FE_OFN953_n_2055), .o(TIMEBOOST_net_10454) );
in01s01 g61959_u0 ( .a(FE_OFN1097_g64577_p), .o(g61959_sb) );
na02s01 g61959_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q), .b(FE_OFN1097_g64577_p), .o(g61959_db) );
na02s01 TIMEBOOST_cell_37045 ( .a(TIMEBOOST_net_10134), .b(n_574), .o(TIMEBOOST_net_6813) );
na02f02 TIMEBOOST_cell_53398 ( .a(TIMEBOOST_net_16916), .b(FE_OFN1797_n_2299), .o(TIMEBOOST_net_14570) );
in01m01 g61961_u0 ( .a(FE_OFN1094_g64577_p), .o(g61961_sb) );
na04s02 TIMEBOOST_cell_46274 ( .a(TIMEBOOST_net_10320), .b(g65782_db), .c(g61808_sb), .d(g61808_db), .o(n_8178) );
in01s01 g61962_u0 ( .a(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61962_sb) );
na02s01 TIMEBOOST_cell_54039 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_17237) );
in01s01 TIMEBOOST_cell_73889 ( .a(TIMEBOOST_net_23453), .o(TIMEBOOST_net_23454) );
na03f02 TIMEBOOST_cell_73312 ( .a(TIMEBOOST_net_9945), .b(FE_OFN1139_g64577_p), .c(g62747_sb), .o(n_5486) );
in01f01 g61963_u0 ( .a(FE_OFN1095_g64577_p), .o(g61963_sb) );
na03f02 TIMEBOOST_cell_46083 ( .a(FE_OFN2059_n_13447), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_395), .o(TIMEBOOST_net_12916) );
na03s02 TIMEBOOST_cell_46892 ( .a(TIMEBOOST_net_12951), .b(g58238_sb), .c(TIMEBOOST_net_13116), .o(TIMEBOOST_net_9530) );
in01s01 TIMEBOOST_cell_45877 ( .a(conf_wb_err_addr_in_943), .o(TIMEBOOST_net_13838) );
na02s01 g61964_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61964_db) );
in01s01 TIMEBOOST_cell_73857 ( .a(TIMEBOOST_net_23421), .o(TIMEBOOST_net_23422) );
in01m01 g61965_u0 ( .a(FE_OFN1095_g64577_p), .o(g61965_sb) );
na04f04 TIMEBOOST_cell_73617 ( .a(FE_OFN1244_n_4092), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q), .c(TIMEBOOST_net_15241), .d(g62922_sb), .o(n_6037) );
na02f01 g61965_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q), .b(FE_OFN1095_g64577_p), .o(g61965_db) );
na02s04 TIMEBOOST_cell_68116 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_79), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_21266) );
na02f04 TIMEBOOST_cell_71441 ( .a(TIMEBOOST_net_22928), .b(FE_RN_567_0), .o(FE_RN_569_0) );
na03f02 TIMEBOOST_cell_66779 ( .a(n_3850), .b(g63121_sb), .c(TIMEBOOST_net_7706), .o(n_5014) );
na02f02 TIMEBOOST_cell_49838 ( .a(TIMEBOOST_net_15136), .b(g63038_sb), .o(n_5172) );
na02s01 TIMEBOOST_cell_38224 ( .a(n_2648), .b(g65236_sb), .o(TIMEBOOST_net_10724) );
in01s01 TIMEBOOST_cell_73945 ( .a(TIMEBOOST_net_23509), .o(TIMEBOOST_net_23510) );
na03f02 TIMEBOOST_cell_66360 ( .a(TIMEBOOST_net_20615), .b(FE_OFN1235_n_6391), .c(g63009_sb), .o(n_5864) );
na03f06 TIMEBOOST_cell_64348 ( .a(n_16520), .b(n_15370), .c(n_1299), .o(n_8660) );
na02m02 TIMEBOOST_cell_4154 ( .a(g61923_sb), .b(g61968_db), .o(TIMEBOOST_net_637) );
na02s01 TIMEBOOST_cell_37043 ( .a(TIMEBOOST_net_10133), .b(n_574), .o(TIMEBOOST_net_6812) );
na02s01 g61969_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q), .b(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61969_db) );
na02m04 TIMEBOOST_cell_69040 ( .a(g65098_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q), .o(TIMEBOOST_net_21728) );
na02s04 TIMEBOOST_cell_43834 ( .a(TIMEBOOST_net_12811), .b(g58437_sb), .o(n_9412) );
na02s02 g58326_u2 ( .a(FE_OFN270_n_9836), .b(FE_OFN1657_n_9502), .o(g58326_db) );
na02m01 TIMEBOOST_cell_54041 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q), .b(n_8272), .o(TIMEBOOST_net_17238) );
na02f02 TIMEBOOST_cell_51196 ( .a(TIMEBOOST_net_15815), .b(g62892_sb), .o(n_6093) );
na02m02 TIMEBOOST_cell_4156 ( .a(g61943_sb), .b(g61972_db), .o(TIMEBOOST_net_638) );
na04f04 TIMEBOOST_cell_33813 ( .a(n_2192), .b(g61700_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q), .d(FE_OFN2081_n_8176), .o(n_8428) );
na02m02 TIMEBOOST_cell_4158 ( .a(g61923_sb), .b(g61973_db), .o(TIMEBOOST_net_639) );
na02s01 g58309_u2 ( .a(FE_OFN260_n_9860), .b(FE_OFN1654_n_9502), .o(g58309_db) );
na02f02 TIMEBOOST_cell_49842 ( .a(TIMEBOOST_net_15138), .b(g63066_sb), .o(n_5118) );
na02m02 TIMEBOOST_cell_4142 ( .a(g61943_sb), .b(g61974_db), .o(TIMEBOOST_net_631) );
na02m02 TIMEBOOST_cell_63003 ( .a(TIMEBOOST_net_20448), .b(g57936_sb), .o(TIMEBOOST_net_14358) );
na02s02 g58291_u2 ( .a(FE_OFN270_n_9836), .b(FE_OFN1690_n_9528), .o(g58291_db) );
na03f02 TIMEBOOST_cell_73383 ( .a(TIMEBOOST_net_16708), .b(FE_OFN1301_n_5763), .c(g62060_sb), .o(n_7750) );
na02s02 g58286_u2 ( .a(FE_OFN268_n_9880), .b(FE_OFN1687_n_9528), .o(g58286_db) );
na02m02 TIMEBOOST_cell_4144 ( .a(g61943_sb), .b(g61976_db), .o(TIMEBOOST_net_632) );
na03m02 TIMEBOOST_cell_69010 ( .a(n_3785), .b(g64889_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q), .o(TIMEBOOST_net_21713) );
na02f02 TIMEBOOST_cell_70015 ( .a(TIMEBOOST_net_22215), .b(g61802_sb), .o(n_8191) );
na03s02 TIMEBOOST_cell_67150 ( .a(TIMEBOOST_net_10235), .b(g65688_sb), .c(TIMEBOOST_net_20325), .o(n_8411) );
na02f01 g58280_u2 ( .a(FE_OFN262_n_9851), .b(FE_OFN1690_n_9528), .o(g58280_db) );
na03f20 TIMEBOOST_cell_31902 ( .a(n_657), .b(n_47), .c(n_15302), .o(n_1514) );
na02s01 TIMEBOOST_cell_54043 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q), .o(TIMEBOOST_net_17239) );
na02m01 TIMEBOOST_cell_62558 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_20226) );
na02f02 TIMEBOOST_cell_71039 ( .a(TIMEBOOST_net_22727), .b(g62928_sb), .o(n_6025) );
na02m02 TIMEBOOST_cell_4146 ( .a(g61885_sb), .b(g61980_db), .o(TIMEBOOST_net_633) );
na02s01 TIMEBOOST_cell_45427 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q), .o(TIMEBOOST_net_13608) );
na02m02 TIMEBOOST_cell_4148 ( .a(g61943_sb), .b(g61981_db), .o(TIMEBOOST_net_634) );
na02s01 TIMEBOOST_cell_45587 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q), .o(TIMEBOOST_net_13688) );
na03f02 TIMEBOOST_cell_66361 ( .a(g62971_sb), .b(FE_OFN1234_n_6391), .c(TIMEBOOST_net_21010), .o(n_5940) );
na02s01 g61983_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(g61983_db) );
na02m02 TIMEBOOST_cell_68273 ( .a(TIMEBOOST_net_21344), .b(g65678_sb), .o(n_2211) );
na02m02 TIMEBOOST_cell_25352 ( .a(TIMEBOOST_net_6780), .b(n_940), .o(TIMEBOOST_net_342) );
na02m02 TIMEBOOST_cell_4150 ( .a(g61923_sb), .b(g61985_db), .o(TIMEBOOST_net_635) );
na02f01 TIMEBOOST_cell_25354 ( .a(TIMEBOOST_net_6781), .b(n_1993), .o(TIMEBOOST_net_228) );
na03f02 TIMEBOOST_cell_66895 ( .a(FE_OFN1747_n_12004), .b(n_12010), .c(TIMEBOOST_net_13567), .o(n_12712) );
na03f02 TIMEBOOST_cell_73817 ( .a(TIMEBOOST_net_16551), .b(FE_OFN1773_n_13800), .c(FE_OFN1768_n_14054), .o(g53155_p) );
na02f02 TIMEBOOST_cell_49850 ( .a(TIMEBOOST_net_15142), .b(g62806_sb), .o(n_5368) );
na03f02 TIMEBOOST_cell_65705 ( .a(TIMEBOOST_net_16367), .b(g64236_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q), .o(TIMEBOOST_net_17316) );
na02m02 TIMEBOOST_cell_4138 ( .a(g61923_sb), .b(g61987_db), .o(TIMEBOOST_net_629) );
na02s01 TIMEBOOST_cell_52711 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q), .b(pci_target_unit_fifos_pcir_control_in_192), .o(TIMEBOOST_net_16573) );
na02f40 TIMEBOOST_cell_62394 ( .a(wbm_adr_o_3_), .b(wbm_adr_o_4_), .o(TIMEBOOST_net_20144) );
na02m02 TIMEBOOST_cell_69566 ( .a(FE_OFN953_n_2055), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q), .o(TIMEBOOST_net_21991) );
na03f01 TIMEBOOST_cell_67975 ( .a(TIMEBOOST_net_15230), .b(FE_OFN1179_n_3476), .c(g60618_sb), .o(n_4836) );
na03m02 TIMEBOOST_cell_65726 ( .a(TIMEBOOST_net_306), .b(g64873_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q), .o(TIMEBOOST_net_20973) );
no02s01 TIMEBOOST_cell_25362 ( .a(TIMEBOOST_net_6785), .b(n_692), .o(g65573_p) );
in01s01 g61990_u0 ( .a(n_8069), .o(g61990_sb) );
na04f04 TIMEBOOST_cell_24797 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q), .b(g58805_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q), .d(FE_OFN2158_n_16439), .o(n_8636) );
na02s01 g61990_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q), .b(n_8069), .o(g61990_db) );
na04f02 TIMEBOOST_cell_72705 ( .a(n_3764), .b(g64939_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q), .d(g64939_db), .o(TIMEBOOST_net_17024) );
in01f02 g61991_u0 ( .a(FE_OFN2212_n_8407), .o(g61991_sb) );
na02m01 TIMEBOOST_cell_62470 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q), .b(pci_target_unit_fifos_pciw_control_in_155), .o(TIMEBOOST_net_20182) );
na02m01 TIMEBOOST_cell_48103 ( .a(FE_OFN576_n_9902), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q), .o(TIMEBOOST_net_14269) );
in01s01 g61992_u0 ( .a(n_8069), .o(g61992_sb) );
na02m02 TIMEBOOST_cell_69253 ( .a(TIMEBOOST_net_21834), .b(g65799_sb), .o(n_1590) );
na02s01 g61992_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q), .b(n_8069), .o(g61992_db) );
na02s02 TIMEBOOST_cell_38439 ( .a(TIMEBOOST_net_10831), .b(g57920_db), .o(n_9891) );
in01f01 g61993_u0 ( .a(FE_OFN699_n_7845), .o(g61993_sb) );
na03f04 TIMEBOOST_cell_66972 ( .a(FE_OCP_RBN1973_n_12381), .b(TIMEBOOST_net_16043), .c(n_11831), .o(n_12723) );
na02s02 TIMEBOOST_cell_38405 ( .a(TIMEBOOST_net_10814), .b(g58087_db), .o(n_9709) );
na02f02 TIMEBOOST_cell_70410 ( .a(n_4062), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q), .o(TIMEBOOST_net_22413) );
in01s01 g61994_u0 ( .a(n_8272), .o(g61994_sb) );
na02s01 TIMEBOOST_cell_43468 ( .a(TIMEBOOST_net_12628), .b(FE_OFN1044_n_2037), .o(TIMEBOOST_net_10809) );
na02m01 TIMEBOOST_cell_62454 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_147), .o(TIMEBOOST_net_20174) );
na03f02 TIMEBOOST_cell_584 ( .a(n_3848), .b(g63124_sb), .c(g63124_db), .o(n_5006) );
in01s01 g61995_u0 ( .a(FE_OFN702_n_7845), .o(g61995_sb) );
na04m02 TIMEBOOST_cell_72767 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q), .b(FE_OFN630_n_4454), .c(n_4498), .d(g65027_sb), .o(TIMEBOOST_net_7630) );
na03f02 TIMEBOOST_cell_72655 ( .a(pci_target_unit_fifos_pciw_addr_data_in_127), .b(FE_OFN928_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q), .o(TIMEBOOST_net_22102) );
na02m04 TIMEBOOST_cell_72306 ( .a(FE_OFN272_n_9828), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q), .o(TIMEBOOST_net_23361) );
na02s01 g61996_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q), .b(n_8232), .o(g61996_db) );
na02s01 TIMEBOOST_cell_51537 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q), .o(TIMEBOOST_net_15986) );
in01s01 g61997_u0 ( .a(n_8119), .o(g61997_sb) );
na02f02 TIMEBOOST_cell_71041 ( .a(TIMEBOOST_net_22728), .b(g62423_sb), .o(n_6749) );
na02m01 g61997_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q), .b(n_8119), .o(g61997_db) );
in01m01 g61998_u0 ( .a(FE_OFN699_n_7845), .o(g61998_sb) );
na02m02 TIMEBOOST_cell_70393 ( .a(TIMEBOOST_net_22404), .b(g61815_sb), .o(n_8161) );
na02f02 TIMEBOOST_cell_63164 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q), .b(n_4911), .o(TIMEBOOST_net_20529) );
in01s01 g61999_u0 ( .a(n_8232), .o(g61999_sb) );
na04m04 TIMEBOOST_cell_67903 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(FE_OFN1057_n_4727), .c(g64251_sb), .d(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q), .o(n_3922) );
na02m01 g61999_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q), .b(n_8232), .o(g61999_db) );
na02s01 TIMEBOOST_cell_38425 ( .a(TIMEBOOST_net_10824), .b(g57965_db), .o(TIMEBOOST_net_9455) );
na02m02 TIMEBOOST_cell_68103 ( .a(TIMEBOOST_net_21259), .b(g54219_sb), .o(TIMEBOOST_net_14030) );
in01s01 g62000_u0 ( .a(FE_OFN2258_n_8060), .o(g62000_sb) );
na02m01 g62000_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q), .b(FE_OFN2258_n_8060), .o(g62000_db) );
na04m08 TIMEBOOST_cell_65277 ( .a(g65042_sb), .b(FE_OFN649_n_4497), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q), .d(n_4473), .o(n_4327) );
in01f01 g62001_u0 ( .a(FE_OFN717_n_8176), .o(g62001_sb) );
na02s02 TIMEBOOST_cell_48578 ( .a(TIMEBOOST_net_14506), .b(FE_OFN1689_n_9528), .o(TIMEBOOST_net_10804) );
na02m02 TIMEBOOST_cell_52452 ( .a(TIMEBOOST_net_16443), .b(g58295_db), .o(n_9510) );
in01m01 g62002_u0 ( .a(FE_OFN702_n_7845), .o(g62002_sb) );
na03f02 TIMEBOOST_cell_51259 ( .a(n_1935), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q), .c(FE_OFN2084_n_8407), .o(TIMEBOOST_net_15847) );
na02s01 TIMEBOOST_cell_62859 ( .a(TIMEBOOST_net_20376), .b(g58159_sb), .o(TIMEBOOST_net_14650) );
in01s01 g62003_u0 ( .a(n_8232), .o(g62003_sb) );
na02f02 TIMEBOOST_cell_37971 ( .a(TIMEBOOST_net_10597), .b(g58388_db), .o(n_9443) );
na02m01 g62003_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q), .b(n_8232), .o(g62003_db) );
na02s01 g62004_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q), .b(n_8176), .o(g62004_db) );
na04f02 TIMEBOOST_cell_67905 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q), .b(g65967_sb), .c(g65967_db), .d(TIMEBOOST_net_20882), .o(n_7873) );
in01f02 g62005_u0 ( .a(FE_OFN712_n_8140), .o(g62005_sb) );
na02s01 TIMEBOOST_cell_42808 ( .a(TIMEBOOST_net_12298), .b(FE_OFN935_n_2292), .o(TIMEBOOST_net_10237) );
na02s01 TIMEBOOST_cell_62858 ( .a(FE_OFN235_n_9834), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q), .o(TIMEBOOST_net_20376) );
in01f01 g62006_u0 ( .a(FE_OFN706_n_8119), .o(g62006_sb) );
na03f02 TIMEBOOST_cell_72766 ( .a(n_4488), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q), .c(TIMEBOOST_net_10801), .o(TIMEBOOST_net_20970) );
no04f04 TIMEBOOST_cell_73685 ( .a(TIMEBOOST_net_8576), .b(FE_RN_127_0), .c(TIMEBOOST_net_736), .d(n_7824), .o(g53077_p) );
na03f02 TIMEBOOST_cell_72800 ( .a(n_4498), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q), .c(TIMEBOOST_net_16255), .o(TIMEBOOST_net_17149) );
in01s01 g62007_u0 ( .a(n_8069), .o(g62007_sb) );
na02f02 TIMEBOOST_cell_44694 ( .a(TIMEBOOST_net_13241), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_11588) );
na02s01 g62007_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q), .b(n_8069), .o(g62007_db) );
na03f06 TIMEBOOST_cell_73136 ( .a(TIMEBOOST_net_17278), .b(FE_OFN1075_n_4740), .c(g64117_sb), .o(n_4043) );
na02m02 TIMEBOOST_cell_63332 ( .a(n_4472), .b(n_28), .o(TIMEBOOST_net_20613) );
na02m01 g62008_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q), .b(n_8407), .o(g62008_db) );
in01f01 g62009_u0 ( .a(FE_OFN713_n_8140), .o(g62009_sb) );
na02s01 TIMEBOOST_cell_38580 ( .a(g58144_sb), .b(FE_OFN215_n_9856), .o(TIMEBOOST_net_10902) );
in01m02 g62010_u0 ( .a(FE_OFN706_n_8119), .o(g62010_sb) );
na02s01 TIMEBOOST_cell_38582 ( .a(FE_OFN213_n_9124), .b(g58143_sb), .o(TIMEBOOST_net_10903) );
na03m02 TIMEBOOST_cell_73122 ( .a(g65376_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q), .c(TIMEBOOST_net_14703), .o(TIMEBOOST_net_13077) );
na02m04 TIMEBOOST_cell_53335 ( .a(TIMEBOOST_net_12370), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q), .o(TIMEBOOST_net_16885) );
in01s02 g62011_u0 ( .a(FE_OFN704_n_8069), .o(g62011_sb) );
na02f01 TIMEBOOST_cell_52744 ( .a(TIMEBOOST_net_16589), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_14530) );
na02f01 TIMEBOOST_cell_63037 ( .a(TIMEBOOST_net_20465), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_15124) );
na02f02 TIMEBOOST_cell_70958 ( .a(TIMEBOOST_net_17408), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_22687) );
in01f01 g62012_u0 ( .a(FE_OFN712_n_8140), .o(g62012_sb) );
na03f02 TIMEBOOST_cell_73750 ( .a(n_12099), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q), .o(TIMEBOOST_net_23035) );
na02m01 g62012_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q), .b(n_8140), .o(g62012_db) );
na02s01 TIMEBOOST_cell_62557 ( .a(TIMEBOOST_net_20225), .b(g58164_sb), .o(TIMEBOOST_net_16689) );
in01f02 g62013_u0 ( .a(FE_OFN712_n_8140), .o(g62013_sb) );
na03f02 TIMEBOOST_cell_73230 ( .a(TIMEBOOST_net_14883), .b(g63544_sb), .c(g63544_db), .o(TIMEBOOST_net_8808) );
na02f04 TIMEBOOST_cell_70205 ( .a(TIMEBOOST_net_22310), .b(g54150_sb), .o(n_13450) );
in01s01 TIMEBOOST_cell_73939 ( .a(TIMEBOOST_net_23503), .o(TIMEBOOST_net_23504) );
in01f01 g62014_u0 ( .a(FE_OFN2084_n_8407), .o(g62014_sb) );
na02s01 TIMEBOOST_cell_18008 ( .a(TIMEBOOST_net_5367), .b(n_4686), .o(TIMEBOOST_net_125) );
na02m06 TIMEBOOST_cell_42869 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q), .o(TIMEBOOST_net_12329) );
in01f01 g62015_u0 ( .a(FE_OFN709_n_8232), .o(g62015_sb) );
na02s01 TIMEBOOST_cell_62556 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q), .b(FE_OFN515_n_9697), .o(TIMEBOOST_net_20225) );
na03f02 TIMEBOOST_cell_34747 ( .a(TIMEBOOST_net_9401), .b(FE_OFN1387_n_8567), .c(g57190_sb), .o(n_11562) );
na03f02 TIMEBOOST_cell_34749 ( .a(TIMEBOOST_net_9402), .b(FE_OFN1381_n_8567), .c(g57389_sb), .o(n_10376) );
in01f02 g62016_u0 ( .a(FE_OFN712_n_8140), .o(g62016_sb) );
na02s02 TIMEBOOST_cell_38584 ( .a(FE_OFN241_n_9830), .b(g58092_sb), .o(TIMEBOOST_net_10904) );
na02m04 TIMEBOOST_cell_68556 ( .a(FE_OFN622_n_4409), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q), .o(TIMEBOOST_net_21486) );
na03f02 TIMEBOOST_cell_34751 ( .a(TIMEBOOST_net_9403), .b(FE_OFN1412_n_8567), .c(g57574_sb), .o(n_11177) );
in01f02 g62017_u0 ( .a(FE_OFN2212_n_8407), .o(g62017_sb) );
na02s01 TIMEBOOST_cell_52712 ( .a(TIMEBOOST_net_16573), .b(FE_OFN2111_n_2248), .o(TIMEBOOST_net_14328) );
na03m02 TIMEBOOST_cell_65522 ( .a(g58294_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q), .c(TIMEBOOST_net_11082), .o(TIMEBOOST_net_9359) );
in01f01 g62018_u0 ( .a(FE_OFN2084_n_8407), .o(g62018_sb) );
na02m02 g52460_u1 ( .a(g52460_sb), .b(wbs_adr_i_15_), .o(g52460_da) );
na02f01 TIMEBOOST_cell_26077 ( .a(pci_target_unit_pcit_if_strd_addr_in_710), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_7143) );
in01f02 g62019_u0 ( .a(FE_OFN2212_n_8407), .o(g62019_sb) );
na02m01 TIMEBOOST_cell_38586 ( .a(g58089_sb), .b(FE_OFN235_n_9834), .o(TIMEBOOST_net_10905) );
na03f02 TIMEBOOST_cell_35052 ( .a(TIMEBOOST_net_9604), .b(FE_OFN1441_n_9372), .c(g58473_sb), .o(n_9371) );
na02s01 TIMEBOOST_cell_48537 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q), .b(g65812_sb), .o(TIMEBOOST_net_14486) );
in01m02 g62020_u0 ( .a(FE_OFN1812_n_7845), .o(g62020_sb) );
na02s01 TIMEBOOST_cell_43463 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q), .o(TIMEBOOST_net_12626) );
na02s01 TIMEBOOST_cell_25364 ( .a(TIMEBOOST_net_6786), .b(g57780_sb), .o(TIMEBOOST_net_420) );
na02m02 TIMEBOOST_cell_4140 ( .a(g61923_sb), .b(g62021_db), .o(TIMEBOOST_net_630) );
in01m01 g62022_u0 ( .a(FE_OFN699_n_7845), .o(g62022_sb) );
na03m02 TIMEBOOST_cell_72883 ( .a(n_8272), .b(g61752_sb), .c(TIMEBOOST_net_14739), .o(n_8311) );
na02s02 TIMEBOOST_cell_49791 ( .a(FE_OFN243_n_9116), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q), .o(TIMEBOOST_net_15113) );
in01m01 g62023_u0 ( .a(FE_OFN719_n_8060), .o(g62023_sb) );
na02s01 TIMEBOOST_cell_38588 ( .a(FE_OFN207_n_9865), .b(g58138_sb), .o(TIMEBOOST_net_10906) );
na02f02 TIMEBOOST_cell_17994 ( .a(TIMEBOOST_net_5360), .b(g67040_sb), .o(n_1681) );
in01m01 g62024_u0 ( .a(FE_OFN720_n_8060), .o(g62024_sb) );
na02f02 TIMEBOOST_cell_49770 ( .a(TIMEBOOST_net_15102), .b(g61714_sb), .o(n_8397) );
in01s01 TIMEBOOST_cell_45977 ( .a(pci_target_unit_fifos_pcir_data_in_169), .o(TIMEBOOST_net_13938) );
in01m01 g62025_u0 ( .a(FE_OFN701_n_7845), .o(g62025_sb) );
na02m02 TIMEBOOST_cell_69907 ( .a(TIMEBOOST_net_22161), .b(TIMEBOOST_net_14714), .o(TIMEBOOST_net_17117) );
na02s02 TIMEBOOST_cell_38415 ( .a(TIMEBOOST_net_10819), .b(g57952_db), .o(n_9857) );
na02s02 TIMEBOOST_cell_49793 ( .a(FE_OFN243_n_9116), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q), .o(TIMEBOOST_net_15114) );
in01m01 g62026_u0 ( .a(FE_OFN720_n_8060), .o(g62026_sb) );
na02s01 TIMEBOOST_cell_45443 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q), .o(TIMEBOOST_net_13616) );
in01s01 TIMEBOOST_cell_45947 ( .a(pci_target_unit_fifos_pcir_data_in_159), .o(TIMEBOOST_net_13908) );
na03f02 TIMEBOOST_cell_73384 ( .a(TIMEBOOST_net_16701), .b(FE_OFN1301_n_5763), .c(g62048_sb), .o(n_7762) );
in01m01 g62027_u0 ( .a(FE_OFN699_n_7845), .o(g62027_sb) );
na02m02 TIMEBOOST_cell_62802 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_135), .o(TIMEBOOST_net_20348) );
na02m01 TIMEBOOST_cell_49794 ( .a(TIMEBOOST_net_15114), .b(FE_OFN1803_n_9690), .o(TIMEBOOST_net_12872) );
na03f02 TIMEBOOST_cell_73338 ( .a(TIMEBOOST_net_22420), .b(FE_OFN877_g64577_p), .c(g62814_sb), .o(n_5349) );
in01f01 g62028_u0 ( .a(FE_OFN702_n_7845), .o(g62028_sb) );
na02s02 TIMEBOOST_cell_38590 ( .a(g58074_sb), .b(FE_OFN213_n_9124), .o(TIMEBOOST_net_10907) );
in01m01 g62029_u0 ( .a(FE_OFN702_n_7845), .o(g62029_sb) );
na03f01 TIMEBOOST_cell_64528 ( .a(n_3755), .b(FE_OFN615_n_4501), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q), .o(TIMEBOOST_net_14421) );
in01m01 g62030_u0 ( .a(FE_OFN1700_n_5751), .o(g62030_sb) );
na02m02 g62030_u1 ( .a(wbm_adr_o_23_), .b(g62030_sb), .o(g62030_da) );
na02f02 g62030_u2 ( .a(n_3135), .b(FE_OFN1699_n_5751), .o(g62030_db) );
na04f04 TIMEBOOST_cell_67693 ( .a(TIMEBOOST_net_16857), .b(FE_OFN2200_n_10256), .c(g52596_sb), .d(TIMEBOOST_net_703), .o(n_11875) );
in01f02 g62031_u0 ( .a(FE_OFN1145_n_15261), .o(g62031_sb) );
na02m01 TIMEBOOST_cell_62626 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q), .b(n_8272), .o(TIMEBOOST_net_20260) );
in01f01 g62032_u0 ( .a(FE_OFN1300_n_5763), .o(g62032_sb) );
na03f02 TIMEBOOST_cell_73717 ( .a(n_12010), .b(TIMEBOOST_net_13551), .c(FE_OFN1746_n_12004), .o(n_12633) );
na03m02 TIMEBOOST_cell_72649 ( .a(TIMEBOOST_net_21491), .b(g65071_sb), .c(TIMEBOOST_net_21681), .o(TIMEBOOST_net_17441) );
na02m01 TIMEBOOST_cell_25370 ( .a(TIMEBOOST_net_6789), .b(n_2299), .o(TIMEBOOST_net_109) );
in01f02 g62033_u0 ( .a(FE_OFN1143_n_15261), .o(g62033_sb) );
na02s02 TIMEBOOST_cell_49413 ( .a(FE_OFN270_n_9836), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q), .o(TIMEBOOST_net_14924) );
na02f02 TIMEBOOST_cell_3637 ( .a(TIMEBOOST_net_378), .b(n_8538), .o(n_8659) );
in01f01 g62034_u0 ( .a(FE_OFN1302_n_5763), .o(g62034_sb) );
na02m08 g52465_u1 ( .a(g52461_sb), .b(wbs_adr_i_19_), .o(g52465_da) );
in01s01 TIMEBOOST_cell_63567 ( .a(TIMEBOOST_net_20747), .o(TIMEBOOST_net_20746) );
in01f02 g62035_u0 ( .a(FE_OFN1301_n_5763), .o(g62035_sb) );
na03m02 TIMEBOOST_cell_72890 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q), .b(g64306_sb), .c(TIMEBOOST_net_12792), .o(n_3869) );
na02m01 TIMEBOOST_cell_25376 ( .a(TIMEBOOST_net_6792), .b(n_2299), .o(TIMEBOOST_net_107) );
in01f02 g62036_u0 ( .a(FE_OFN1301_n_5763), .o(g62036_sb) );
na03s02 TIMEBOOST_cell_72889 ( .a(g65819_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q), .c(TIMEBOOST_net_10696), .o(TIMEBOOST_net_14591) );
na02s01 TIMEBOOST_cell_25380 ( .a(TIMEBOOST_net_6794), .b(n_1349), .o(n_1963) );
na03f04 TIMEBOOST_cell_46033 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q), .b(n_7822), .c(pci_target_unit_pcit_if_pcir_fifo_data_in_772), .o(TIMEBOOST_net_12849) );
in01f02 g62037_u0 ( .a(FE_OFN1301_n_5763), .o(g62037_sb) );
na03f02 TIMEBOOST_cell_66817 ( .a(TIMEBOOST_net_17102), .b(FE_OFN1310_n_6624), .c(g62407_sb), .o(n_6785) );
na02m01 TIMEBOOST_cell_48599 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q), .b(n_3783), .o(TIMEBOOST_net_14517) );
in01f01 g62038_u0 ( .a(FE_OFN1302_n_5763), .o(g62038_sb) );
na04f04 TIMEBOOST_cell_73385 ( .a(configuration_pci_err_data_527), .b(FE_OFN1186_n_3476), .c(wbm_dat_o_26_), .d(g60658_sb), .o(n_5663) );
in01f01 g62039_u0 ( .a(FE_OFN1302_n_5763), .o(g62039_sb) );
na02m02 TIMEBOOST_cell_54336 ( .a(TIMEBOOST_net_17385), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_15349) );
in01s01 TIMEBOOST_cell_73844 ( .a(n_727), .o(TIMEBOOST_net_23409) );
na02m10 TIMEBOOST_cell_45313 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q), .o(TIMEBOOST_net_13551) );
in01f01 g62040_u0 ( .a(FE_OFN1302_n_5763), .o(g62040_sb) );
na02s02 TIMEBOOST_cell_69884 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(g64200_sb), .o(TIMEBOOST_net_22150) );
in01f02 g62041_u0 ( .a(FE_OFN1301_n_5763), .o(g62041_sb) );
na02m01 TIMEBOOST_cell_54083 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_139), .o(TIMEBOOST_net_17259) );
in01s03 TIMEBOOST_cell_63566 ( .a(TIMEBOOST_net_20746), .o(wbs_adr_i_28_) );
in01f01 g62042_u0 ( .a(FE_OFN1302_n_5763), .o(g62042_sb) );
na03f02 TIMEBOOST_cell_66457 ( .a(TIMEBOOST_net_17110), .b(FE_OFN1317_n_6624), .c(g62484_sb), .o(n_6620) );
na03f04 TIMEBOOST_cell_66870 ( .a(n_12228), .b(FE_OFN1749_n_12004), .c(TIMEBOOST_net_21083), .o(n_12623) );
in01f02 g62043_u0 ( .a(FE_OFN1299_n_5763), .o(g62043_sb) );
na02s01 TIMEBOOST_cell_45395 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q), .o(TIMEBOOST_net_13592) );
in01f01 g62044_u0 ( .a(FE_OFN1300_n_5763), .o(g62044_sb) );
na02f01 TIMEBOOST_cell_54084 ( .a(TIMEBOOST_net_17259), .b(FE_OFN1032_n_4732), .o(TIMEBOOST_net_14754) );
na02s01 TIMEBOOST_cell_25412 ( .a(TIMEBOOST_net_6810), .b(FE_OFN946_n_2248), .o(TIMEBOOST_net_152) );
na02s01 TIMEBOOST_cell_25414 ( .a(TIMEBOOST_net_6811), .b(FE_OFN946_n_2248), .o(TIMEBOOST_net_147) );
in01f01 g62045_u0 ( .a(FE_OFN1302_n_5763), .o(g62045_sb) );
na02s02 TIMEBOOST_cell_48833 ( .a(FE_OFN231_n_9839), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q), .o(TIMEBOOST_net_14634) );
na02f01 TIMEBOOST_cell_25416 ( .a(TIMEBOOST_net_6812), .b(g67051_sb), .o(n_1503) );
na02f01 TIMEBOOST_cell_25418 ( .a(TIMEBOOST_net_6813), .b(g67051_sb), .o(n_1444) );
in01f02 g62046_u0 ( .a(FE_OFN1299_n_5763), .o(g62046_sb) );
na04f80 TIMEBOOST_cell_35542 ( .a(pci_trdy_i), .b(g67082_sb), .c(output_backup_trdy_out_reg_Q), .d(parchk_pci_trdy_en_in), .o(n_1192) );
na02s02 TIMEBOOST_cell_52816 ( .a(TIMEBOOST_net_16625), .b(g64226_sb), .o(n_4516) );
na02m20 TIMEBOOST_cell_48689 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_123), .o(TIMEBOOST_net_14562) );
in01f01 g62047_u0 ( .a(FE_OFN1302_n_5763), .o(g62047_sb) );
na03m02 TIMEBOOST_cell_67353 ( .a(n_1858), .b(g61859_db), .c(g61859_sb), .o(n_8121) );
in01f02 g62048_u0 ( .a(FE_OFN1301_n_5763), .o(g62048_sb) );
na02s01 TIMEBOOST_cell_25426 ( .a(TIMEBOOST_net_6817), .b(g56934_sb), .o(TIMEBOOST_net_691) );
na02m02 TIMEBOOST_cell_52919 ( .a(TIMEBOOST_net_13043), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_16677) );
in01f02 g62049_u0 ( .a(FE_OFN1301_n_5763), .o(g62049_sb) );
na02s01 TIMEBOOST_cell_25428 ( .a(TIMEBOOST_net_6818), .b(g57797_sb), .o(TIMEBOOST_net_713) );
na02s01 TIMEBOOST_cell_64198 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q), .o(TIMEBOOST_net_21085) );
in01f02 g62050_u0 ( .a(FE_OFN1301_n_5763), .o(g62050_sb) );
na02s01 TIMEBOOST_cell_25430 ( .a(TIMEBOOST_net_6819), .b(g56934_sb), .o(TIMEBOOST_net_769) );
na02f06 TIMEBOOST_cell_25432 ( .a(TIMEBOOST_net_6820), .b(n_2256), .o(TIMEBOOST_net_121) );
in01f02 g62051_u0 ( .a(FE_OFN1299_n_5763), .o(g62051_sb) );
in01s01 TIMEBOOST_cell_72353 ( .a(TIMEBOOST_net_23386), .o(TIMEBOOST_net_23385) );
in01f02 g62052_u0 ( .a(FE_OFN1301_n_5763), .o(g62052_sb) );
na02m20 TIMEBOOST_cell_52353 ( .a(pci_target_unit_pcit_if_strd_addr_in_702), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66), .o(TIMEBOOST_net_16394) );
na03s01 TIMEBOOST_cell_64416 ( .a(TIMEBOOST_net_20794), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_391), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q), .o(TIMEBOOST_net_16802) );
in01f01 g62053_u0 ( .a(FE_OFN1302_n_5763), .o(g62053_sb) );
na02s01 TIMEBOOST_cell_31841 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__Q), .b(wbu_sel_in_314), .o(TIMEBOOST_net_10025) );
na02f04 TIMEBOOST_cell_45230 ( .a(TIMEBOOST_net_13509), .b(FE_RN_456_0), .o(FE_RN_457_0) );
na02m10 TIMEBOOST_cell_45231 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q), .o(TIMEBOOST_net_13510) );
in01f02 g62054_u0 ( .a(FE_OFN1302_n_5763), .o(g62054_sb) );
na02m06 TIMEBOOST_cell_72120 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q), .o(TIMEBOOST_net_23268) );
in01f02 g62055_u0 ( .a(FE_OFN1299_n_5763), .o(g62055_sb) );
na02m02 TIMEBOOST_cell_69024 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q), .b(FE_OFN639_n_4669), .o(TIMEBOOST_net_21720) );
na03f04 TIMEBOOST_cell_70164 ( .a(FE_OFN1074_n_4740), .b(pci_target_unit_fifos_pciw_addr_data_in_145), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q), .o(TIMEBOOST_net_22290) );
na03m02 TIMEBOOST_cell_73137 ( .a(TIMEBOOST_net_23257), .b(FE_OFN1077_n_4740), .c(g64084_sb), .o(TIMEBOOST_net_15028) );
in01f02 g62056_u0 ( .a(FE_OFN1301_n_5763), .o(g62056_sb) );
na02m02 TIMEBOOST_cell_50040 ( .a(TIMEBOOST_net_15237), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_13297) );
na03m02 TIMEBOOST_cell_72631 ( .a(g65026_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q), .c(TIMEBOOST_net_10401), .o(TIMEBOOST_net_17464) );
in01f02 g62057_u0 ( .a(FE_OFN1302_n_5763), .o(g62057_sb) );
na02m02 TIMEBOOST_cell_53855 ( .a(TIMEBOOST_net_7597), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q), .o(TIMEBOOST_net_17145) );
na02s03 TIMEBOOST_cell_72020 ( .a(TIMEBOOST_net_12451), .b(FE_OFN955_n_1699), .o(TIMEBOOST_net_23218) );
in01s01 TIMEBOOST_cell_73978 ( .a(wbm_dat_i_9_), .o(TIMEBOOST_net_23543) );
in01f01 g62058_u0 ( .a(FE_OFN2079_n_8069), .o(g62058_sb) );
na02s02 TIMEBOOST_cell_42777 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q), .b(n_8831), .o(TIMEBOOST_net_12283) );
na02f02 TIMEBOOST_cell_49882 ( .a(TIMEBOOST_net_15158), .b(g63110_sb), .o(n_5036) );
na03f02 TIMEBOOST_cell_73386 ( .a(TIMEBOOST_net_16442), .b(FE_OFN1184_n_3476), .c(g60608_sb), .o(n_4846) );
in01f02 g62059_u0 ( .a(FE_OFN1299_n_5763), .o(g62059_sb) );
na02m04 TIMEBOOST_cell_68648 ( .a(g64808_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q), .o(TIMEBOOST_net_21532) );
na04f04 TIMEBOOST_cell_42527 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_787), .c(FE_OFN2135_n_13124), .d(g54352_sb), .o(n_13089) );
na02m02 TIMEBOOST_cell_53207 ( .a(n_1423), .b(TIMEBOOST_net_686), .o(TIMEBOOST_net_16821) );
in01f02 g62060_u0 ( .a(FE_OFN1301_n_5763), .o(g62060_sb) );
in01s01 TIMEBOOST_cell_67775 ( .a(pci_target_unit_fifos_pcir_data_in_188), .o(TIMEBOOST_net_21202) );
in01s01 TIMEBOOST_cell_73946 ( .a(wbm_dat_i_23_), .o(TIMEBOOST_net_23511) );
na03f02 TIMEBOOST_cell_66222 ( .a(TIMEBOOST_net_20527), .b(FE_OFN1264_n_4095), .c(g62903_sb), .o(n_6071) );
in01f01 g62061_u0 ( .a(FE_OFN1300_n_5763), .o(g62061_sb) );
na02m02 TIMEBOOST_cell_71478 ( .a(TIMEBOOST_net_16444), .b(g52404_sb), .o(TIMEBOOST_net_22947) );
na02f02 TIMEBOOST_cell_70551 ( .a(TIMEBOOST_net_22483), .b(g63031_sb), .o(n_5185) );
in01f01 g62062_u0 ( .a(FE_OFN1300_n_5763), .o(g62062_sb) );
na03f02 TIMEBOOST_cell_66818 ( .a(TIMEBOOST_net_17171), .b(FE_OFN1345_n_8567), .c(g57115_sb), .o(n_11631) );
na03m02 TIMEBOOST_cell_64526 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q), .b(n_3783), .c(FE_OFN612_n_4501), .o(TIMEBOOST_net_16240) );
in01f02 g62063_u0 ( .a(FE_OFN1301_n_5763), .o(g62063_sb) );
na02f02 TIMEBOOST_cell_53858 ( .a(TIMEBOOST_net_17146), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_15387) );
na03f01 TIMEBOOST_cell_64525 ( .a(n_3752), .b(n_3616), .c(FE_OFN618_n_4490), .o(TIMEBOOST_net_14389) );
na02m01 TIMEBOOST_cell_72008 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q), .b(FE_OFN644_n_4677), .o(TIMEBOOST_net_23212) );
in01f02 g62064_u0 ( .a(FE_OFN1302_n_5763), .o(g62064_sb) );
na04f06 TIMEBOOST_cell_20897 ( .a(n_1343), .b(n_1344), .c(n_1253), .d(n_1341), .o(n_2401) );
na02s01 TIMEBOOST_cell_44047 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q), .o(TIMEBOOST_net_12918) );
in01f02 g62065_u0 ( .a(FE_OFN1301_n_5763), .o(g62065_sb) );
na03f02 TIMEBOOST_cell_34917 ( .a(TIMEBOOST_net_9513), .b(FE_OFN1382_n_8567), .c(g57437_sb), .o(n_11297) );
na03m02 TIMEBOOST_cell_71898 ( .a(n_3752), .b(g64833_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q), .o(TIMEBOOST_net_23157) );
na03m04 TIMEBOOST_cell_72707 ( .a(g64811_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q), .c(TIMEBOOST_net_16266), .o(TIMEBOOST_net_17565) );
in01s01 g62066_u0 ( .a(FE_OFN2079_n_8069), .o(g62066_sb) );
na03f02 TIMEBOOST_cell_72112 ( .a(FE_OFN1049_n_16657), .b(TIMEBOOST_net_16617), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q), .o(TIMEBOOST_net_23264) );
na02s01 TIMEBOOST_cell_44015 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(FE_OFN1041_n_2037), .o(TIMEBOOST_net_12902) );
in01f02 g62067_u0 ( .a(FE_OFN1700_n_5751), .o(g62067_sb) );
in01s01 TIMEBOOST_cell_45926 ( .a(TIMEBOOST_net_13886), .o(TIMEBOOST_net_13887) );
na02f06 TIMEBOOST_cell_3455 ( .a(TIMEBOOST_net_287), .b(n_3378), .o(n_8750) );
in01f02 g62068_u0 ( .a(FE_OFN1699_n_5751), .o(g62068_sb) );
in01s01 TIMEBOOST_cell_45878 ( .a(TIMEBOOST_net_13838), .o(TIMEBOOST_net_13839) );
na02f04 g62068_u2 ( .a(n_2720), .b(FE_OFN1699_n_5751), .o(g62068_db) );
na02s06 TIMEBOOST_cell_43083 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q), .o(TIMEBOOST_net_12436) );
in01s01 g62069_u0 ( .a(FE_OFN2079_n_8069), .o(g62069_sb) );
na02s01 TIMEBOOST_cell_43131 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q), .o(TIMEBOOST_net_12460) );
na04m02 TIMEBOOST_cell_72722 ( .a(g65063_sb), .b(g65063_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q), .d(n_4452), .o(TIMEBOOST_net_17545) );
na02m02 TIMEBOOST_cell_51953 ( .a(FE_OFN917_n_4725), .b(TIMEBOOST_net_12378), .o(TIMEBOOST_net_16194) );
in01s01 g62070_u0 ( .a(FE_OFN2079_n_8069), .o(g62070_sb) );
na03f02 TIMEBOOST_cell_66459 ( .a(TIMEBOOST_net_16773), .b(FE_OFN1311_n_6624), .c(g62425_sb), .o(n_6747) );
na02f02 TIMEBOOST_cell_70638 ( .a(TIMEBOOST_net_20914), .b(FE_OCPN1909_n_16497), .o(TIMEBOOST_net_22527) );
in01f02 g62071_u0 ( .a(FE_OFN2079_n_8069), .o(g62071_sb) );
na02m08 TIMEBOOST_cell_43033 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_148), .o(TIMEBOOST_net_12411) );
na03f02 TIMEBOOST_cell_67970 ( .a(TIMEBOOST_net_13222), .b(n_2843), .c(n_3236), .o(n_4808) );
in01s01 TIMEBOOST_cell_67750 ( .a(TIMEBOOST_net_21176), .o(TIMEBOOST_net_21177) );
in01f02 g62072_u0 ( .a(n_5633), .o(g62072_sb) );
na02m01 TIMEBOOST_cell_53057 ( .a(configuration_pci_err_addr_499), .b(wbm_adr_o_29_), .o(TIMEBOOST_net_16746) );
na04f04 TIMEBOOST_cell_67695 ( .a(TIMEBOOST_net_16866), .b(FE_OFN2200_n_10256), .c(g52607_sb), .d(TIMEBOOST_net_697), .o(n_11864) );
in01f04 g62073_u0 ( .a(FE_OFN1174_n_5592), .o(g62073_sb) );
na02m01 TIMEBOOST_cell_37638 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q), .b(FE_OFN666_n_4495), .o(TIMEBOOST_net_10431) );
in01s01 TIMEBOOST_cell_64264 ( .a(pci_target_unit_fifos_pcir_data_in_170), .o(TIMEBOOST_net_21120) );
na02m08 TIMEBOOST_cell_52525 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q), .o(TIMEBOOST_net_16480) );
in01f02 g62074_u0 ( .a(FE_OFN1170_n_5592), .o(g62074_sb) );
na03f02 TIMEBOOST_cell_66966 ( .a(FE_OCPN1866_n_12377), .b(TIMEBOOST_net_8609), .c(FE_OFN1756_n_12681), .o(n_12668) );
na03f02 TIMEBOOST_cell_73231 ( .a(TIMEBOOST_net_12928), .b(g64165_sb), .c(TIMEBOOST_net_17308), .o(TIMEBOOST_net_22582) );
in01f02 g62075_u0 ( .a(FE_OFN1163_n_5615), .o(g62075_sb) );
na03f02 TIMEBOOST_cell_72583 ( .a(TIMEBOOST_net_21436), .b(g64750_sb), .c(TIMEBOOST_net_22103), .o(TIMEBOOST_net_17411) );
na02m02 TIMEBOOST_cell_68160 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q), .b(FE_OFN2055_n_8831), .o(TIMEBOOST_net_21288) );
in01f02 g62076_u0 ( .a(FE_OFN1174_n_5592), .o(g62076_sb) );
na04f04 TIMEBOOST_cell_67442 ( .a(n_4477), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q), .c(FE_OFN1236_n_6391), .d(g62402_sb), .o(n_6795) );
in01f02 g62077_u0 ( .a(n_5633), .o(g62077_sb) );
na03m02 TIMEBOOST_cell_67391 ( .a(wbs_adr_i_28_), .b(g52462_sb), .c(FE_OFN1021_n_11877), .o(TIMEBOOST_net_706) );
na04f06 TIMEBOOST_cell_73138 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q), .b(FE_OFN1074_n_4740), .c(pci_target_unit_fifos_pciw_addr_data_in_123), .d(g64094_sb), .o(n_4061) );
na02s02 TIMEBOOST_cell_48379 ( .a(g58338_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q), .o(TIMEBOOST_net_14407) );
in01f02 g62078_u0 ( .a(n_5633), .o(g62078_sb) );
na03f02 TIMEBOOST_cell_1091 ( .a(n_4077), .b(g63124_sb), .c(g62724_db), .o(n_5534) );
na03f02 TIMEBOOST_cell_73659 ( .a(TIMEBOOST_net_22422), .b(n_3921), .c(g63142_sb), .o(n_4963) );
na03f02 TIMEBOOST_cell_66461 ( .a(TIMEBOOST_net_20612), .b(g54173_sb), .c(TIMEBOOST_net_646), .o(n_13496) );
in01f02 g62079_u0 ( .a(FE_OFN1163_n_5615), .o(g62079_sb) );
na02f01 TIMEBOOST_cell_69438 ( .a(n_4442), .b(n_38), .o(TIMEBOOST_net_21927) );
na03m02 TIMEBOOST_cell_72554 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN685_n_4417), .c(TIMEBOOST_net_21713), .o(TIMEBOOST_net_17558) );
in01f02 g62080_u0 ( .a(FE_OFN1169_n_5592), .o(g62080_sb) );
na03m02 TIMEBOOST_cell_72469 ( .a(FE_OFN576_n_9902), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q), .c(g58075_sb), .o(TIMEBOOST_net_17266) );
na02m08 TIMEBOOST_cell_52527 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q), .o(TIMEBOOST_net_16481) );
na03f02 TIMEBOOST_cell_64347 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q), .b(n_12595), .c(pci_target_unit_pcit_if_pcir_fifo_data_in_795), .o(TIMEBOOST_net_20914) );
in01f02 g62081_u0 ( .a(FE_OFN1169_n_5592), .o(g62081_sb) );
na02f01 TIMEBOOST_cell_42878 ( .a(TIMEBOOST_net_12333), .b(FE_OFN959_n_2299), .o(TIMEBOOST_net_10317) );
na02m02 TIMEBOOST_cell_68848 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q), .o(TIMEBOOST_net_21632) );
na02m02 TIMEBOOST_cell_68891 ( .a(TIMEBOOST_net_21653), .b(n_4493), .o(TIMEBOOST_net_16213) );
in01f02 g62082_u0 ( .a(FE_OFN1173_n_5592), .o(g62082_sb) );
na02m01 TIMEBOOST_cell_38002 ( .a(g58082_sb), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_10613) );
na04m08 TIMEBOOST_cell_67478 ( .a(g58105_db), .b(FE_OFN239_n_9832), .c(g58105_sb), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q), .o(TIMEBOOST_net_16849) );
in01f02 g62083_u0 ( .a(FE_OFN1173_n_5592), .o(g62083_sb) );
na02f02 TIMEBOOST_cell_70845 ( .a(TIMEBOOST_net_22630), .b(g62038_sb), .o(n_7777) );
na02f01 TIMEBOOST_cell_68161 ( .a(TIMEBOOST_net_21288), .b(wbu_addr_in_275), .o(TIMEBOOST_net_12304) );
in01f02 g62084_u0 ( .a(FE_OFN1165_n_5615), .o(g62084_sb) );
na03f02 TIMEBOOST_cell_70626 ( .a(TIMEBOOST_net_20417), .b(TIMEBOOST_net_7219), .c(FE_OFN877_g64577_p), .o(TIMEBOOST_net_22521) );
na02s01 TIMEBOOST_cell_52529 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q), .o(TIMEBOOST_net_16482) );
na02m01 TIMEBOOST_cell_69605 ( .a(TIMEBOOST_net_22010), .b(FE_OFN1031_n_4732), .o(TIMEBOOST_net_20413) );
in01f02 g62085_u0 ( .a(FE_OFN1173_n_5592), .o(g62085_sb) );
na02s01 TIMEBOOST_cell_42992 ( .a(TIMEBOOST_net_12390), .b(FE_OFN950_n_2055), .o(TIMEBOOST_net_10461) );
na04m02 TIMEBOOST_cell_67313 ( .a(g64801_sb), .b(n_4479), .c(g64801_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q), .o(TIMEBOOST_net_20610) );
in01f02 g62086_u0 ( .a(FE_OFN1173_n_5592), .o(g62086_sb) );
na02m02 TIMEBOOST_cell_54613 ( .a(n_3760), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q), .o(TIMEBOOST_net_17524) );
na03f02 TIMEBOOST_cell_66304 ( .a(TIMEBOOST_net_20986), .b(g52440_sb), .c(TIMEBOOST_net_15556), .o(n_14812) );
in01f02 g62087_u0 ( .a(FE_OFN1173_n_5592), .o(g62087_sb) );
na04f02 TIMEBOOST_cell_73618 ( .a(TIMEBOOST_net_21060), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .c(n_8747), .d(g58622_sb), .o(n_8854) );
na02m04 TIMEBOOST_cell_68484 ( .a(g64772_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q), .o(TIMEBOOST_net_21450) );
in01f02 g62088_u0 ( .a(FE_OFN1173_n_5592), .o(g62088_sb) );
na02s01 TIMEBOOST_cell_38592 ( .a(g58066_sb), .b(FE_OFN252_n_9868), .o(TIMEBOOST_net_10908) );
na03f02 TIMEBOOST_cell_73619 ( .a(TIMEBOOST_net_23376), .b(n_8747), .c(g58630_sb), .o(n_8851) );
in01f02 g62089_u0 ( .a(FE_OFN1164_n_5615), .o(g62089_sb) );
na02m10 TIMEBOOST_cell_28997 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q), .o(TIMEBOOST_net_8603) );
in01f02 g62090_u0 ( .a(n_5633), .o(g62090_sb) );
na02m02 TIMEBOOST_cell_48316 ( .a(TIMEBOOST_net_14375), .b(g58316_sb), .o(TIMEBOOST_net_11211) );
na03f02 TIMEBOOST_cell_73461 ( .a(TIMEBOOST_net_8852), .b(FE_OFN1215_n_4151), .c(g62559_sb), .o(n_6443) );
na03m02 TIMEBOOST_cell_73123 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q), .b(g64261_sb), .c(g64261_db), .o(n_3912) );
in01f02 g62091_u0 ( .a(FE_OFN1164_n_5615), .o(g62091_sb) );
na02s02 TIMEBOOST_cell_28185 ( .a(TIMEBOOST_net_21193), .b(g65733_sb), .o(TIMEBOOST_net_8197) );
na04f02 TIMEBOOST_cell_73620 ( .a(TIMEBOOST_net_16821), .b(n_11), .c(n_8747), .d(g58598_sb), .o(n_8855) );
na02m02 TIMEBOOST_cell_63978 ( .a(n_263), .b(n_4902), .o(TIMEBOOST_net_20975) );
in01f02 g62092_u0 ( .a(FE_OFN1173_n_5592), .o(g62092_sb) );
no02f02 TIMEBOOST_cell_28943 ( .a(FE_RN_361_0), .b(FE_OFN1706_n_4868), .o(TIMEBOOST_net_8576) );
na04f06 TIMEBOOST_cell_64296 ( .a(n_1698), .b(n_1061), .c(n_2648), .d(FE_RN_305_0), .o(TIMEBOOST_net_216) );
na03f02 TIMEBOOST_cell_47278 ( .a(FE_OFN1733_n_16317), .b(TIMEBOOST_net_13576), .c(FE_OFN1738_n_11019), .o(n_12651) );
in01f02 g62093_u0 ( .a(FE_OFN1168_n_5592), .o(g62093_sb) );
na03f02 TIMEBOOST_cell_64295 ( .a(n_2411), .b(n_1227), .c(n_2929), .o(TIMEBOOST_net_317) );
na03f02 TIMEBOOST_cell_47280 ( .a(FE_OFN1736_n_16317), .b(TIMEBOOST_net_13578), .c(FE_OFN1742_n_11019), .o(n_12517) );
in01f02 g62094_u0 ( .a(n_5633), .o(g62094_sb) );
na03f02 TIMEBOOST_cell_66628 ( .a(TIMEBOOST_net_8540), .b(FE_OCPN1847_n_14981), .c(g59110_sb), .o(n_8693) );
na02f02 TIMEBOOST_cell_50684 ( .a(TIMEBOOST_net_15559), .b(g62846_sb), .o(n_5279) );
na02m04 TIMEBOOST_cell_45471 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q), .o(TIMEBOOST_net_13630) );
in01f02 g62095_u0 ( .a(n_5633), .o(g62095_sb) );
na03f02 TIMEBOOST_cell_65966 ( .a(TIMEBOOST_net_20447), .b(g65906_da), .c(g61873_sb), .o(n_8087) );
na02m01 TIMEBOOST_cell_42882 ( .a(TIMEBOOST_net_12335), .b(FE_OFN904_n_4736), .o(TIMEBOOST_net_10323) );
in01f02 g62096_u0 ( .a(FE_OFN1168_n_5592), .o(g62096_sb) );
na02f01 TIMEBOOST_cell_37304 ( .a(n_2376), .b(FE_OFN989_n_574), .o(TIMEBOOST_net_10264) );
na02m01 TIMEBOOST_cell_52979 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q), .b(wishbone_slave_unit_pcim_sm_data_in_665), .o(TIMEBOOST_net_16707) );
na03f02 TIMEBOOST_cell_34891 ( .a(TIMEBOOST_net_9416), .b(FE_OFN1397_n_8567), .c(g57247_sb), .o(n_10424) );
in01f02 g62097_u0 ( .a(FE_OFN1168_n_5592), .o(g62097_sb) );
na02s01 TIMEBOOST_cell_52537 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_16486) );
na03f04 TIMEBOOST_cell_64294 ( .a(n_1968), .b(n_2872), .c(n_1969), .o(TIMEBOOST_net_265) );
in01f02 g62098_u0 ( .a(FE_OFN1168_n_5592), .o(g62098_sb) );
na03m04 TIMEBOOST_cell_72632 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q), .c(TIMEBOOST_net_12742), .o(TIMEBOOST_net_17498) );
na02s01 TIMEBOOST_cell_52539 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q), .o(TIMEBOOST_net_16487) );
in01f02 g62099_u0 ( .a(FE_OFN1163_n_5615), .o(g62099_sb) );
na03f02 TIMEBOOST_cell_47282 ( .a(FE_OFN1734_n_16317), .b(TIMEBOOST_net_13580), .c(FE_OFN1739_n_11019), .o(n_12680) );
in01f02 g62100_u0 ( .a(FE_OFN1168_n_5592), .o(g62100_sb) );
na02f04 TIMEBOOST_cell_47715 ( .a(n_1481), .b(n_2914), .o(TIMEBOOST_net_14075) );
na02f01 TIMEBOOST_cell_50005 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_), .b(FE_OFN1117_g64577_p), .o(TIMEBOOST_net_15220) );
na02s01 TIMEBOOST_cell_52541 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q), .o(TIMEBOOST_net_16488) );
in01f02 g62101_u0 ( .a(n_5633), .o(g62101_sb) );
na03m04 TIMEBOOST_cell_73105 ( .a(TIMEBOOST_net_22058), .b(g65350_sb), .c(TIMEBOOST_net_23277), .o(TIMEBOOST_net_20581) );
na03f02 TIMEBOOST_cell_34833 ( .a(TIMEBOOST_net_9445), .b(FE_OFN1413_n_8567), .c(g57466_sb), .o(n_10343) );
in01f02 g62102_u0 ( .a(FE_OFN1164_n_5615), .o(g62102_sb) );
na02s01 TIMEBOOST_cell_52543 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q), .o(TIMEBOOST_net_16489) );
na02s01 TIMEBOOST_cell_52545 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q), .o(TIMEBOOST_net_16490) );
in01f02 g62103_u0 ( .a(FE_OFN1164_n_5615), .o(g62103_sb) );
na03s02 TIMEBOOST_cell_41936 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q), .b(g58277_sb), .c(g58277_db), .o(n_9525) );
na02m02 TIMEBOOST_cell_64098 ( .a(n_323), .b(n_4903), .o(TIMEBOOST_net_21035) );
na03f02 TIMEBOOST_cell_67977 ( .a(TIMEBOOST_net_8840), .b(FE_OFN1183_n_3476), .c(g60615_sb), .o(n_4839) );
in01f02 g62104_u0 ( .a(FE_OFN1163_n_5615), .o(g62104_sb) );
na02s01 TIMEBOOST_cell_68514 ( .a(n_2541), .b(g66398_sb), .o(TIMEBOOST_net_21465) );
na02s02 TIMEBOOST_cell_72100 ( .a(pci_target_unit_fifos_pciw_addr_data_in_128), .b(g64090_sb), .o(TIMEBOOST_net_23258) );
in01f02 g62105_u0 ( .a(FE_OFN1174_n_5592), .o(g62105_sb) );
na03m02 TIMEBOOST_cell_73106 ( .a(TIMEBOOST_net_10708), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q), .c(TIMEBOOST_net_16343), .o(TIMEBOOST_net_17403) );
na02s01 TIMEBOOST_cell_52547 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q), .o(TIMEBOOST_net_16491) );
in01f01 g62106_u0 ( .a(n_5633), .o(g62106_sb) );
na03f02 TIMEBOOST_cell_69120 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(g63543_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q), .o(TIMEBOOST_net_21768) );
na02f02 g62106_u2 ( .a(configuration_wb_err_data_575), .b(n_5633), .o(g62106_db) );
na02m02 TIMEBOOST_cell_25621 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54), .b(pci_target_unit_pcit_if_strd_addr_in_690), .o(TIMEBOOST_net_6915) );
in01f02 g62107_u0 ( .a(FE_OFN1174_n_5592), .o(g62107_sb) );
na02m06 TIMEBOOST_cell_28565 ( .a(configuration_pci_err_addr_473), .b(wbm_adr_o_3_), .o(TIMEBOOST_net_8387) );
na02f02 TIMEBOOST_cell_63951 ( .a(TIMEBOOST_net_20961), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_15474) );
in01f02 g62108_u0 ( .a(FE_OFN1174_n_5592), .o(g62108_sb) );
na03f02 TIMEBOOST_cell_73621 ( .a(TIMEBOOST_net_23377), .b(n_8747), .c(g58631_sb), .o(n_8850) );
na03f02 TIMEBOOST_cell_67980 ( .a(TIMEBOOST_net_20968), .b(FE_OFN1284_n_4097), .c(g62539_sb), .o(n_6490) );
na02s01 TIMEBOOST_cell_52549 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q), .o(TIMEBOOST_net_16492) );
in01f02 g62109_u0 ( .a(FE_OFN1169_n_5592), .o(g62109_sb) );
na03f02 TIMEBOOST_cell_73387 ( .a(TIMEBOOST_net_16736), .b(FE_OFN1185_n_3476), .c(g60610_sb), .o(n_4844) );
na03f02 TIMEBOOST_cell_47286 ( .a(FE_OFN1734_n_16317), .b(TIMEBOOST_net_13583), .c(FE_OFN1739_n_11019), .o(n_12696) );
na02s01 TIMEBOOST_cell_52551 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q), .o(TIMEBOOST_net_16493) );
in01f02 g62110_u0 ( .a(FE_OFN1165_n_5615), .o(g62110_sb) );
na04s02 TIMEBOOST_cell_67844 ( .a(TIMEBOOST_net_12392), .b(g65684_sb), .c(g61743_sb), .d(g61743_db), .o(n_8331) );
na03f02 TIMEBOOST_cell_67979 ( .a(TIMEBOOST_net_8842), .b(FE_OFN1183_n_3476), .c(g60604_sb), .o(n_4851) );
in01f01 g62111_u0 ( .a(n_5633), .o(g62111_sb) );
na02s01 TIMEBOOST_cell_48556 ( .a(TIMEBOOST_net_14495), .b(g65855_sb), .o(n_1873) );
na02f01 g62111_u2 ( .a(configuration_wb_err_addr_542), .b(n_5633), .o(g62111_db) );
na03f02 TIMEBOOST_cell_73818 ( .a(TIMEBOOST_net_16549), .b(FE_OFN1775_n_13800), .c(FE_OFN1768_n_14054), .o(g53242_p) );
in01f04 g62112_u0 ( .a(FE_OFN1171_n_5592), .o(g62112_sb) );
na02m02 TIMEBOOST_cell_71934 ( .a(FE_OFN644_n_4677), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q), .o(TIMEBOOST_net_23175) );
na02s01 TIMEBOOST_cell_52553 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q), .o(TIMEBOOST_net_16494) );
in01f01 g62113_u0 ( .a(FE_OFN1170_n_5592), .o(g62113_sb) );
na04m01 TIMEBOOST_cell_72418 ( .a(FE_OFN276_n_9941), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q), .c(g57795_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_), .o(TIMEBOOST_net_21313) );
na02m06 TIMEBOOST_cell_69034 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q), .b(g65295_sb), .o(TIMEBOOST_net_21725) );
in01f01 g62114_u0 ( .a(n_5633), .o(g62114_sb) );
na02f01 TIMEBOOST_cell_18273 ( .a(n_3449), .b(n_7608), .o(TIMEBOOST_net_5500) );
na02f02 g62114_u2 ( .a(configuration_wb_err_addr_545), .b(n_5633), .o(g62114_db) );
in01f01 g62115_u0 ( .a(FE_OFN1166_n_5615), .o(g62115_sb) );
na02s01 TIMEBOOST_cell_52555 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q), .o(TIMEBOOST_net_16495) );
na02s01 TIMEBOOST_cell_50031 ( .a(wbm_dat_o_25_), .b(configuration_pci_err_data_526), .o(TIMEBOOST_net_15233) );
in01f02 g62116_u0 ( .a(n_5633), .o(g62116_sb) );
na03f02 TIMEBOOST_cell_66378 ( .a(TIMEBOOST_net_17407), .b(FE_OFN1270_n_4095), .c(g62693_sb), .o(n_6162) );
in01s02 TIMEBOOST_cell_67777 ( .a(pci_target_unit_fifos_pcir_data_in_178), .o(TIMEBOOST_net_21204) );
na02s06 TIMEBOOST_cell_47557 ( .a(wbs_dat_i_24_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q), .o(TIMEBOOST_net_13996) );
in01f02 g62117_u0 ( .a(FE_OFN1166_n_5615), .o(g62117_sb) );
na04f04 TIMEBOOST_cell_42478 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q), .b(n_13179), .c(FE_OFN1331_n_13547), .d(g53908_sb), .o(n_13533) );
in01f02 g62118_u0 ( .a(FE_OFN1171_n_5592), .o(g62118_sb) );
na02s01 TIMEBOOST_cell_45087 ( .a(g61868_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_13438) );
na03f02 TIMEBOOST_cell_67982 ( .a(TIMEBOOST_net_20981), .b(FE_OFN1293_n_4098), .c(g62639_sb), .o(n_6271) );
na04f04 TIMEBOOST_cell_42482 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q), .b(n_13228), .c(FE_OFN1332_n_13547), .d(g53910_sb), .o(n_13531) );
in01f01 g62119_u0 ( .a(n_5633), .o(g62119_sb) );
na04f04 TIMEBOOST_cell_42484 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q), .b(n_13180), .c(FE_OFN1331_n_13547), .d(g53907_sb), .o(n_13534) );
na02f01 g62119_u2 ( .a(configuration_wb_err_addr_550), .b(n_5633), .o(g62119_db) );
na02m08 TIMEBOOST_cell_52557 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q), .o(TIMEBOOST_net_16496) );
in01f02 g62120_u0 ( .a(FE_OFN1170_n_5592), .o(g62120_sb) );
na03s01 TIMEBOOST_cell_64714 ( .a(pci_target_unit_del_sync_addr_in_225), .b(g66406_sb), .c(g66418_db), .o(n_2514) );
na02m02 TIMEBOOST_cell_50032 ( .a(TIMEBOOST_net_15233), .b(FE_OFN1186_n_3476), .o(TIMEBOOST_net_13291) );
na03s02 TIMEBOOST_cell_69644 ( .a(TIMEBOOST_net_14272), .b(TIMEBOOST_net_10293), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q), .o(TIMEBOOST_net_22030) );
in01f01 g62121_u0 ( .a(FE_OFN1171_n_5592), .o(g62121_sb) );
na03f02 TIMEBOOST_cell_67981 ( .a(TIMEBOOST_net_17575), .b(FE_OFN1268_n_4095), .c(g62680_sb), .o(n_6179) );
in01f01 g62122_u0 ( .a(FE_OFN1172_n_5592), .o(g62122_sb) );
na02m01 TIMEBOOST_cell_37644 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q), .b(FE_OFN904_n_4736), .o(TIMEBOOST_net_10434) );
na02s01 TIMEBOOST_cell_52559 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q), .o(TIMEBOOST_net_16497) );
na03f02 TIMEBOOST_cell_73388 ( .a(TIMEBOOST_net_16437), .b(FE_OFN1184_n_3476), .c(g60616_sb), .o(n_4838) );
in01f02 g62123_u0 ( .a(FE_OFN1171_n_5592), .o(g62123_sb) );
na02f01 TIMEBOOST_cell_37646 ( .a(FE_OFN902_n_4736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q), .o(TIMEBOOST_net_10435) );
na02s01 TIMEBOOST_cell_52561 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q), .o(TIMEBOOST_net_16498) );
no02s01 TIMEBOOST_cell_52563 ( .a(FE_RN_717_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377), .o(TIMEBOOST_net_16499) );
in01f02 g62124_u0 ( .a(n_5633), .o(g62124_sb) );
na02m02 TIMEBOOST_cell_68930 ( .a(n_4444), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q), .o(TIMEBOOST_net_21673) );
na02m01 TIMEBOOST_cell_42884 ( .a(TIMEBOOST_net_12336), .b(FE_OFN904_n_4736), .o(TIMEBOOST_net_10324) );
na03f02 TIMEBOOST_cell_34913 ( .a(TIMEBOOST_net_9489), .b(FE_OFN1414_n_8567), .c(g57327_sb), .o(n_11423) );
in01f02 g62125_u0 ( .a(FE_OFN1170_n_5592), .o(g62125_sb) );
na03f02 TIMEBOOST_cell_72974 ( .a(TIMEBOOST_net_20348), .b(FE_OFN1055_n_4727), .c(g64233_sb), .o(n_3939) );
na02s02 TIMEBOOST_cell_68248 ( .a(n_8884), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q), .o(TIMEBOOST_net_21332) );
na02s01 TIMEBOOST_cell_50039 ( .a(configuration_pci_err_data_523), .b(wbm_dat_o_22_), .o(TIMEBOOST_net_15237) );
in01f02 g62126_u0 ( .a(FE_OFN1170_n_5592), .o(g62126_sb) );
na02m01 TIMEBOOST_cell_68892 ( .a(n_4479), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q), .o(TIMEBOOST_net_21654) );
in01f02 g62127_u0 ( .a(FE_OFN1172_n_5592), .o(g62127_sb) );
na02s01 TIMEBOOST_cell_69782 ( .a(FE_OFN548_n_9477), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q), .o(TIMEBOOST_net_22099) );
na02s01 TIMEBOOST_cell_52565 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q), .o(TIMEBOOST_net_16500) );
na03m02 TIMEBOOST_cell_68836 ( .a(g64978_sb), .b(n_4645), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q), .o(TIMEBOOST_net_21626) );
in01f02 g62128_u0 ( .a(FE_OFN1171_n_5592), .o(g62128_sb) );
na02s01 TIMEBOOST_cell_52567 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_16501) );
in01f02 g62129_u0 ( .a(FE_OFN1166_n_5615), .o(g62129_sb) );
na02m01 TIMEBOOST_cell_37181 ( .a(TIMEBOOST_net_10202), .b(n_4730), .o(TIMEBOOST_net_178) );
na02m02 TIMEBOOST_cell_49207 ( .a(n_8892), .b(FE_OFN1671_n_9477), .o(TIMEBOOST_net_14821) );
in01f02 g62130_u0 ( .a(FE_OFN1171_n_5592), .o(g62130_sb) );
na02s02 TIMEBOOST_cell_38396 ( .a(g58130_sb), .b(FE_OFN241_n_9830), .o(TIMEBOOST_net_10810) );
na03f02 TIMEBOOST_cell_73389 ( .a(TIMEBOOST_net_16727), .b(FE_OFN1184_n_3476), .c(g60649_sb), .o(n_5676) );
in01f02 g62131_u0 ( .a(FE_OFN1171_n_5592), .o(g62131_sb) );
na02f02 TIMEBOOST_cell_70209 ( .a(TIMEBOOST_net_22312), .b(n_3269), .o(TIMEBOOST_net_7603) );
na02s01 TIMEBOOST_cell_52569 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q), .o(TIMEBOOST_net_16502) );
na03f01 TIMEBOOST_cell_68722 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q), .c(FE_OFN1626_n_4438), .o(TIMEBOOST_net_21569) );
in01f02 g62132_u0 ( .a(n_5633), .o(g62132_sb) );
na03m02 TIMEBOOST_cell_65561 ( .a(TIMEBOOST_net_10705), .b(g65288_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q), .o(TIMEBOOST_net_17412) );
na02f02 TIMEBOOST_cell_44855 ( .a(TIMEBOOST_net_8843), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_13322) );
in01f02 g62133_u0 ( .a(n_5633), .o(g62133_sb) );
na03f02 TIMEBOOST_cell_44291 ( .a(TIMEBOOST_net_10958), .b(g65252_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q), .o(TIMEBOOST_net_13040) );
na02s01 TIMEBOOST_cell_43095 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q), .o(TIMEBOOST_net_12442) );
in01f01 g62134_u0 ( .a(n_5633), .o(g62134_sb) );
na03f02 TIMEBOOST_cell_66575 ( .a(TIMEBOOST_net_13060), .b(FE_OFN1112_g64577_p), .c(g63072_sb), .o(n_5106) );
na02f02 g62134_u2 ( .a(configuration_wb_err_addr_535), .b(n_5633), .o(g62134_db) );
in01f02 g62135_u0 ( .a(FE_OFN1166_n_5615), .o(g62135_sb) );
na03m02 TIMEBOOST_cell_69776 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(FE_OFN927_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q), .o(TIMEBOOST_net_22096) );
na02m01 TIMEBOOST_cell_50043 ( .a(configuration_pci_err_addr_500), .b(wbm_adr_o_30_), .o(TIMEBOOST_net_15239) );
na02s01 TIMEBOOST_cell_52571 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q), .o(TIMEBOOST_net_16503) );
in01f02 g62136_u0 ( .a(FE_OFN1171_n_5592), .o(g62136_sb) );
na02s01 TIMEBOOST_cell_52573 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q), .o(TIMEBOOST_net_16504) );
in01f02 g62137_u0 ( .a(FE_OFN1171_n_5592), .o(g62137_sb) );
na02m10 TIMEBOOST_cell_52805 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_144), .o(TIMEBOOST_net_16620) );
na02s01 TIMEBOOST_cell_52575 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_16505) );
in01f02 g62138_u0 ( .a(FE_OFN1170_n_5592), .o(g62138_sb) );
na02f02 TIMEBOOST_cell_42994 ( .a(TIMEBOOST_net_12391), .b(g58777_sb), .o(n_9849) );
na02s01 TIMEBOOST_cell_38400 ( .a(g58233_sb), .b(FE_OFN213_n_9124), .o(TIMEBOOST_net_10812) );
in01f04 g62139_u0 ( .a(FE_OFN1171_n_5592), .o(g62139_sb) );
na02m01 TIMEBOOST_cell_42886 ( .a(TIMEBOOST_net_12337), .b(FE_OFN904_n_4736), .o(TIMEBOOST_net_10325) );
na03f02 TIMEBOOST_cell_73718 ( .a(n_12001), .b(TIMEBOOST_net_13555), .c(FE_OFN1747_n_12004), .o(n_12704) );
na02s02 TIMEBOOST_cell_38404 ( .a(FE_OFN233_n_9876), .b(g58087_sb), .o(TIMEBOOST_net_10814) );
in01f01 g62140_u0 ( .a(FE_OFN1166_n_5615), .o(g62140_sb) );
in01s01 TIMEBOOST_cell_73979 ( .a(TIMEBOOST_net_23543), .o(TIMEBOOST_net_23544) );
na02s01 TIMEBOOST_cell_52577 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q), .o(TIMEBOOST_net_16506) );
na02s02 TIMEBOOST_cell_38406 ( .a(FE_OFN221_n_9846), .b(g58080_sb), .o(TIMEBOOST_net_10815) );
in01f04 g62141_u0 ( .a(FE_OFN1174_n_5592), .o(g62141_sb) );
na02s01 TIMEBOOST_cell_38408 ( .a(FE_OFN252_n_9868), .b(g58037_sb), .o(TIMEBOOST_net_10816) );
na02m04 TIMEBOOST_cell_50047 ( .a(TIMEBOOST_net_10617), .b(g65308_sb), .o(TIMEBOOST_net_15241) );
in01m02 g62143_u0 ( .a(n_2035), .o(n_2281) );
in01s01 g62144_u0 ( .a(n_1694), .o(n_1695) );
in01f01 g62145_u0 ( .a(n_1692), .o(n_1693) );
na02f10 g62193_u0 ( .a(n_15931), .b(n_1698), .o(n_7427) );
na02f10 g62194_u0 ( .a(n_15931), .b(n_2044), .o(n_7420) );
na02f20 g62195_u0 ( .a(n_15931), .b(n_1061), .o(n_7410) );
na02f02 g62196_u0 ( .a(n_7466), .b(FE_OCPN1854_n_2071), .o(n_7437) );
oa12f02 g62197_u0 ( .a(configuration_wb_err_cs_bit8), .b(n_3282), .c(n_8440), .o(n_7743) );
na02f20 g62198_u0 ( .a(FE_OFN1158_n_15325), .b(n_1061), .o(n_7015) );
na02f04 g62199_u0 ( .a(n_7809), .b(FE_OCPN1854_n_2071), .o(n_7810) );
na02f08 g62200_u0 ( .a(n_7803), .b(FE_OCPN1854_n_2071), .o(n_7804) );
oa12m02 g62201_u0 ( .a(configuration_isr_bit_2975), .b(n_3800), .c(n_8440), .o(n_7742) );
na02f10 g62202_u0 ( .a(n_7466), .b(n_1698), .o(n_7467) );
oa12f02 g62203_u0 ( .a(configuration_status_bit8), .b(n_3257), .c(n_8440), .o(n_7740) );
oa12f01 g62204_u0 ( .a(configuration_status_bit_322), .b(n_3256), .c(n_8440), .o(n_7739) );
na02f20 g62205_u0 ( .a(n_16916), .b(n_1698), .o(n_7283) );
na02f10 g62207_u0 ( .a(n_16916), .b(n_2044), .o(n_7273) );
na02f20 g62208_u0 ( .a(FE_OFN1159_n_15325), .b(n_1698), .o(n_7012) );
na02f20 g62209_u0 ( .a(FE_OFN1159_n_15325), .b(n_2044), .o(n_7007) );
na02f20 g62210_u0 ( .a(n_16916), .b(n_1061), .o(n_7293) );
oa12s01 g62211_u0 ( .a(configuration_status_bit_435), .b(n_3255), .c(n_8440), .o(n_7738) );
oa12m03 g62212_u0 ( .a(configuration_status_bit_379), .b(n_3258), .c(n_8440), .o(n_7737) );
oa12s02 g62213_u0 ( .a(configuration_status_bit_351), .b(n_3262), .c(n_8440), .o(n_7735) );
oa12f01 g62214_u0 ( .a(configuration_status_bit_407), .b(n_3254), .c(n_8440), .o(n_7734) );
na02f10 g62215_u0 ( .a(n_7795), .b(FE_OCPN1854_n_2071), .o(n_7796) );
no02f40 g62217_u0 ( .a(n_4686), .b(n_4685), .o(n_4853) );
in01f02 g62218_u0 ( .a(n_4815), .o(n_4816) );
no02f20 g62219_u0 ( .a(n_2708), .b(n_4685), .o(g62219_p) );
in01f20 g62219_u1 ( .a(g62219_p), .o(n_4815) );
na02f10 g62220_u0 ( .a(n_1390), .b(n_2680), .o(g62220_p) );
in01f08 g62220_u1 ( .a(g62220_p), .o(n_2970) );
na02f10 g62221_u0 ( .a(n_2463), .b(n_2738), .o(g62221_p) );
in01f08 g62221_u1 ( .a(g62221_p), .o(n_2873) );
na02f01 g62222_u0 ( .a(FE_OCP_RBN2222_n_15347), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_6944) );
na02f06 g62223_u0 ( .a(wishbone_slave_unit_wishbone_slave_do_del_request), .b(FE_OCP_RBN2220_n_15347), .o(g62223_p) );
in01f04 g62223_u1 ( .a(g62223_p), .o(n_4814) );
na03f02 g62224_u0 ( .a(n_15435), .b(n_2898), .c(n_15436), .o(n_4188) );
na02m04 g62225_u0 ( .a(FE_OFN1169_n_5592), .b(configuration_wb_err_cs_bit9), .o(n_4813) );
na02m04 TIMEBOOST_cell_52807 ( .a(pci_target_unit_pcit_if_strd_addr_in_699), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63), .o(TIMEBOOST_net_16621) );
na02f10 g62254_u0 ( .a(n_3342), .b(n_3341), .o(g62254_p) );
in01f10 g62254_u1 ( .a(g62254_p), .o(n_3476) );
na02f01 TIMEBOOST_cell_44292 ( .a(TIMEBOOST_net_13040), .b(FE_OFN1128_g64577_p), .o(TIMEBOOST_net_11318) );
oa12f02 g62258_u0 ( .a(n_4123), .b(n_2972), .c(n_2127), .o(n_4812) );
na02f02 g62259_u0 ( .a(FE_OFN2079_n_8069), .b(n_8876), .o(n_7733) );
no02s01 g62260_u0 ( .a(n_2721), .b(FE_OFN778_n_4152), .o(n_3162) );
ao12f01 g62261_u0 ( .a(configuration_sync_pci_err_cs_8_del_bit_reg_Q), .b(n_4721), .c(n_4743), .o(n_7574) );
na02f02 g62262_u0 ( .a(n_3436), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_7078) );
na02f06 g62263_u0 ( .a(FE_OFN2079_n_8069), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .o(n_7731) );
na02f06 g62264_u0 ( .a(n_2461), .b(n_2680), .o(g62264_p) );
in01f06 g62264_u1 ( .a(g62264_p), .o(n_2462) );
na02f04 g62265_u0 ( .a(FE_OFN1171_n_5592), .b(configuration_wb_err_addr), .o(n_4811) );
no02f02 g62267_u0 ( .a(n_7398), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_7725) );
na02f04 g62273_u0 ( .a(n_1111), .b(n_13825), .o(n_6942) );
na02f04 g62274_u0 ( .a(wishbone_slave_unit_pcim_sm_be_in_558), .b(n_13825), .o(n_6941) );
na02f04 g62275_u0 ( .a(wishbone_slave_unit_pcim_sm_be_in_559), .b(n_13825), .o(n_6940) );
in01f04 g62277_u0 ( .a(n_2460), .o(n_2735) );
no02f20 g62278_u0 ( .a(n_1639), .b(n_2011), .o(n_2460) );
no02f02 g62279_u0 ( .a(n_2940), .b(FE_OFN1142_n_15261), .o(n_3339) );
na03f02 TIMEBOOST_cell_66075 ( .a(n_3857), .b(g63112_sb), .c(TIMEBOOST_net_7714), .o(n_5031) );
no02f04 g62281_u0 ( .a(n_2941), .b(FE_OFN1144_n_15261), .o(n_3338) );
no02f02 g62282_u0 ( .a(n_3136), .b(FE_OFN1145_n_15261), .o(n_3468) );
ao12s01 g62283_u0 ( .a(configuration_sync_isr_2_del_bit_reg_Q), .b(n_3799), .c(n_4743), .o(n_7571) );
na03s02 TIMEBOOST_cell_65250 ( .a(TIMEBOOST_net_20270), .b(FE_OFN1793_n_9904), .c(g58053_sb), .o(n_9735) );
na02f08 g62285_u0 ( .a(n_3160), .b(wishbone_slave_unit_pcim_if_del_we_in), .o(g62285_p) );
in01f04 g62285_u1 ( .a(g62285_p), .o(n_3391) );
no02f04 g62286_u0 ( .a(FE_OFN1172_n_5592), .b(n_16763), .o(n_4809) );
na03f01 TIMEBOOST_cell_64521 ( .a(n_3747), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q), .c(FE_OFN1642_n_4671), .o(TIMEBOOST_net_20293) );
no02f02 g62288_u0 ( .a(n_2943), .b(n_692), .o(n_3337) );
no02f02 g62289_u0 ( .a(n_16163), .b(pci_target_unit_wishbone_master_retried), .o(TIMEBOOST_net_10068) );
no02f01 g62290_u0 ( .a(n_2010), .b(FE_OFN778_n_4152), .o(n_2980) );
na02f01 TIMEBOOST_cell_52826 ( .a(TIMEBOOST_net_16630), .b(FE_OFN1076_n_4740), .o(TIMEBOOST_net_14874) );
na02f01 g62293_u0 ( .a(n_7350), .b(n_7569), .o(n_8503) );
na02f10 g62294_u0 ( .a(n_15920), .b(n_15347), .o(n_15014) );
na02m01 TIMEBOOST_cell_50041 ( .a(wbm_adr_o_7_), .b(configuration_pci_err_addr_477), .o(TIMEBOOST_net_15238) );
na02s01 TIMEBOOST_cell_45315 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q), .o(TIMEBOOST_net_13552) );
na04f04 TIMEBOOST_cell_42463 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q), .b(n_13167), .c(FE_OFN1331_n_13547), .d(g53925_sb), .o(n_13520) );
na02m02 TIMEBOOST_cell_71978 ( .a(FE_OFN653_n_4508), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q), .o(TIMEBOOST_net_23197) );
na04m06 TIMEBOOST_cell_67209 ( .a(g64989_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q), .c(FE_OFN684_n_4417), .d(n_4498), .o(n_4359) );
na04m08 TIMEBOOST_cell_67211 ( .a(g64997_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q), .c(FE_OFN689_n_4438), .d(n_4444), .o(n_4354) );
na02m02 TIMEBOOST_cell_72117 ( .a(TIMEBOOST_net_23266), .b(g64113_sb), .o(n_4739) );
na02m01 TIMEBOOST_cell_37554 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q), .b(FE_OFN623_n_4409), .o(TIMEBOOST_net_10389) );
na02f06 g62312_u0 ( .a(n_1970), .b(n_2738), .o(g62312_p) );
in01f04 g62312_u1 ( .a(g62312_p), .o(n_2456) );
ao22f04 g62314_u0 ( .a(n_2264), .b(n_2727), .c(n_2711), .d(n_2430), .o(n_4197) );
oa12f01 g62316_u0 ( .a(n_5545), .b(n_5546), .c(pci_target_unit_fifos_pciw_inTransactionCount_1_), .o(n_5548) );
oa12f01 g62317_u0 ( .a(n_5545), .b(pci_target_unit_fifos_inGreyCount_0_), .c(n_5546), .o(n_5547) );
no02f01 g62318_u0 ( .a(n_1557), .b(n_4680), .o(g62318_p) );
in01f02 g62318_u1 ( .a(g62318_p), .o(n_4681) );
na02f01 g62319_u0 ( .a(n_3450), .b(n_4718), .o(g62319_p) );
in01f01 g62319_u1 ( .a(g62319_p), .o(n_4679) );
ao12f04 g62320_u0 ( .a(n_2956), .b(n_1445), .c(FE_OCP_RBN2239_g74749_p), .o(n_4165) );
ao12f02 g62321_u0 ( .a(n_3157), .b(n_1335), .c(wbm_rty_i), .o(n_3159) );
ao12s01 g62322_u0 ( .a(n_1714), .b(n_1226), .c(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(n_2034) );
in01s01 TIMEBOOST_cell_46005 ( .a(TIMEBOOST_net_13966), .o(TIMEBOOST_net_13863) );
oa12f01 g62325_u0 ( .a(n_7136), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_), .c(FE_OFN1192_n_6935), .o(n_7137) );
in01f01 g62326_u0 ( .a(FE_OFN1192_n_6935), .o(g62326_sb) );
na02s04 TIMEBOOST_cell_64016 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q), .o(TIMEBOOST_net_20994) );
na02f02 g62326_u2 ( .a(n_1510), .b(FE_OFN1192_n_6935), .o(g62326_db) );
na02f02 TIMEBOOST_cell_3266 ( .a(n_16495), .b(n_1774), .o(TIMEBOOST_net_193) );
ao12f02 g62327_u0 ( .a(n_3157), .b(n_2291), .c(wbm_rty_i), .o(n_3158) );
ao12f04 g62328_u0 ( .a(n_3157), .b(n_2396), .c(wbm_rty_i), .o(n_3156) );
ao12m06 g62329_u0 ( .a(n_1808), .b(n_4675), .c(n_4674), .o(n_4896) );
in01f02 g62330_u0 ( .a(n_7400), .o(n_7135) );
no02f04 g62331_u0 ( .a(n_4793), .b(n_3811), .o(n_7400) );
oa12f01 g62332_u0 ( .a(n_1099), .b(n_2728), .c(n_2959), .o(n_3333) );
in01f02 g62333_u0 ( .a(FE_OFN1269_n_4095), .o(g62333_sb) );
na02m02 TIMEBOOST_cell_68968 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q), .b(FE_OFN1643_n_4671), .o(TIMEBOOST_net_21692) );
na02m02 TIMEBOOST_cell_69756 ( .a(n_4444), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q), .o(TIMEBOOST_net_22086) );
in01m02 g62334_u0 ( .a(FE_OFN1269_n_4095), .o(g62334_sb) );
in01s01 TIMEBOOST_cell_73890 ( .a(n_8291), .o(TIMEBOOST_net_23455) );
na03f02 TIMEBOOST_cell_66516 ( .a(TIMEBOOST_net_16800), .b(FE_OFN1331_n_13547), .c(g53922_sb), .o(n_13522) );
in01s01 TIMEBOOST_cell_45974 ( .a(TIMEBOOST_net_13934), .o(TIMEBOOST_net_13935) );
in01f01 g62335_u0 ( .a(FE_OFN1275_n_4096), .o(g62335_sb) );
na02f02 TIMEBOOST_cell_71482 ( .a(n_1675), .b(FE_OFN1697_n_5751), .o(TIMEBOOST_net_22949) );
na03f02 TIMEBOOST_cell_73674 ( .a(TIMEBOOST_net_17507), .b(FE_OFN1233_n_6391), .c(g62532_sb), .o(n_6509) );
in01f02 g62336_u0 ( .a(FE_OFN1257_n_4143), .o(g62336_sb) );
na02s01 TIMEBOOST_cell_37452 ( .a(TIMEBOOST_net_23394), .b(g65691_sb), .o(TIMEBOOST_net_10338) );
na04m02 TIMEBOOST_cell_67829 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q), .b(n_8272), .c(n_1719), .d(g61903_sb), .o(n_8017) );
in01f02 g62337_u0 ( .a(FE_OFN1231_n_6391), .o(g62337_sb) );
na03s02 TIMEBOOST_cell_67907 ( .a(TIMEBOOST_net_7105), .b(FE_OFN775_n_15366), .c(g65893_sb), .o(n_2584) );
na02s02 TIMEBOOST_cell_53534 ( .a(TIMEBOOST_net_16984), .b(TIMEBOOST_net_12430), .o(TIMEBOOST_net_9416) );
in01f02 g62338_u0 ( .a(FE_OFN1231_n_6391), .o(g62338_sb) );
na03f02 TIMEBOOST_cell_66463 ( .a(TIMEBOOST_net_17017), .b(FE_OFN1224_n_6391), .c(g62517_sb), .o(n_6543) );
na02m06 TIMEBOOST_cell_71986 ( .a(FE_OFN636_n_4669), .b(n_4273), .o(TIMEBOOST_net_23201) );
na03f02 TIMEBOOST_cell_34742 ( .a(TIMEBOOST_net_9360), .b(FE_OFN1374_n_8567), .c(g57525_sb), .o(n_11216) );
in01f02 g62339_u0 ( .a(FE_OFN2064_n_6391), .o(g62339_sb) );
na02s02 TIMEBOOST_cell_44198 ( .a(TIMEBOOST_net_12993), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9473) );
in01f01 g62340_u0 ( .a(FE_OFN1275_n_4096), .o(g62340_sb) );
na03s02 TIMEBOOST_cell_67488 ( .a(TIMEBOOST_net_14674), .b(g58229_sb), .c(TIMEBOOST_net_14850), .o(TIMEBOOST_net_9538) );
in01f02 g62341_u0 ( .a(FE_OFN1295_n_4098), .o(g62341_sb) );
na02f02 TIMEBOOST_cell_72235 ( .a(TIMEBOOST_net_23325), .b(TIMEBOOST_net_14646), .o(TIMEBOOST_net_9341) );
na02f02 TIMEBOOST_cell_49766 ( .a(TIMEBOOST_net_15100), .b(g61902_sb), .o(n_8019) );
in01f02 g62342_u0 ( .a(FE_OFN1259_n_4143), .o(g62342_sb) );
na02m04 TIMEBOOST_cell_72119 ( .a(TIMEBOOST_net_23267), .b(FE_OFN923_n_4740), .o(TIMEBOOST_net_22282) );
na04f04 TIMEBOOST_cell_65120 ( .a(FE_OFN1655_n_9502), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q), .c(g58337_sb), .d(FE_OFN247_n_9112), .o(n_9019) );
in01m01 g62343_u0 ( .a(FE_OFN1219_n_6886), .o(g62343_sb) );
na02s01 TIMEBOOST_cell_44049 ( .a(FE_OFN554_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q), .o(TIMEBOOST_net_12919) );
na02s01 TIMEBOOST_cell_51541 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q), .o(TIMEBOOST_net_15988) );
in01f01 g62344_u0 ( .a(FE_OFN1275_n_4096), .o(g62344_sb) );
na03f02 TIMEBOOST_cell_66448 ( .a(TIMEBOOST_net_17121), .b(FE_OFN1314_n_6624), .c(g62666_sb), .o(n_6206) );
na02m01 TIMEBOOST_cell_68390 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q), .b(n_4677), .o(TIMEBOOST_net_21403) );
in01f02 g62345_u0 ( .a(FE_OFN1311_n_6624), .o(g62345_sb) );
na03f02 TIMEBOOST_cell_66498 ( .a(TIMEBOOST_net_17377), .b(FE_OFN1206_n_6356), .c(g62476_sb), .o(n_6636) );
na02f01 TIMEBOOST_cell_39481 ( .a(TIMEBOOST_net_11352), .b(g62836_sb), .o(n_5300) );
na03f02 TIMEBOOST_cell_73232 ( .a(TIMEBOOST_net_23364), .b(FE_OFN2084_n_8407), .c(g61780_sb), .o(n_8246) );
in01f02 g62346_u0 ( .a(FE_OFN1231_n_6391), .o(g62346_sb) );
na02f02 TIMEBOOST_cell_49918 ( .a(TIMEBOOST_net_15176), .b(g62737_sb), .o(TIMEBOOST_net_11340) );
na02s01 TIMEBOOST_cell_52416 ( .a(TIMEBOOST_net_16425), .b(FE_OFN201_n_9230), .o(TIMEBOOST_net_11461) );
na02m01 TIMEBOOST_cell_43097 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_133), .o(TIMEBOOST_net_12443) );
in01m02 g62347_u0 ( .a(FE_OFN1219_n_6886), .o(g62347_sb) );
na02s02 TIMEBOOST_cell_72021 ( .a(TIMEBOOST_net_23218), .b(g65704_sb), .o(n_1613) );
na03m02 TIMEBOOST_cell_69698 ( .a(FE_OFN1677_n_4655), .b(g65348_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q), .o(TIMEBOOST_net_22057) );
na04m04 TIMEBOOST_cell_72603 ( .a(TIMEBOOST_net_21471), .b(FE_OFN640_n_4669), .c(g65374_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q), .o(TIMEBOOST_net_17436) );
in01f02 g62348_u0 ( .a(n_6319), .o(g62348_sb) );
na02m10 TIMEBOOST_cell_53045 ( .a(configuration_pci_err_data_524), .b(wbm_dat_o_23_), .o(TIMEBOOST_net_16740) );
in01f02 g62349_u0 ( .a(FE_OFN1269_n_4095), .o(g62349_sb) );
na02s01 TIMEBOOST_cell_31845 ( .a(wbu_sel_in), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q), .o(TIMEBOOST_net_10027) );
na02m02 TIMEBOOST_cell_63157 ( .a(TIMEBOOST_net_20525), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_15531) );
na02s02 TIMEBOOST_cell_49297 ( .a(g58218_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_14866) );
in01f02 g62350_u0 ( .a(FE_OFN1278_n_4097), .o(g62350_sb) );
na03m02 TIMEBOOST_cell_64519 ( .a(n_3744), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q), .c(FE_OFN624_n_4409), .o(TIMEBOOST_net_10386) );
na03s02 TIMEBOOST_cell_65505 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q), .b(FE_OFN699_n_7845), .c(n_1903), .o(TIMEBOOST_net_14775) );
na03m04 TIMEBOOST_cell_72824 ( .a(g65053_sb), .b(n_17), .c(TIMEBOOST_net_16241), .o(TIMEBOOST_net_17556) );
in01f02 g62351_u0 ( .a(FE_OFN1322_n_6436), .o(g62351_sb) );
na02m02 TIMEBOOST_cell_70481 ( .a(TIMEBOOST_net_22448), .b(g59097_sb), .o(TIMEBOOST_net_670) );
in01f04 g62352_u0 ( .a(FE_OFN1250_n_4093), .o(g62352_sb) );
na04f10 TIMEBOOST_cell_20925 ( .a(n_1508), .b(pci_target_unit_wishbone_master_read_bound), .c(n_2000), .d(n_1535), .o(n_3304) );
na02m02 TIMEBOOST_cell_68275 ( .a(TIMEBOOST_net_21345), .b(TIMEBOOST_net_14157), .o(n_2213) );
na02m06 TIMEBOOST_cell_38842 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q), .b(n_13447), .o(TIMEBOOST_net_11033) );
in01f01 g62353_u0 ( .a(FE_OFN1261_n_4143), .o(g62353_sb) );
na03m02 TIMEBOOST_cell_67216 ( .a(FE_OFN562_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q), .c(TIMEBOOST_net_14358), .o(TIMEBOOST_net_9353) );
na03s02 TIMEBOOST_cell_46896 ( .a(TIMEBOOST_net_12957), .b(g58047_sb), .c(n_15569), .o(TIMEBOOST_net_9372) );
in01f01 g62354_u0 ( .a(FE_OFN1261_n_4143), .o(g62354_sb) );
na03f02 TIMEBOOST_cell_34921 ( .a(TIMEBOOST_net_9492), .b(FE_OFN1380_n_8567), .c(g57304_sb), .o(n_10404) );
in01f02 g62355_u0 ( .a(FE_OFN1232_n_6391), .o(g62355_sb) );
na04f04 TIMEBOOST_cell_73313 ( .a(n_3906), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q), .c(FE_OFN1132_g64577_p), .d(g63119_sb), .o(n_5018) );
in01m01 g62356_u0 ( .a(FE_OFN1218_n_6886), .o(g62356_sb) );
in01f02 g62357_u0 ( .a(FE_OFN1284_n_4097), .o(g62357_sb) );
na02s02 TIMEBOOST_cell_25329 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_73), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6769) );
na02s01 TIMEBOOST_cell_42892 ( .a(TIMEBOOST_net_12340), .b(FE_OFN941_n_2047), .o(TIMEBOOST_net_10354) );
na02s01 TIMEBOOST_cell_42894 ( .a(TIMEBOOST_net_12341), .b(FE_OFN941_n_2047), .o(TIMEBOOST_net_10339) );
in01f02 g62358_u0 ( .a(FE_OFN1273_n_4096), .o(g62358_sb) );
no03f10 TIMEBOOST_cell_20929 ( .a(FE_RN_428_0), .b(FE_RN_764_0), .c(FE_RN_430_0), .o(FE_RN_462_0) );
na03f02 TIMEBOOST_cell_67092 ( .a(FE_OFN1596_n_13741), .b(n_13903), .c(TIMEBOOST_net_13800), .o(n_14428) );
in01f02 g62359_u0 ( .a(FE_OFN1216_n_4151), .o(g62359_sb) );
na02f01 TIMEBOOST_cell_48124 ( .a(TIMEBOOST_net_14279), .b(g66001_db), .o(n_2147) );
na03f02 TIMEBOOST_cell_47290 ( .a(FE_OFN1734_n_16317), .b(TIMEBOOST_net_13586), .c(FE_OFN1739_n_11019), .o(n_12607) );
na02m02 TIMEBOOST_cell_38618 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q), .b(g65401_sb), .o(TIMEBOOST_net_10921) );
in01f02 g62360_u0 ( .a(FE_OFN1282_n_4097), .o(g62360_sb) );
na02m02 TIMEBOOST_cell_49760 ( .a(TIMEBOOST_net_15097), .b(g61878_sb), .o(n_8073) );
na02s01 TIMEBOOST_cell_49231 ( .a(FE_OFN1021_n_11877), .b(wbu_addr_in_269), .o(TIMEBOOST_net_14833) );
na02f01 TIMEBOOST_cell_68050 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q), .b(n_8831), .o(TIMEBOOST_net_21233) );
in01f01 g62361_u0 ( .a(FE_OFN1246_n_4093), .o(g62361_sb) );
in01f01 g62362_u0 ( .a(FE_OFN1274_n_4096), .o(g62362_sb) );
na02m01 TIMEBOOST_cell_51931 ( .a(n_4677), .b(n_3764), .o(TIMEBOOST_net_16183) );
in01f02 g62363_u0 ( .a(n_6431), .o(g62363_sb) );
in01s06 TIMEBOOST_cell_67734 ( .a(TIMEBOOST_net_21161), .o(TIMEBOOST_net_21160) );
na04m02 TIMEBOOST_cell_72709 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q), .b(g64854_sb), .c(FE_OFN1626_n_4438), .d(TIMEBOOST_net_20355), .o(TIMEBOOST_net_13374) );
in01f02 g62364_u0 ( .a(FE_OFN1258_n_4143), .o(g62364_sb) );
na03s02 TIMEBOOST_cell_72507 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q), .b(FE_OFN517_n_9697), .c(TIMEBOOST_net_14178), .o(TIMEBOOST_net_12982) );
na04f06 TIMEBOOST_cell_42134 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q), .b(g63533_sb), .c(g63533_db), .d(TIMEBOOST_net_625), .o(n_5642) );
na02f04 TIMEBOOST_cell_51671 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q), .b(FE_OCP_RBN1976_n_12381), .o(TIMEBOOST_net_16053) );
in01f02 g62365_u0 ( .a(FE_OFN1222_n_6391), .o(g62365_sb) );
na02m01 TIMEBOOST_cell_62812 ( .a(n_3792), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q), .o(TIMEBOOST_net_20353) );
na03f02 TIMEBOOST_cell_66412 ( .a(n_3846), .b(g63126_sb), .c(g63126_db), .o(n_5001) );
in01m01 g62366_u0 ( .a(FE_OFN1192_n_6935), .o(g62366_sb) );
na02f10 TIMEBOOST_cell_3271 ( .a(TIMEBOOST_net_195), .b(n_2562), .o(n_3388) );
na02f01 g62366_u2 ( .a(n_3765), .b(FE_OFN1192_n_6935), .o(g62366_db) );
na04s02 TIMEBOOST_cell_72905 ( .a(TIMEBOOST_net_12493), .b(g65694_sb), .c(g61775_sb), .d(g61775_db), .o(n_8258) );
in01f02 g62367_u0 ( .a(FE_OFN2063_n_6391), .o(g62367_sb) );
na02s01 TIMEBOOST_cell_45445 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q), .o(TIMEBOOST_net_13617) );
na04f02 TIMEBOOST_cell_73462 ( .a(n_3721), .b(FE_OFN1222_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q), .d(g62513_sb), .o(n_6553) );
in01f02 g62368_u0 ( .a(n_6287), .o(g62368_sb) );
na02f02 TIMEBOOST_cell_26215 ( .a(conf_wb_err_addr_in_956), .b(g53937_sb), .o(TIMEBOOST_net_7212) );
na02f02 TIMEBOOST_cell_49854 ( .a(TIMEBOOST_net_15144), .b(g62838_sb), .o(n_5298) );
in01f02 g62369_u0 ( .a(FE_OFN1293_n_4098), .o(g62369_sb) );
na02m02 TIMEBOOST_cell_53581 ( .a(n_4359), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q), .o(TIMEBOOST_net_17008) );
na03m02 TIMEBOOST_cell_65076 ( .a(n_3785), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q), .c(FE_OFN619_n_4490), .o(TIMEBOOST_net_16237) );
na03f02 TIMEBOOST_cell_67984 ( .a(TIMEBOOST_net_20956), .b(FE_OFN1293_n_4098), .c(g62369_sb), .o(n_6865) );
in01f02 g62370_u0 ( .a(FE_OFN1230_n_6391), .o(g62370_sb) );
na02m04 TIMEBOOST_cell_26207 ( .a(FE_OFN2071_n_15978), .b(conf_wb_err_addr_in_953), .o(TIMEBOOST_net_7208) );
na03f02 TIMEBOOST_cell_72733 ( .a(TIMEBOOST_net_14311), .b(FE_OFN2108_n_2047), .c(TIMEBOOST_net_17246), .o(TIMEBOOST_net_14593) );
na03f02 TIMEBOOST_cell_67035 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_16534), .c(FE_OFN1600_n_13995), .o(n_14448) );
in01f01 g62371_u0 ( .a(FE_OFN1194_n_6935), .o(g62371_sb) );
in01s01 TIMEBOOST_cell_67784 ( .a(TIMEBOOST_net_21210), .o(TIMEBOOST_net_21211) );
na03f02 TIMEBOOST_cell_67983 ( .a(TIMEBOOST_net_20978), .b(FE_OFN1293_n_4098), .c(g62962_sb), .o(n_5958) );
in01f01 g62372_u0 ( .a(FE_OFN1284_n_4097), .o(g62372_sb) );
na02s01 TIMEBOOST_cell_48128 ( .a(TIMEBOOST_net_14281), .b(g58195_sb), .o(TIMEBOOST_net_12491) );
na03f02 TIMEBOOST_cell_73719 ( .a(n_12001), .b(TIMEBOOST_net_13556), .c(FE_OFN1746_n_12004), .o(n_12666) );
in01m01 g62373_u0 ( .a(FE_OFN1295_n_4098), .o(g62373_sb) );
in01f02 g62374_u0 ( .a(FE_OFN1207_n_6356), .o(g62374_sb) );
na04f02 TIMEBOOST_cell_73622 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q), .b(n_8747), .c(TIMEBOOST_net_9976), .d(g58633_sb), .o(n_8848) );
na03m02 TIMEBOOST_cell_72470 ( .a(TIMEBOOST_net_16571), .b(FE_OFN903_n_4736), .c(g64219_sb), .o(TIMEBOOST_net_13113) );
in01m02 g62375_u0 ( .a(FE_OFN1269_n_4095), .o(g62375_sb) );
na02m02 TIMEBOOST_cell_70745 ( .a(TIMEBOOST_net_22580), .b(g61724_sb), .o(n_8373) );
na03f04 TIMEBOOST_cell_64345 ( .a(n_15755), .b(wbu_map_in_132), .c(n_15065), .o(n_2389) );
na03f02 TIMEBOOST_cell_73675 ( .a(TIMEBOOST_net_17369), .b(FE_OFN1258_n_4143), .c(g62537_sb), .o(n_6495) );
in01f01 g62376_u0 ( .a(FE_OFN1261_n_4143), .o(g62376_sb) );
na02s01 TIMEBOOST_cell_64196 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q), .o(TIMEBOOST_net_21084) );
na02f02 TIMEBOOST_cell_3219 ( .a(TIMEBOOST_net_169), .b(FE_OFN1071_n_15729), .o(n_3084) );
na02s01 TIMEBOOST_cell_30855 ( .a(n_9786), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q), .o(TIMEBOOST_net_9532) );
in01f02 g62377_u0 ( .a(FE_OFN1260_n_4143), .o(g62377_sb) );
na04f04 TIMEBOOST_cell_24954 ( .a(n_10112), .b(n_10116), .c(n_9295), .d(n_9294), .o(n_11847) );
in01f02 g62378_u0 ( .a(FE_OFN1231_n_6391), .o(g62378_sb) );
na02m02 TIMEBOOST_cell_72116 ( .a(TIMEBOOST_net_17249), .b(FE_OFN1049_n_16657), .o(TIMEBOOST_net_23266) );
na03f02 TIMEBOOST_cell_35055 ( .a(TIMEBOOST_net_9607), .b(FE_OFN1439_n_9372), .c(g58474_sb), .o(n_9368) );
in01f02 g62379_u0 ( .a(FE_OFN1230_n_6391), .o(g62379_sb) );
na03f02 TIMEBOOST_cell_35054 ( .a(TIMEBOOST_net_9606), .b(FE_OFN1436_n_9372), .c(g58460_sb), .o(n_8986) );
in01m02 g62380_u0 ( .a(FE_OFN1269_n_4095), .o(g62380_sb) );
na02m01 TIMEBOOST_cell_52148 ( .a(TIMEBOOST_net_16291), .b(g65811_sb), .o(n_1903) );
na04f04 TIMEBOOST_cell_24848 ( .a(wbs_dat_o_20_), .b(g52516_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_119), .d(FE_OFN1472_g52675_p), .o(n_13709) );
na04f04 TIMEBOOST_cell_24850 ( .a(wbs_dat_o_11_), .b(g52505_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_110), .d(FE_OFN2243_g52675_p), .o(n_13822) );
in01f02 g62381_u0 ( .a(FE_OFN2064_n_6391), .o(g62381_sb) );
na02m04 TIMEBOOST_cell_26213 ( .a(g53897_sb), .b(conf_wb_err_addr_in_959), .o(TIMEBOOST_net_7211) );
na03m04 TIMEBOOST_cell_72756 ( .a(n_4476), .b(n_4429), .c(TIMEBOOST_net_12691), .o(TIMEBOOST_net_20583) );
na04f02 TIMEBOOST_cell_73124 ( .a(g64277_da), .b(g64277_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q), .d(FE_OFN1140_g64577_p), .o(TIMEBOOST_net_22456) );
in01f02 g62382_u0 ( .a(n_6554), .o(g62382_sb) );
na02m01 TIMEBOOST_cell_52328 ( .a(TIMEBOOST_net_16381), .b(FE_OFN2021_n_4778), .o(n_7195) );
in01s01 TIMEBOOST_cell_73980 ( .a(n_8843), .o(TIMEBOOST_net_23545) );
na02m08 TIMEBOOST_cell_45625 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q), .o(TIMEBOOST_net_13707) );
in01m01 g62383_u0 ( .a(FE_OFN1218_n_6886), .o(g62383_sb) );
na02m10 TIMEBOOST_cell_52981 ( .a(wishbone_slave_unit_pcim_sm_data_in_638), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q), .o(TIMEBOOST_net_16708) );
na04f04 TIMEBOOST_cell_24852 ( .a(wbs_dat_o_10_), .b(g52503_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_109), .d(FE_OFN2243_g52675_p), .o(n_13823) );
na02m02 g54203_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_11__Q), .b(n_13221), .o(g54203_db) );
in01f01 g62384_u0 ( .a(FE_OFN1284_n_4097), .o(g62384_sb) );
na02f02 TIMEBOOST_cell_50264 ( .a(TIMEBOOST_net_15349), .b(g62343_sb), .o(n_6913) );
na02f08 TIMEBOOST_cell_71833 ( .a(TIMEBOOST_net_23124), .b(parchk_pci_cbe_out_in_1204), .o(n_2566) );
na04f04 TIMEBOOST_cell_24854 ( .a(wbs_dat_o_19_), .b(g52513_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_118), .d(FE_OFN2243_g52675_p), .o(n_13812) );
in01f01 g62385_u0 ( .a(FE_OFN1285_n_4097), .o(g62385_sb) );
na04f04 TIMEBOOST_cell_24856 ( .a(wbs_dat_o_17_), .b(g52511_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_116), .d(FE_OFN2243_g52675_p), .o(n_13712) );
na04f04 TIMEBOOST_cell_24858 ( .a(wbs_dat_o_14_), .b(g52508_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_113), .d(FE_OFN2242_g52675_p), .o(n_13717) );
in01f01 g62386_u0 ( .a(FE_OFN1261_n_4143), .o(g62386_sb) );
na02m01 TIMEBOOST_cell_37532 ( .a(n_3783), .b(n_4671), .o(TIMEBOOST_net_10378) );
na03m02 TIMEBOOST_cell_68696 ( .a(TIMEBOOST_net_20207), .b(FE_OFN916_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q), .o(TIMEBOOST_net_21556) );
in01f01 g62387_u0 ( .a(FE_OFN1273_n_4096), .o(g62387_sb) );
na02f06 TIMEBOOST_cell_3245 ( .a(TIMEBOOST_net_182), .b(n_3013), .o(n_3359) );
na02f02 TIMEBOOST_cell_72121 ( .a(TIMEBOOST_net_23268), .b(FE_OFN923_n_4740), .o(TIMEBOOST_net_22291) );
in01f02 g62388_u0 ( .a(FE_OFN1213_n_4151), .o(g62388_sb) );
na04f02 TIMEBOOST_cell_73623 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q), .b(n_8747), .c(TIMEBOOST_net_9977), .d(g58635_sb), .o(n_8847) );
in01f01 g62389_u0 ( .a(FE_OFN1212_n_4151), .o(g62389_sb) );
in01s01 TIMEBOOST_cell_63535 ( .a(TIMEBOOST_net_20715), .o(TIMEBOOST_net_20714) );
na03f02 TIMEBOOST_cell_33522 ( .a(TIMEBOOST_net_8784), .b(FE_OFN1168_n_5592), .c(g62093_sb), .o(n_5612) );
na02m06 TIMEBOOST_cell_69350 ( .a(g65301_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q), .o(TIMEBOOST_net_21883) );
in01m01 g62390_u0 ( .a(FE_OFN1279_n_4097), .o(g62390_sb) );
na03f02 TIMEBOOST_cell_73510 ( .a(TIMEBOOST_net_13376), .b(n_6287), .c(g62911_sb), .o(n_6056) );
na02m02 TIMEBOOST_cell_38192 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q), .b(g65283_sb), .o(TIMEBOOST_net_10708) );
in01f01 g62391_u0 ( .a(FE_OFN1285_n_4097), .o(g62391_sb) );
na04f04 TIMEBOOST_cell_36850 ( .a(n_9022), .b(g57471_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q), .d(FE_OFN1391_n_8567), .o(n_10342) );
na04f02 TIMEBOOST_cell_24872 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q), .b(g54485_sb), .c(n_13608), .d(n_13617), .o(n_13614) );
na02m02 TIMEBOOST_cell_68697 ( .a(TIMEBOOST_net_21556), .b(g64363_sb), .o(TIMEBOOST_net_13055) );
in01f01 g62392_u0 ( .a(FE_OFN1208_n_6356), .o(g62392_sb) );
na02s01 TIMEBOOST_cell_31843 ( .a(wbu_sel_in_313), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q), .o(TIMEBOOST_net_10026) );
na03f02 TIMEBOOST_cell_24876 ( .a(FE_RN_89_0), .b(n_10644), .c(n_12575), .o(n_12837) );
in01f01 g62393_u0 ( .a(FE_OFN1250_n_4093), .o(g62393_sb) );
na03f02 TIMEBOOST_cell_73819 ( .a(n_13891), .b(TIMEBOOST_net_16554), .c(FE_OFN1593_n_13741), .o(g53258_p) );
na02m01 TIMEBOOST_cell_68644 ( .a(FE_OFN667_n_4495), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q), .o(TIMEBOOST_net_21530) );
in01f01 g62394_u0 ( .a(FE_OFN1275_n_4096), .o(g62394_sb) );
na02m02 TIMEBOOST_cell_50020 ( .a(TIMEBOOST_net_15227), .b(TIMEBOOST_net_11462), .o(TIMEBOOST_net_9379) );
na03f02 TIMEBOOST_cell_73660 ( .a(TIMEBOOST_net_14890), .b(FE_OFN1094_g64577_p), .c(g63048_sb), .o(n_5156) );
na04m04 TIMEBOOST_cell_67215 ( .a(g65008_sb), .b(FE_OFN1625_n_4438), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q), .d(n_4447), .o(n_4349) );
in01f02 g62395_u0 ( .a(FE_OFN1316_n_6624), .o(g62395_sb) );
na03f02 TIMEBOOST_cell_73780 ( .a(TIMEBOOST_net_8111), .b(n_13987), .c(FE_OFN1589_n_13736), .o(n_16252) );
in01f02 g62396_u0 ( .a(n_6431), .o(g62396_sb) );
na02f02 TIMEBOOST_cell_27019 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_8__Q), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_7614) );
na02m02 TIMEBOOST_cell_50598 ( .a(TIMEBOOST_net_15516), .b(g62582_sb), .o(n_6388) );
na02m02 TIMEBOOST_cell_68274 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(g65674_sb), .o(TIMEBOOST_net_21345) );
in01f01 g62397_u0 ( .a(FE_OFN1214_n_4151), .o(g62397_sb) );
na03f02 TIMEBOOST_cell_73390 ( .a(TIMEBOOST_net_16726), .b(FE_OFN1184_n_3476), .c(g60643_sb), .o(n_5686) );
na03m02 TIMEBOOST_cell_72658 ( .a(n_3755), .b(FE_OFN644_n_4677), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q), .o(TIMEBOOST_net_22122) );
in01f02 g62398_u0 ( .a(FE_OFN1260_n_4143), .o(g62398_sb) );
na04f04 TIMEBOOST_cell_36706 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q), .b(g53927_sb), .c(n_13166), .d(FE_OFN1327_n_13547), .o(n_13518) );
na03f02 TIMEBOOST_cell_66205 ( .a(TIMEBOOST_net_20969), .b(FE_OFN1200_n_4090), .c(g63094_sb), .o(n_5856) );
na02f02 TIMEBOOST_cell_70836 ( .a(TIMEBOOST_net_16698), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_22626) );
in01m01 g62399_u0 ( .a(FE_OFN1193_n_6935), .o(g62399_sb) );
na02f02 TIMEBOOST_cell_52934 ( .a(TIMEBOOST_net_16684), .b(g63097_sb), .o(n_5060) );
na02s01 TIMEBOOST_cell_48573 ( .a(FE_OFN219_n_9853), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q), .o(TIMEBOOST_net_14504) );
na02s02 TIMEBOOST_cell_48571 ( .a(FE_OFN223_n_9844), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q), .o(TIMEBOOST_net_14503) );
in01f02 g62400_u0 ( .a(n_6645), .o(g62400_sb) );
na03f02 TIMEBOOST_cell_73511 ( .a(TIMEBOOST_net_13372), .b(n_6287), .c(g62664_sb), .o(n_6211) );
na02s01 TIMEBOOST_cell_44201 ( .a(g57911_sb), .b(g57911_db), .o(TIMEBOOST_net_12995) );
na04f04 TIMEBOOST_cell_67658 ( .a(TIMEBOOST_net_7548), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q), .c(FE_OFN1248_n_4093), .d(g62918_sb), .o(n_6043) );
in01f02 g62401_u0 ( .a(FE_OFN1313_n_6624), .o(g62401_sb) );
na02m01 TIMEBOOST_cell_69620 ( .a(n_4645), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q), .o(TIMEBOOST_net_22018) );
na02s02 TIMEBOOST_cell_39799 ( .a(g58438_db), .b(TIMEBOOST_net_11511), .o(n_9201) );
in01f02 g62402_u0 ( .a(FE_OFN1236_n_6391), .o(g62402_sb) );
na02m10 TIMEBOOST_cell_45243 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q), .o(TIMEBOOST_net_13516) );
na02f02 TIMEBOOST_cell_71129 ( .a(TIMEBOOST_net_22772), .b(g62440_sb), .o(n_6716) );
na02f06 TIMEBOOST_cell_71835 ( .a(TIMEBOOST_net_23125), .b(parchk_pci_cbe_out_in_1203), .o(n_2171) );
in01f02 g62403_u0 ( .a(FE_OFN1232_n_6391), .o(g62403_sb) );
na02f10 TIMEBOOST_cell_69682 ( .a(n_13763), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_394), .o(TIMEBOOST_net_22049) );
no03f02 TIMEBOOST_cell_3482 ( .a(n_1635), .b(n_1697), .c(g59232_BP), .o(TIMEBOOST_net_301) );
in01f02 g62404_u0 ( .a(n_6319), .o(g62404_sb) );
na02m02 TIMEBOOST_cell_63327 ( .a(TIMEBOOST_net_20610), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_15496) );
na04f02 TIMEBOOST_cell_36837 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q), .b(FE_OFN1394_n_8567), .c(n_9130), .d(g57063_sb), .o(n_10503) );
na03f02 TIMEBOOST_cell_34865 ( .a(TIMEBOOST_net_9329), .b(FE_OFN1400_n_8567), .c(g57206_sb), .o(n_11551) );
in01m01 g62405_u0 ( .a(FE_OFN1219_n_6886), .o(g62405_sb) );
na02s01 TIMEBOOST_cell_69783 ( .a(TIMEBOOST_net_22099), .b(FE_OFN215_n_9856), .o(TIMEBOOST_net_17015) );
na02s02 TIMEBOOST_cell_48567 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q), .o(TIMEBOOST_net_14501) );
na02s02 TIMEBOOST_cell_48563 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q), .o(TIMEBOOST_net_14499) );
in01f02 g62406_u0 ( .a(FE_OFN1235_n_6391), .o(g62406_sb) );
no02f02 TIMEBOOST_cell_3483 ( .a(TIMEBOOST_net_301), .b(n_7715), .o(g59232_p) );
na02s02 TIMEBOOST_cell_3484 ( .a(pci_target_unit_del_sync_comp_cycle_count_14_), .b(pci_target_unit_del_sync_comp_cycle_count_15_), .o(TIMEBOOST_net_302) );
in01f02 g62407_u0 ( .a(FE_OFN1310_n_6624), .o(g62407_sb) );
na03f02 TIMEBOOST_cell_73055 ( .a(TIMEBOOST_net_22030), .b(FE_OFN2084_n_8407), .c(g61819_sb), .o(n_8152) );
na02f02 TIMEBOOST_cell_3741 ( .a(TIMEBOOST_net_430), .b(n_17049), .o(n_4881) );
in01s01 TIMEBOOST_cell_73947 ( .a(TIMEBOOST_net_23511), .o(TIMEBOOST_net_23512) );
in01f02 g62408_u0 ( .a(FE_OFN1310_n_6624), .o(g62408_sb) );
na02m02 TIMEBOOST_cell_53418 ( .a(TIMEBOOST_net_16926), .b(g64158_sb), .o(TIMEBOOST_net_8797) );
na02f02 TIMEBOOST_cell_3743 ( .a(TIMEBOOST_net_431), .b(n_17040), .o(n_4878) );
na03f02 TIMEBOOST_cell_65513 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q), .b(FE_OFN714_n_8140), .c(n_1946), .o(TIMEBOOST_net_14872) );
in01f04 g62409_u0 ( .a(FE_OFN1234_n_6391), .o(g62409_sb) );
na02f06 TIMEBOOST_cell_3485 ( .a(n_3025), .b(TIMEBOOST_net_302), .o(n_3463) );
na02s02 TIMEBOOST_cell_3486 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q), .o(TIMEBOOST_net_303) );
in01m01 g62410_u0 ( .a(FE_OFN1270_n_4095), .o(g62410_sb) );
na03f02 TIMEBOOST_cell_73233 ( .a(TIMEBOOST_net_23363), .b(FE_OFN2084_n_8407), .c(g61788_sb), .o(n_8226) );
na02f04 TIMEBOOST_cell_51672 ( .a(n_16402), .b(TIMEBOOST_net_16053), .o(n_16403) );
in01f01 g62411_u0 ( .a(FE_OFN1272_n_4096), .o(g62411_sb) );
na02s01 TIMEBOOST_cell_43443 ( .a(pci_target_unit_fifos_pcir_data_in), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q), .o(TIMEBOOST_net_12616) );
in01f01 g62412_u0 ( .a(FE_OFN1202_n_4090), .o(g62412_sb) );
na02f02 TIMEBOOST_cell_28006 ( .a(n_13901), .b(TIMEBOOST_net_8107), .o(TIMEBOOST_net_762) );
na04f04 TIMEBOOST_cell_24657 ( .a(n_9726), .b(g57207_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q), .d(FE_OFN1427_n_8567), .o(n_11549) );
in01f01 g62413_u0 ( .a(FE_OFN1253_n_4143), .o(g62413_sb) );
na04f04 TIMEBOOST_cell_24659 ( .a(n_9223), .b(g57199_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q), .d(FE_OFN1427_n_8567), .o(n_10835) );
na02s02 TIMEBOOST_cell_38551 ( .a(TIMEBOOST_net_10887), .b(g57945_db), .o(n_9867) );
in01f01 g62414_u0 ( .a(FE_OFN1214_n_4151), .o(g62414_sb) );
na02s01 TIMEBOOST_cell_68192 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q), .b(g65907_db), .o(TIMEBOOST_net_21304) );
na03f02 TIMEBOOST_cell_73661 ( .a(TIMEBOOST_net_13058), .b(FE_OFN1118_g64577_p), .c(g63030_sb), .o(n_5188) );
in01m01 g62415_u0 ( .a(FE_OFN1219_n_6886), .o(g62415_sb) );
na02m01 TIMEBOOST_cell_68512 ( .a(pci_target_unit_del_sync_addr_in_223), .b(g66397_sb), .o(TIMEBOOST_net_21464) );
in01s04 TIMEBOOST_cell_17853 ( .a(TIMEBOOST_net_5264), .o(n_3280) );
in01f02 g62416_u0 ( .a(FE_OFN1316_n_6624), .o(g62416_sb) );
na03f02 TIMEBOOST_cell_47292 ( .a(FE_OFN1736_n_16317), .b(TIMEBOOST_net_13588), .c(FE_OFN1742_n_11019), .o(n_12613) );
in01s01 TIMEBOOST_cell_72354 ( .a(pci_target_unit_fifos_pcir_data_in_167), .o(TIMEBOOST_net_23387) );
na03m02 TIMEBOOST_cell_64518 ( .a(n_3749), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q), .c(FE_OFN682_n_4460), .o(TIMEBOOST_net_10541) );
in01f02 g62417_u0 ( .a(FE_OFN1253_n_4143), .o(g62417_sb) );
na02m04 TIMEBOOST_cell_68742 ( .a(FE_OFN660_n_4392), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q), .o(TIMEBOOST_net_21579) );
na04f04 TIMEBOOST_cell_24590 ( .a(n_9488), .b(g57464_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q), .d(FE_OFN2177_n_8567), .o(n_11268) );
in01m01 g62418_u0 ( .a(FE_OFN1241_n_4092), .o(g62418_sb) );
na04f04 TIMEBOOST_cell_24592 ( .a(n_9431), .b(g57450_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q), .d(FE_OFN2168_n_8567), .o(n_11284) );
na04f04 TIMEBOOST_cell_24594 ( .a(n_8553), .b(g58595_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q), .d(FE_OFN2184_n_8567), .o(n_8957) );
in01f01 g62419_u0 ( .a(FE_OFN1243_n_4092), .o(g62419_sb) );
na03m02 TIMEBOOST_cell_65184 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q), .b(g64289_sb), .c(TIMEBOOST_net_14667), .o(TIMEBOOST_net_13060) );
na04f04 TIMEBOOST_cell_24596 ( .a(n_9405), .b(g57594_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q), .d(FE_OFN1427_n_8567), .o(n_11159) );
na04f04 TIMEBOOST_cell_24598 ( .a(n_9200), .b(g57586_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q), .d(FE_OFN2170_n_8567), .o(n_10799) );
in01f01 g62420_u0 ( .a(FE_OFN1268_n_4095), .o(g62420_sb) );
na02m02 TIMEBOOST_cell_38317 ( .a(TIMEBOOST_net_10770), .b(g58389_db), .o(n_9007) );
na04f04 TIMEBOOST_cell_24600 ( .a(n_9419), .b(g57573_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q), .d(FE_OFN2180_n_8567), .o(n_11178) );
na04f04 TIMEBOOST_cell_24558 ( .a(n_9206), .b(g57553_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q), .d(FE_OFN1416_n_8567), .o(n_10807) );
in01f02 g62421_u0 ( .a(n_6554), .o(g62421_sb) );
na02m01 TIMEBOOST_cell_68196 ( .a(n_2299), .b(TIMEBOOST_net_12338), .o(TIMEBOOST_net_21306) );
na02f01 TIMEBOOST_cell_63027 ( .a(TIMEBOOST_net_20460), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_15189) );
na02s01 TIMEBOOST_cell_48813 ( .a(FE_OFN235_n_9834), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_14624) );
in01f01 g62422_u0 ( .a(FE_OFN1244_n_4092), .o(g62422_sb) );
na04f04 TIMEBOOST_cell_24602 ( .a(n_9426), .b(g57563_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q), .d(FE_OFN2188_n_8567), .o(n_11188) );
na04f04 TIMEBOOST_cell_24622 ( .a(n_9872), .b(g57058_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q), .d(FE_OFN2174_n_8567), .o(n_11679) );
in01m01 g62423_u0 ( .a(FE_OFN1224_n_6391), .o(g62423_sb) );
na02f02 TIMEBOOST_cell_70247 ( .a(TIMEBOOST_net_22331), .b(g61841_sb), .o(n_6969) );
in01f02 g62424_u0 ( .a(FE_OFN1252_n_4143), .o(g62424_sb) );
na02f01 TIMEBOOST_cell_37212 ( .a(TIMEBOOST_net_5353), .b(n_1813), .o(TIMEBOOST_net_10218) );
na04f04 TIMEBOOST_cell_24624 ( .a(n_9110), .b(g57109_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q), .d(FE_OFN2167_n_8567), .o(n_10478) );
na02s01 g58449_u2 ( .a(FE_OFN233_n_9876), .b(FE_OFN1648_n_9428), .o(g58449_db) );
in01f02 g62425_u0 ( .a(FE_OFN1311_n_6624), .o(g62425_sb) );
na03f02 TIMEBOOST_cell_34864 ( .a(TIMEBOOST_net_9511), .b(FE_OFN1385_n_8567), .c(g57053_sb), .o(n_11683) );
na03s01 TIMEBOOST_cell_69170 ( .a(g61924_sb), .b(g61924_db), .c(g65865_db), .o(TIMEBOOST_net_21793) );
na02m01 TIMEBOOST_cell_52183 ( .a(configuration_wb_err_cs_bit_569), .b(parchk_pci_cbe_out_in_1203), .o(TIMEBOOST_net_16309) );
in01f02 g62426_u0 ( .a(FE_OFN1223_n_6391), .o(g62426_sb) );
na02f02 TIMEBOOST_cell_71081 ( .a(TIMEBOOST_net_22748), .b(g62412_sb), .o(n_6774) );
na02f02 TIMEBOOST_cell_53622 ( .a(TIMEBOOST_net_17028), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_15477) );
na02f08 TIMEBOOST_cell_3276 ( .a(n_2681), .b(n_2680), .o(TIMEBOOST_net_198) );
in01f02 g62427_u0 ( .a(FE_OFN1316_n_6624), .o(g62427_sb) );
na03m02 TIMEBOOST_cell_65737 ( .a(TIMEBOOST_net_20856), .b(n_1585), .c(g61927_sb), .o(n_7969) );
na02f02 TIMEBOOST_cell_69445 ( .a(TIMEBOOST_net_21930), .b(TIMEBOOST_net_14434), .o(TIMEBOOST_net_17133) );
na02f02 TIMEBOOST_cell_3750 ( .a(n_7712), .b(n_8452), .o(TIMEBOOST_net_435) );
in01f01 g62428_u0 ( .a(FE_OFN1224_n_6391), .o(g62428_sb) );
na02f06 TIMEBOOST_cell_3277 ( .a(TIMEBOOST_net_198), .b(n_2461), .o(n_2991) );
na04f04 TIMEBOOST_cell_24174 ( .a(n_9509), .b(g57436_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q), .d(FE_OFN1402_n_8567), .o(n_11300) );
in01m01 g62429_u0 ( .a(FE_OFN1219_n_6886), .o(g62429_sb) );
na02f02 TIMEBOOST_cell_40617 ( .a(TIMEBOOST_net_11920), .b(n_12858), .o(n_14806) );
na02s01 g58445_u2 ( .a(FE_OFN254_n_9825), .b(FE_OFN523_n_9428), .o(g58445_db) );
na03f02 TIMEBOOST_cell_66854 ( .a(TIMEBOOST_net_17588), .b(n_14971), .c(g58655_sb), .o(n_9234) );
in01m02 g62430_u0 ( .a(FE_OFN1269_n_4095), .o(g62430_sb) );
na03m02 TIMEBOOST_cell_73036 ( .a(TIMEBOOST_net_12606), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q), .c(TIMEBOOST_net_8728), .o(TIMEBOOST_net_17390) );
na02m01 TIMEBOOST_cell_47883 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN938_n_2292), .o(TIMEBOOST_net_14159) );
na02s02 TIMEBOOST_cell_47923 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q), .b(pci_target_unit_fifos_pcir_data_in_164), .o(TIMEBOOST_net_14179) );
in01f02 g62431_u0 ( .a(FE_OFN2063_n_6391), .o(g62431_sb) );
na02f06 TIMEBOOST_cell_3487 ( .a(TIMEBOOST_net_303), .b(n_3074), .o(n_3462) );
na03s02 TIMEBOOST_cell_72685 ( .a(TIMEBOOST_net_14151), .b(g65878_db), .c(TIMEBOOST_net_20340), .o(n_7879) );
in01f02 g62432_u0 ( .a(FE_OFN1235_n_6391), .o(g62432_sb) );
na03m04 TIMEBOOST_cell_72686 ( .a(g64999_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q), .c(TIMEBOOST_net_10567), .o(TIMEBOOST_net_20579) );
na03m02 TIMEBOOST_cell_68804 ( .a(TIMEBOOST_net_20213), .b(FE_OFN916_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_21610) );
in01f04 g62433_u0 ( .a(FE_OFN1313_n_6624), .o(g62433_sb) );
na02f06 TIMEBOOST_cell_3751 ( .a(TIMEBOOST_net_435), .b(n_16167), .o(n_12956) );
na02f02 TIMEBOOST_cell_70557 ( .a(TIMEBOOST_net_22486), .b(g62812_sb), .o(n_5354) );
in01f02 g62434_u0 ( .a(n_6554), .o(g62434_sb) );
na04m02 TIMEBOOST_cell_73234 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(g64109_sb), .c(TIMEBOOST_net_16411), .d(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q), .o(TIMEBOOST_net_22420) );
na02s01 TIMEBOOST_cell_30975 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_17__Q), .b(FE_OFN219_n_9853), .o(TIMEBOOST_net_9592) );
na03f02 TIMEBOOST_cell_49899 ( .a(n_3910), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q), .c(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_15167) );
in01f02 g62435_u0 ( .a(n_6645), .o(g62435_sb) );
na03f02 TIMEBOOST_cell_73488 ( .a(TIMEBOOST_net_23334), .b(g61855_db), .c(TIMEBOOST_net_23348), .o(n_14825) );
na03f02 TIMEBOOST_cell_67037 ( .a(FE_OFN1602_n_13995), .b(TIMEBOOST_net_16539), .c(FE_OCPN2219_n_13997), .o(n_14439) );
na02f01 TIMEBOOST_cell_69352 ( .a(wbu_latency_tim_val_in_247), .b(n_6986), .o(TIMEBOOST_net_21884) );
in01m01 g62436_u0 ( .a(FE_OFN1241_n_4092), .o(g62436_sb) );
na03m02 TIMEBOOST_cell_66282 ( .a(g60635_sb), .b(TIMEBOOST_net_10050), .c(TIMEBOOST_net_5515), .o(n_5701) );
na03f02 TIMEBOOST_cell_73147 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q), .b(FE_OFN1076_n_4740), .c(TIMEBOOST_net_23298), .o(TIMEBOOST_net_17312) );
in01f02 g62437_u0 ( .a(FE_OFN1283_n_4097), .o(g62437_sb) );
na02m01 TIMEBOOST_cell_54089 ( .a(n_4479), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q), .o(TIMEBOOST_net_17262) );
na03f02 TIMEBOOST_cell_73235 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(g63538_sb), .c(g63538_db), .o(n_4617) );
in01m01 g62438_u0 ( .a(FE_OFN1241_n_4092), .o(g62438_sb) );
na04f04 TIMEBOOST_cell_24604 ( .a(n_9430), .b(g57561_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q), .d(FE_OFN1428_n_8567), .o(n_11191) );
na03f02 TIMEBOOST_cell_66736 ( .a(TIMEBOOST_net_16836), .b(FE_OFN1305_n_13124), .c(g54338_sb), .o(n_12980) );
in01f02 g62439_u0 ( .a(FE_OFN1310_n_6624), .o(g62439_sb) );
na03m04 TIMEBOOST_cell_63716 ( .a(n_4465), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q), .c(FE_OFN652_n_4508), .o(TIMEBOOST_net_20844) );
na02m01 TIMEBOOST_cell_26273 ( .a(wbu_addr_in_250), .b(FE_OFN1021_n_11877), .o(TIMEBOOST_net_7241) );
in01f02 g62440_u0 ( .a(FE_OFN1278_n_4097), .o(g62440_sb) );
na02f02 TIMEBOOST_cell_71576 ( .a(FE_OFN2209_n_11027), .b(TIMEBOOST_net_8605), .o(TIMEBOOST_net_22996) );
in01f02 g62441_u0 ( .a(FE_OFN2064_n_6391), .o(g62441_sb) );
na02m01 TIMEBOOST_cell_48117 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q), .b(FE_OFN665_n_4495), .o(TIMEBOOST_net_14276) );
in01f01 g62442_u0 ( .a(FE_OFN1261_n_4143), .o(g62442_sb) );
na02f01 TIMEBOOST_cell_48000 ( .a(TIMEBOOST_net_14217), .b(FE_OFN614_n_4501), .o(TIMEBOOST_net_12603) );
in01f02 TIMEBOOST_cell_17852 ( .a(TIMEBOOST_net_5263), .o(TIMEBOOST_net_5262) );
in01s01 TIMEBOOST_cell_73891 ( .a(TIMEBOOST_net_23455), .o(TIMEBOOST_net_23456) );
in01f01 g62443_u0 ( .a(FE_OFN1247_n_4093), .o(g62443_sb) );
na03f20 TIMEBOOST_cell_23950 ( .a(g75160_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .c(g75160_db), .o(n_16533) );
in01f04 g62444_u0 ( .a(FE_OFN1323_n_6436), .o(g62444_sb) );
na02s01 TIMEBOOST_cell_52723 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q), .o(TIMEBOOST_net_16579) );
na02f02 TIMEBOOST_cell_3756 ( .a(n_2904), .b(n_3034), .o(TIMEBOOST_net_438) );
in01f01 g62445_u0 ( .a(FE_OFN1212_n_4151), .o(g62445_sb) );
na02m02 TIMEBOOST_cell_71993 ( .a(TIMEBOOST_net_23204), .b(TIMEBOOST_net_16605), .o(TIMEBOOST_net_13232) );
in01f02 g62446_u0 ( .a(FE_OFN1311_n_6624), .o(g62446_sb) );
in01m01 TIMEBOOST_cell_31887 ( .a(conf_wb_err_addr_in_953), .o(TIMEBOOST_net_10051) );
na02f02 TIMEBOOST_cell_3757 ( .a(TIMEBOOST_net_438), .b(n_4119), .o(n_4856) );
na03f04 TIMEBOOST_cell_73165 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q), .b(g64288_sb), .c(g64288_db), .o(n_3885) );
in01f02 g62447_u0 ( .a(n_6431), .o(g62447_sb) );
na03m04 TIMEBOOST_cell_72540 ( .a(g64759_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q), .c(TIMEBOOST_net_14195), .o(TIMEBOOST_net_17070) );
na02s01 TIMEBOOST_cell_31011 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_4__Q), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_9610) );
in01f02 g62448_u0 ( .a(FE_OFN1215_n_4151), .o(g62448_sb) );
na02s01 TIMEBOOST_cell_47703 ( .a(n_2515), .b(g66417_db), .o(TIMEBOOST_net_14069) );
na02m01 TIMEBOOST_cell_69624 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q), .o(TIMEBOOST_net_22020) );
in01s01 TIMEBOOST_cell_73910 ( .a(n_2501), .o(TIMEBOOST_net_23475) );
in01f02 g62449_u0 ( .a(FE_OFN1293_n_4098), .o(g62449_sb) );
na03m02 TIMEBOOST_cell_65152 ( .a(TIMEBOOST_net_14388), .b(g65337_sb), .c(TIMEBOOST_net_17262), .o(TIMEBOOST_net_13240) );
na03f02 TIMEBOOST_cell_73668 ( .a(TIMEBOOST_net_13088), .b(FE_OFN1116_g64577_p), .c(g62772_sb), .o(n_5450) );
in01m01 g62450_u0 ( .a(FE_OFN1222_n_6391), .o(g62450_sb) );
na02f06 TIMEBOOST_cell_3279 ( .a(TIMEBOOST_net_199), .b(n_2694), .o(n_3147) );
na02f04 TIMEBOOST_cell_49368 ( .a(TIMEBOOST_net_14901), .b(g54311_db), .o(n_13018) );
na02f02 TIMEBOOST_cell_3280 ( .a(n_2427), .b(n_2431), .o(TIMEBOOST_net_200) );
in01f02 g62451_u0 ( .a(FE_OFN1317_n_6624), .o(g62451_sb) );
in01s01 TIMEBOOST_cell_67716 ( .a(TIMEBOOST_net_21142), .o(TIMEBOOST_net_21143) );
na02m01 TIMEBOOST_cell_44017 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(FE_OFN1042_n_2037), .o(TIMEBOOST_net_12903) );
in01f02 g62452_u0 ( .a(FE_OFN1285_n_4097), .o(g62452_sb) );
na03f02 TIMEBOOST_cell_68008 ( .a(TIMEBOOST_net_17445), .b(FE_OFN1293_n_4098), .c(g62949_sb), .o(n_5983) );
na02m10 TIMEBOOST_cell_52655 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q), .o(TIMEBOOST_net_16545) );
na03f02 TIMEBOOST_cell_66899 ( .a(FE_OFN1747_n_12004), .b(TIMEBOOST_net_15999), .c(n_11977), .o(n_12622) );
in01f02 g62453_u0 ( .a(FE_OFN1319_n_6436), .o(g62453_sb) );
in01s01 TIMEBOOST_cell_73858 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_), .o(TIMEBOOST_net_23423) );
in01m01 g62454_u0 ( .a(FE_OFN1208_n_6356), .o(g62454_sb) );
na02s01 TIMEBOOST_cell_70434 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q), .b(TIMEBOOST_net_16966), .o(TIMEBOOST_net_22425) );
in01f02 g62455_u0 ( .a(FE_OFN1232_n_6391), .o(g62455_sb) );
na02m02 TIMEBOOST_cell_50669 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q), .b(g58290_sb), .o(TIMEBOOST_net_15552) );
na02f01 TIMEBOOST_cell_3494 ( .a(FE_OFN2093_n_2301), .b(FE_OCPN1838_n_1238), .o(TIMEBOOST_net_307) );
in01m01 g62456_u0 ( .a(FE_OFN1193_n_6935), .o(g62456_sb) );
na04f02 TIMEBOOST_cell_72667 ( .a(TIMEBOOST_net_21519), .b(FE_OFN930_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q), .d(g64317_sb), .o(TIMEBOOST_net_13067) );
in01s01 TIMEBOOST_cell_73981 ( .a(TIMEBOOST_net_23545), .o(TIMEBOOST_net_23546) );
in01f02 g62457_u0 ( .a(FE_OFN2063_n_6391), .o(g62457_sb) );
na02f01 TIMEBOOST_cell_3495 ( .a(TIMEBOOST_net_307), .b(n_2725), .o(n_3363) );
na02f02 TIMEBOOST_cell_69841 ( .a(TIMEBOOST_net_22128), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_11039) );
in01f02 g62458_u0 ( .a(FE_OFN1212_n_4151), .o(g62458_sb) );
na02s02 TIMEBOOST_cell_52476 ( .a(TIMEBOOST_net_16455), .b(g57933_sb), .o(TIMEBOOST_net_9511) );
na02f02 TIMEBOOST_cell_71611 ( .a(TIMEBOOST_net_23013), .b(n_11823), .o(n_12515) );
na03f02 TIMEBOOST_cell_73512 ( .a(TIMEBOOST_net_13363), .b(n_6645), .c(g62924_sb), .o(n_6033) );
in01f02 g62459_u0 ( .a(FE_OFN1285_n_4097), .o(g62459_sb) );
na04f04 TIMEBOOST_cell_24798 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q), .b(g58804_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q), .d(FE_OFN2157_n_16439), .o(n_8637) );
na04f04 TIMEBOOST_cell_24800 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q), .b(g58802_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q), .d(FE_OFN2153_n_16439), .o(n_8640) );
in01f02 g62460_u0 ( .a(FE_OFN1225_n_6391), .o(g62460_sb) );
na04f04 TIMEBOOST_cell_24802 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q), .b(g58835_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q), .d(FE_OFN2153_n_16439), .o(n_8602) );
na02s01 TIMEBOOST_cell_51543 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q), .o(TIMEBOOST_net_15989) );
in01f02 g62461_u0 ( .a(FE_OFN1232_n_6391), .o(g62461_sb) );
na02f02 TIMEBOOST_cell_44139 ( .a(n_3982), .b(g62835_db), .o(TIMEBOOST_net_12964) );
na02f01 TIMEBOOST_cell_38013 ( .a(TIMEBOOST_net_10618), .b(g65312_sb), .o(n_3568) );
na02f01 TIMEBOOST_cell_45090 ( .a(TIMEBOOST_net_13439), .b(g63070_sb), .o(n_5110) );
in01f02 g62462_u0 ( .a(FE_OFN1204_n_4090), .o(g62462_sb) );
na03f02 TIMEBOOST_cell_66467 ( .a(TIMEBOOST_net_16789), .b(FE_OFN1311_n_6624), .c(g62345_sb), .o(n_6910) );
na02f01 TIMEBOOST_cell_3220 ( .a(n_15065), .b(wbu_map_in_131), .o(TIMEBOOST_net_170) );
na03f02 TIMEBOOST_cell_66077 ( .a(n_2057), .b(g63397_sb), .c(TIMEBOOST_net_7515), .o(n_4130) );
in01m02 g62463_u0 ( .a(FE_OFN1294_n_4098), .o(g62463_sb) );
na03f02 TIMEBOOST_cell_66468 ( .a(TIMEBOOST_net_17114), .b(FE_OFN1323_n_6436), .c(g62558_sb), .o(n_6446) );
in01f02 TIMEBOOST_cell_17848 ( .a(TIMEBOOST_net_5259), .o(TIMEBOOST_net_5258) );
na03m02 TIMEBOOST_cell_72473 ( .a(TIMEBOOST_net_16144), .b(FE_OFN904_n_4736), .c(g64120_sb), .o(TIMEBOOST_net_20468) );
in01f02 g62464_u0 ( .a(FE_OFN1213_n_4151), .o(g62464_sb) );
na03f02 TIMEBOOST_cell_34799 ( .a(TIMEBOOST_net_9549), .b(FE_OFN1403_n_8567), .c(g57097_sb), .o(n_10485) );
na03f02 TIMEBOOST_cell_73236 ( .a(n_2261), .b(g63196_sb), .c(TIMEBOOST_net_22883), .o(n_13505) );
na03f04 TIMEBOOST_cell_73237 ( .a(n_2710), .b(n_2301), .c(n_3027), .o(TIMEBOOST_net_15730) );
in01f02 g62465_u0 ( .a(FE_OFN1235_n_6391), .o(g62465_sb) );
in01s01 TIMEBOOST_cell_73845 ( .a(TIMEBOOST_net_23409), .o(TIMEBOOST_net_23410) );
na02s06 TIMEBOOST_cell_53047 ( .a(configuration_pci_err_data_508), .b(wbm_dat_o_7_), .o(TIMEBOOST_net_16741) );
na03f40 TIMEBOOST_cell_64293 ( .a(n_994), .b(n_1165), .c(n_1669), .o(n_2011) );
in01m02 g62466_u0 ( .a(FE_OFN1219_n_6886), .o(g62466_sb) );
na03m02 TIMEBOOST_cell_65371 ( .a(TIMEBOOST_net_20344), .b(g65014_sb), .c(n_4343), .o(TIMEBOOST_net_13243) );
na03f02 TIMEBOOST_cell_73820 ( .a(n_13891), .b(TIMEBOOST_net_16555), .c(FE_OFN1596_n_13741), .o(g53238_p) );
in01f02 g62467_u0 ( .a(FE_OFN1260_n_4143), .o(g62467_sb) );
na02s01 TIMEBOOST_cell_37233 ( .a(TIMEBOOST_net_10228), .b(g65853_sb), .o(n_1567) );
na02s01 TIMEBOOST_cell_45397 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q), .o(TIMEBOOST_net_13593) );
na02m02 TIMEBOOST_cell_49208 ( .a(TIMEBOOST_net_14821), .b(g58367_da), .o(n_9459) );
in01m01 g62468_u0 ( .a(FE_OFN1193_n_6935), .o(g62468_sb) );
na02f08 TIMEBOOST_cell_3281 ( .a(TIMEBOOST_net_200), .b(n_2437), .o(n_2432) );
na02f06 TIMEBOOST_cell_49367 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_787), .b(g54311_sb), .o(TIMEBOOST_net_14901) );
na02f01 TIMEBOOST_cell_44296 ( .a(TIMEBOOST_net_13042), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_11311) );
in01f02 g62469_u0 ( .a(FE_OFN2064_n_6391), .o(g62469_sb) );
na02m08 TIMEBOOST_cell_53009 ( .a(wbm_adr_o_5_), .b(configuration_pci_err_addr_475), .o(TIMEBOOST_net_16722) );
in01f02 g62470_u0 ( .a(FE_OFN1208_n_6356), .o(g62470_sb) );
na03f02 TIMEBOOST_cell_66726 ( .a(TIMEBOOST_net_17397), .b(FE_OFN1204_n_4090), .c(g62462_sb), .o(n_6672) );
na02s01 TIMEBOOST_cell_18172 ( .a(TIMEBOOST_net_5449), .b(g65893_sb), .o(n_2590) );
in01s01 TIMEBOOST_cell_17897 ( .a(TIMEBOOST_net_5308), .o(wbs_sel_i_0_) );
in01f01 g62471_u0 ( .a(FE_OFN1261_n_4143), .o(g62471_sb) );
na02s01 TIMEBOOST_cell_42865 ( .a(FE_OFN601_n_9687), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q), .o(TIMEBOOST_net_12327) );
na02s04 TIMEBOOST_cell_17921 ( .a(pci_target_unit_del_sync_comp_cycle_count_7_), .b(pci_target_unit_del_sync_comp_cycle_count_4_), .o(TIMEBOOST_net_5324) );
in01f02 g62472_u0 ( .a(n_6645), .o(g62472_sb) );
in01s01 TIMEBOOST_cell_31883 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .o(TIMEBOOST_net_10047) );
na02s02 TIMEBOOST_cell_47816 ( .a(TIMEBOOST_net_14125), .b(TIMEBOOST_net_10229), .o(TIMEBOOST_net_9561) );
in01f02 g62473_u0 ( .a(FE_OFN1234_n_6391), .o(g62473_sb) );
na02m01 TIMEBOOST_cell_68170 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_402), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q), .o(TIMEBOOST_net_21293) );
in01f01 g62474_u0 ( .a(FE_OFN1275_n_4096), .o(g62474_sb) );
na02f10 TIMEBOOST_cell_62882 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_785), .o(TIMEBOOST_net_20388) );
na02m02 TIMEBOOST_cell_44981 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_402), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_13385) );
na02m01 TIMEBOOST_cell_17918 ( .a(TIMEBOOST_net_5322), .b(n_9), .o(TIMEBOOST_net_275) );
in01f02 g62475_u0 ( .a(n_6319), .o(g62475_sb) );
in01s01 TIMEBOOST_cell_31884 ( .a(TIMEBOOST_net_10047), .o(TIMEBOOST_net_10048) );
na02f02 TIMEBOOST_cell_51376 ( .a(TIMEBOOST_net_15905), .b(n_4871), .o(n_4873) );
in01f02 g62476_u0 ( .a(FE_OFN1206_n_6356), .o(g62476_sb) );
na04s02 TIMEBOOST_cell_33454 ( .a(g57987_sb), .b(FE_OFN264_n_9849), .c(g57987_db), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q), .o(TIMEBOOST_net_9427) );
in01s01 TIMEBOOST_cell_17896 ( .a(TIMEBOOST_net_5306), .o(TIMEBOOST_net_5307) );
in01s01 TIMEBOOST_cell_17895 ( .a(parchk_pci_cbe_en_in), .o(TIMEBOOST_net_5306) );
in01f02 g62477_u0 ( .a(FE_OFN1311_n_6624), .o(g62477_sb) );
na03s02 TIMEBOOST_cell_41736 ( .a(g58340_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q), .c(g58340_db), .o(n_9480) );
na04f04 TIMEBOOST_cell_67668 ( .a(TIMEBOOST_net_15243), .b(FE_OFN1202_n_4090), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q), .d(g62587_sb), .o(n_6376) );
in01f02 g62478_u0 ( .a(n_6232), .o(g62478_sb) );
na04m04 TIMEBOOST_cell_67666 ( .a(TIMEBOOST_net_21026), .b(FE_OFN580_n_9531), .c(g58385_sb), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q), .o(TIMEBOOST_net_9512) );
in01f01 g62479_u0 ( .a(FE_OFN1222_n_6391), .o(g62479_sb) );
na03f02 TIMEBOOST_cell_34767 ( .a(TIMEBOOST_net_9362), .b(FE_OFN1377_n_8567), .c(g57164_sb), .o(n_10838) );
na03m02 TIMEBOOST_cell_73166 ( .a(g64266_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q), .c(TIMEBOOST_net_14744), .o(TIMEBOOST_net_8331) );
in01f02 g62480_u0 ( .a(FE_OFN1222_n_6391), .o(g62480_sb) );
na03f02 TIMEBOOST_cell_34802 ( .a(TIMEBOOST_net_9507), .b(FE_OFN1411_n_8567), .c(g57287_sb), .o(n_11466) );
na03m02 TIMEBOOST_cell_72791 ( .a(TIMEBOOST_net_23163), .b(g65029_sb), .c(TIMEBOOST_net_21853), .o(TIMEBOOST_net_17115) );
na02m02 TIMEBOOST_cell_68591 ( .a(TIMEBOOST_net_21503), .b(TIMEBOOST_net_14121), .o(TIMEBOOST_net_17384) );
in01f02 g62481_u0 ( .a(FE_OFN1317_n_6624), .o(g62481_sb) );
na03f02 TIMEBOOST_cell_73238 ( .a(n_3345), .b(g59383_sb), .c(TIMEBOOST_net_15802), .o(n_13511) );
in01f02 g62482_u0 ( .a(FE_OFN1288_n_4098), .o(g62482_sb) );
na02s02 TIMEBOOST_cell_17923 ( .a(pci_target_unit_del_sync_comp_cycle_count_14_), .b(pci_target_unit_del_sync_comp_cycle_count_13_), .o(TIMEBOOST_net_5325) );
na04m08 TIMEBOOST_cell_67514 ( .a(g57985_db), .b(FE_OFN262_n_9851), .c(g57985_sb), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q), .o(TIMEBOOST_net_17171) );
in01f02 g62483_u0 ( .a(FE_OFN1293_n_4098), .o(g62483_sb) );
na02f02 TIMEBOOST_cell_53872 ( .a(TIMEBOOST_net_17153), .b(FE_OFN1258_n_4143), .o(TIMEBOOST_net_15375) );
na03m02 TIMEBOOST_cell_64517 ( .a(n_3744), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q), .c(FE_OFN643_n_4677), .o(TIMEBOOST_net_10702) );
na02s01 TIMEBOOST_cell_45601 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q), .o(TIMEBOOST_net_13695) );
in01f02 g62484_u0 ( .a(FE_OFN1317_n_6624), .o(g62484_sb) );
na03f08 TIMEBOOST_cell_64304 ( .a(n_15014), .b(n_1432), .c(TIMEBOOST_net_5319), .o(n_5742) );
na03m02 TIMEBOOST_cell_72830 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q), .b(n_3785), .c(FE_OFN631_n_4454), .o(TIMEBOOST_net_16245) );
in01f01 g62485_u0 ( .a(FE_OFN1258_n_4143), .o(g62485_sb) );
na02f08 TIMEBOOST_cell_37221 ( .a(TIMEBOOST_net_10222), .b(n_3123), .o(FE_RN_273_0) );
na03s02 TIMEBOOST_cell_41738 ( .a(g58428_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q), .c(g58428_db), .o(n_9419) );
na03m06 TIMEBOOST_cell_70150 ( .a(FE_OFN1075_n_4740), .b(TIMEBOOST_net_16946), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q), .o(TIMEBOOST_net_22283) );
in01f02 g62486_u0 ( .a(FE_OFN1317_n_6624), .o(g62486_sb) );
na03f02 TIMEBOOST_cell_73624 ( .a(TIMEBOOST_net_16815), .b(n_16748), .c(g52653_sb), .o(n_14733) );
na02s02 TIMEBOOST_cell_48541 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q), .b(g65978_sb), .o(TIMEBOOST_net_14488) );
na03f02 TIMEBOOST_cell_68916 ( .a(g64826_sb), .b(n_4488), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q), .o(TIMEBOOST_net_21666) );
in01f02 g62487_u0 ( .a(FE_OFN1268_n_4095), .o(g62487_sb) );
in01f01 g62488_u0 ( .a(FE_OFN1294_n_4098), .o(g62488_sb) );
na04f04 TIMEBOOST_cell_73167 ( .a(n_1889), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q), .c(FE_OFN710_n_8232), .d(g61892_sb), .o(n_8044) );
na03m06 TIMEBOOST_cell_64516 ( .a(n_3780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q), .c(FE_OFN622_n_4409), .o(TIMEBOOST_net_14248) );
in01m01 g62489_u0 ( .a(FE_OFN1193_n_6935), .o(g62489_sb) );
na02m10 TIMEBOOST_cell_52983 ( .a(wishbone_slave_unit_pcim_sm_data_in_653), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q), .o(TIMEBOOST_net_16709) );
na02s01 TIMEBOOST_cell_47853 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q), .o(TIMEBOOST_net_14144) );
na03f02 TIMEBOOST_cell_71292 ( .a(n_4209), .b(FE_OFN1700_n_5751), .c(g52447_db), .o(TIMEBOOST_net_22854) );
in01f01 g62490_u0 ( .a(FE_OFN1248_n_4093), .o(g62490_sb) );
na03m04 TIMEBOOST_cell_72610 ( .a(TIMEBOOST_net_23151), .b(FE_OFN615_n_4501), .c(TIMEBOOST_net_21742), .o(TIMEBOOST_net_17525) );
na02s01 TIMEBOOST_cell_48085 ( .a(FE_OFN223_n_9844), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q), .o(TIMEBOOST_net_14260) );
na02f02 TIMEBOOST_cell_42932 ( .a(g65904_db), .b(TIMEBOOST_net_12360), .o(n_2177) );
in01f02 g62491_u0 ( .a(n_6232), .o(g62491_sb) );
in01s01 TIMEBOOST_cell_31885 ( .a(wbm_adr_o_9_), .o(TIMEBOOST_net_10049) );
na02m02 TIMEBOOST_cell_31379 ( .a(n_4444), .b(FE_OFN636_n_4669), .o(TIMEBOOST_net_9794) );
na04m08 TIMEBOOST_cell_67225 ( .a(g64937_sb), .b(FE_OFN659_n_4392), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q), .d(n_4498), .o(n_4383) );
in01f02 g62492_u0 ( .a(FE_OFN1241_n_4092), .o(g62492_sb) );
na03s01 TIMEBOOST_cell_64303 ( .a(TIMEBOOST_net_10137), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_384), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q), .o(TIMEBOOST_net_16807) );
in01f02 g62493_u0 ( .a(n_6554), .o(g62493_sb) );
na02f01 TIMEBOOST_cell_44140 ( .a(TIMEBOOST_net_12964), .b(g62835_sb), .o(n_5303) );
na02s01 TIMEBOOST_cell_54023 ( .a(FE_OFN205_n_9140), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q), .o(TIMEBOOST_net_17229) );
na02s03 TIMEBOOST_cell_48910 ( .a(TIMEBOOST_net_14672), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_12771) );
in01f01 g62494_u0 ( .a(FE_OFN1276_n_4096), .o(g62494_sb) );
na02m02 TIMEBOOST_cell_63013 ( .a(TIMEBOOST_net_20453), .b(g58128_db), .o(TIMEBOOST_net_9491) );
na03f02 TIMEBOOST_cell_65850 ( .a(TIMEBOOST_net_14887), .b(g64157_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q), .o(TIMEBOOST_net_20465) );
in01f02 g62495_u0 ( .a(n_6287), .o(g62495_sb) );
na02s01 TIMEBOOST_cell_42957 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q), .o(TIMEBOOST_net_12373) );
na02s01 TIMEBOOST_cell_53373 ( .a(pci_target_unit_fifos_pcir_data_in), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_16904) );
in01m01 g62496_u0 ( .a(FE_OFN1249_n_4093), .o(g62496_sb) );
na03s02 TIMEBOOST_cell_70864 ( .a(FE_OFN252_n_9868), .b(FE_OFN589_n_9692), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_22640) );
na03f02 TIMEBOOST_cell_47429 ( .a(FE_OCP_RBN1996_n_13971), .b(TIMEBOOST_net_13743), .c(FE_OFN1586_n_13736), .o(g53222_p) );
na04m06 TIMEBOOST_cell_72749 ( .a(g64853_sb), .b(n_4479), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q), .d(TIMEBOOST_net_14331), .o(TIMEBOOST_net_13242) );
in01f02 g62497_u0 ( .a(FE_OFN1249_n_4093), .o(g62497_sb) );
na02s01 TIMEBOOST_cell_44202 ( .a(TIMEBOOST_net_12995), .b(FE_OFN268_n_9880), .o(n_9901) );
na04f02 TIMEBOOST_cell_73125 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q), .b(FE_OFN1075_n_4740), .c(pci_target_unit_fifos_pciw_addr_data_in_149), .d(g64209_sb), .o(n_3960) );
in01f04 g62498_u0 ( .a(FE_OFN1313_n_6624), .o(g62498_sb) );
na02s02 TIMEBOOST_cell_30647 ( .a(n_9573), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q), .o(TIMEBOOST_net_9428) );
na04f04 TIMEBOOST_cell_67697 ( .a(TIMEBOOST_net_16864), .b(FE_OFN2198_n_10256), .c(g52609_sb), .d(TIMEBOOST_net_700), .o(n_11862) );
na03s02 TIMEBOOST_cell_21320 ( .a(g58165_sb), .b(FE_OFN245_n_9114), .c(g58165_db), .o(n_9064) );
in01f01 g62499_u0 ( .a(FE_OFN1253_n_4143), .o(g62499_sb) );
na02m02 TIMEBOOST_cell_69434 ( .a(g64886_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q), .o(TIMEBOOST_net_21925) );
na02f02 TIMEBOOST_cell_41232 ( .a(FE_OFN1770_n_14054), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_12228) );
in01m01 g62500_u0 ( .a(FE_OFN1274_n_4096), .o(g62500_sb) );
na03f20 TIMEBOOST_cell_64317 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q), .b(n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_406), .o(TIMEBOOST_net_14856) );
na04f04 TIMEBOOST_cell_67699 ( .a(TIMEBOOST_net_16863), .b(FE_OFN2200_n_10256), .c(g52599_sb), .d(TIMEBOOST_net_707), .o(n_11873) );
in01f02 g62501_u0 ( .a(FE_OFN1310_n_6624), .o(g62501_sb) );
na02s02 TIMEBOOST_cell_62786 ( .a(g61870_sb), .b(g62008_db), .o(TIMEBOOST_net_20340) );
na04f04 TIMEBOOST_cell_25005 ( .a(n_9312), .b(n_10173), .c(n_10176), .d(n_9311), .o(n_12160) );
in01m01 g62502_u0 ( .a(FE_OFN1295_n_4098), .o(g62502_sb) );
in01s01 TIMEBOOST_cell_45927 ( .a(TIMEBOOST_net_13888), .o(n_1064) );
na04f04 TIMEBOOST_cell_24670 ( .a(n_9524), .b(g57415_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q), .d(FE_OFN2185_n_8567), .o(n_11327) );
na04f04 TIMEBOOST_cell_24672 ( .a(n_9218), .b(g57406_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q), .d(FE_OFN2175_n_8567), .o(n_10828) );
in01f04 g62503_u0 ( .a(FE_OFN1250_n_4093), .o(g62503_sb) );
na02f01 TIMEBOOST_cell_29406 ( .a(TIMEBOOST_net_8807), .b(FE_OFN881_g64577_p), .o(TIMEBOOST_net_7413) );
na04f04 TIMEBOOST_cell_24674 ( .a(n_9539), .b(g57402_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q), .d(FE_OFN2173_n_8567), .o(n_11340) );
in01f02 g62504_u0 ( .a(FE_OFN1322_n_6436), .o(g62504_sb) );
na04f04 TIMEBOOST_cell_73314 ( .a(n_4056), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q), .c(FE_OFN1119_g64577_p), .d(g62743_sb), .o(n_5493) );
na02f04 TIMEBOOST_cell_68412 ( .a(n_13447), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q), .o(TIMEBOOST_net_21414) );
na03f02 TIMEBOOST_cell_73446 ( .a(TIMEBOOST_net_20949), .b(FE_OFN1200_n_4090), .c(g62999_sb), .o(n_5884) );
in01f01 g62505_u0 ( .a(FE_OFN1268_n_4095), .o(g62505_sb) );
na02f04 TIMEBOOST_cell_40621 ( .a(TIMEBOOST_net_11922), .b(FE_RN_368_0), .o(FE_RN_369_0) );
na03m02 TIMEBOOST_cell_64515 ( .a(n_3749), .b(FE_OFN1628_n_4438), .c(n_27), .o(TIMEBOOST_net_14714) );
na04f04 TIMEBOOST_cell_24676 ( .a(n_9556), .b(g57379_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q), .d(FE_OFN2185_n_8567), .o(n_11369) );
in01m02 g62506_u0 ( .a(FE_OFN369_n_4092), .o(g62506_sb) );
na02m02 TIMEBOOST_cell_45134 ( .a(TIMEBOOST_net_13461), .b(g62592_sb), .o(n_6369) );
no03f08 TIMEBOOST_cell_24678 ( .a(TIMEBOOST_net_688), .b(n_8819), .c(FE_RN_280_0), .o(n_15611) );
na02s02 TIMEBOOST_cell_49283 ( .a(g58443_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q), .o(TIMEBOOST_net_14859) );
in01f02 g62507_u0 ( .a(FE_OFN1223_n_6391), .o(g62507_sb) );
in01s01 TIMEBOOST_cell_45928 ( .a(TIMEBOOST_net_13889), .o(TIMEBOOST_net_13888) );
na02f02 TIMEBOOST_cell_69353 ( .a(TIMEBOOST_net_21884), .b(g60672_sb), .o(TIMEBOOST_net_5482) );
na03f02 TIMEBOOST_cell_34753 ( .a(TIMEBOOST_net_9405), .b(FE_OFN1390_n_8567), .c(g57459_sb), .o(n_11274) );
in01f02 g62508_u0 ( .a(FE_OFN1243_n_4092), .o(g62508_sb) );
na03m02 TIMEBOOST_cell_72768 ( .a(n_4482), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q), .c(TIMEBOOST_net_12687), .o(TIMEBOOST_net_20542) );
na02s02 TIMEBOOST_cell_44019 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q), .b(FE_OFN539_n_9690), .o(TIMEBOOST_net_12904) );
in01f01 g62509_u0 ( .a(FE_OFN1243_n_4092), .o(g62509_sb) );
in01m01 TIMEBOOST_cell_45885 ( .a(parchk_pci_ad_out_in_1192), .o(TIMEBOOST_net_13846) );
na02m02 TIMEBOOST_cell_68768 ( .a(g64856_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q), .o(TIMEBOOST_net_21592) );
na03f02 TIMEBOOST_cell_34903 ( .a(TIMEBOOST_net_9448), .b(FE_OFN1400_n_8567), .c(g57460_sb), .o(n_10344) );
in01f02 g62510_u0 ( .a(FE_OFN1270_n_4095), .o(g62510_sb) );
na02m02 TIMEBOOST_cell_48802 ( .a(TIMEBOOST_net_14618), .b(TIMEBOOST_net_11079), .o(TIMEBOOST_net_9553) );
na02s01 TIMEBOOST_cell_17917 ( .a(n_692), .b(wishbone_slave_unit_pci_initiator_if_read_count_3_), .o(TIMEBOOST_net_5322) );
na02f08 TIMEBOOST_cell_17916 ( .a(n_2235), .b(TIMEBOOST_net_5321), .o(TIMEBOOST_net_87) );
in01f02 g62511_u0 ( .a(n_6554), .o(g62511_sb) );
na02f01 TIMEBOOST_cell_43506 ( .a(TIMEBOOST_net_12647), .b(g65215_sb), .o(n_2653) );
na03f02 TIMEBOOST_cell_69674 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q), .b(TIMEBOOST_net_14283), .c(g65854_db), .o(TIMEBOOST_net_22045) );
in01f02 g62512_u0 ( .a(FE_OFN1222_n_6391), .o(g62512_sb) );
na03f10 TIMEBOOST_cell_35130 ( .a(g75416_db), .b(FE_OCP_RBN1956_n_16981), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_16970) );
na02m10 TIMEBOOST_cell_45767 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q), .o(TIMEBOOST_net_13778) );
na03f10 TIMEBOOST_cell_36069 ( .a(n_16163), .b(n_3422), .c(n_5722), .o(n_8452) );
in01f02 g62513_u0 ( .a(FE_OFN1222_n_6391), .o(g62513_sb) );
in01s01 TIMEBOOST_cell_45879 ( .a(TIMEBOOST_net_13943), .o(TIMEBOOST_net_13840) );
na02f01 TIMEBOOST_cell_3292 ( .a(n_15762), .b(FE_OFN197_n_2683), .o(TIMEBOOST_net_206) );
in01f02 g62514_u0 ( .a(FE_OFN1244_n_4092), .o(g62514_sb) );
na04f04 TIMEBOOST_cell_67701 ( .a(TIMEBOOST_net_16861), .b(FE_OFN2200_n_10256), .c(g52601_sb), .d(TIMEBOOST_net_710), .o(n_11870) );
na02m02 TIMEBOOST_cell_17915 ( .a(n_1412), .b(n_1674), .o(TIMEBOOST_net_5321) );
na02s02 TIMEBOOST_cell_17914 ( .a(TIMEBOOST_net_5320), .b(n_523), .o(TIMEBOOST_net_168) );
in01f01 g62515_u0 ( .a(FE_OFN1226_n_6391), .o(g62515_sb) );
in01s01 TIMEBOOST_cell_67722 ( .a(TIMEBOOST_net_21148), .o(TIMEBOOST_net_21149) );
in01f03 TIMEBOOST_cell_17846 ( .a(TIMEBOOST_net_5257), .o(TIMEBOOST_net_5256) );
na02s01 TIMEBOOST_cell_17913 ( .a(pci_target_unit_del_sync_comp_cycle_count_10_), .b(pci_target_unit_del_sync_comp_cycle_count_11_), .o(TIMEBOOST_net_5320) );
in01m01 g62516_u0 ( .a(FE_OFN1222_n_6391), .o(g62516_sb) );
na02f01 TIMEBOOST_cell_3293 ( .a(TIMEBOOST_net_206), .b(n_3386), .o(n_4533) );
na02f02 g62516_u2 ( .a(n_3650), .b(FE_OFN1222_n_6391), .o(g62516_db) );
na03f02 TIMEBOOST_cell_67039 ( .a(FE_OFN1606_n_13997), .b(TIMEBOOST_net_16532), .c(FE_OFN1600_n_13995), .o(n_14459) );
in01f02 g62517_u0 ( .a(FE_OFN1224_n_6391), .o(g62517_sb) );
na02m02 TIMEBOOST_cell_68751 ( .a(TIMEBOOST_net_21583), .b(TIMEBOOST_net_10445), .o(TIMEBOOST_net_20587) );
na04m04 TIMEBOOST_cell_67902 ( .a(n_3785), .b(g64950_sb), .c(g64950_db), .d(n_3665), .o(TIMEBOOST_net_17578) );
na02s01 TIMEBOOST_cell_48721 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q), .b(FE_OFN585_n_9692), .o(TIMEBOOST_net_14578) );
in01f02 g62518_u0 ( .a(FE_OFN1314_n_6624), .o(g62518_sb) );
na02m10 TIMEBOOST_cell_53433 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_146), .o(TIMEBOOST_net_16934) );
na02f02 TIMEBOOST_cell_3777 ( .a(TIMEBOOST_net_448), .b(n_7033), .o(n_7504) );
na02m02 TIMEBOOST_cell_54060 ( .a(TIMEBOOST_net_17247), .b(FE_OFN1049_n_16657), .o(TIMEBOOST_net_14717) );
in01f02 g62519_u0 ( .a(FE_OFN1317_n_6624), .o(g62519_sb) );
na02m02 TIMEBOOST_cell_49660 ( .a(TIMEBOOST_net_15047), .b(g61716_sb), .o(n_8393) );
na02f04 TIMEBOOST_cell_3779 ( .a(TIMEBOOST_net_449), .b(n_16970), .o(n_13703) );
in01f02 g62520_u0 ( .a(FE_OFN1316_n_6624), .o(g62520_sb) );
in01s01 TIMEBOOST_cell_67732 ( .a(TIMEBOOST_net_21158), .o(TIMEBOOST_net_21159) );
na04m06 TIMEBOOST_cell_65886 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q), .b(g58009_sb), .c(FE_OFN258_n_9862), .d(g58009_db), .o(TIMEBOOST_net_16845) );
in01f02 g62521_u0 ( .a(FE_OFN1260_n_4143), .o(g62521_sb) );
in01f06 TIMEBOOST_cell_17847 ( .a(TIMEBOOST_net_5258), .o(n_8540) );
na03f02 TIMEBOOST_cell_73821 ( .a(n_13891), .b(TIMEBOOST_net_16556), .c(FE_OCP_RBN1961_FE_OFN1591_n_13741), .o(g53226_p) );
in01f02 g62522_u0 ( .a(FE_OFN1260_n_4143), .o(g62522_sb) );
na02m02 TIMEBOOST_cell_68964 ( .a(g64800_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q), .o(TIMEBOOST_net_21690) );
na02m08 TIMEBOOST_cell_17911 ( .a(n_288), .b(wbu_wb_init_complete_in), .o(TIMEBOOST_net_5319) );
in01f10 TIMEBOOST_cell_17845 ( .a(TIMEBOOST_net_5256), .o(FE_OFN1000_n_15978) );
in01f02 g62523_u0 ( .a(FE_OFN1314_n_6624), .o(g62523_sb) );
na02f02 TIMEBOOST_cell_3783 ( .a(TIMEBOOST_net_451), .b(FE_RN_438_0), .o(FE_RN_439_0) );
na04f04 TIMEBOOST_cell_24176 ( .a(n_9216), .b(g57434_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q), .d(FE_OFN1416_n_8567), .o(n_10821) );
in01m01 g62524_u0 ( .a(FE_OFN1249_n_4093), .o(g62524_sb) );
in01m20 TIMEBOOST_cell_17844 ( .a(TIMEBOOST_net_5255), .o(TIMEBOOST_net_5254) );
in01s01 TIMEBOOST_cell_17879 ( .a(TIMEBOOST_net_5290), .o(wbs_dat_i_12_) );
in01f01 g62525_u0 ( .a(FE_OFN1248_n_4093), .o(g62525_sb) );
na03f04 TIMEBOOST_cell_71824 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .c(g65270_sb), .o(TIMEBOOST_net_23120) );
in01s01 TIMEBOOST_cell_17878 ( .a(TIMEBOOST_net_5289), .o(TIMEBOOST_net_5288) );
in01s01 TIMEBOOST_cell_45978 ( .a(TIMEBOOST_net_13938), .o(TIMEBOOST_net_13939) );
in01f02 g62526_u0 ( .a(FE_OFN1278_n_4097), .o(g62526_sb) );
in01s01 TIMEBOOST_cell_17900 ( .a(TIMEBOOST_net_5311), .o(TIMEBOOST_net_5310) );
in01f02 g62527_u0 ( .a(FE_OFN1282_n_4097), .o(g62527_sb) );
na02s02 TIMEBOOST_cell_70722 ( .a(FE_OFN201_n_9230), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q), .o(TIMEBOOST_net_22569) );
na04f04 TIMEBOOST_cell_24692 ( .a(wishbone_slave_unit_fifos_wbr_be_in_266), .b(g58841_sb), .c(TIMEBOOST_net_13903), .d(FE_OFN1438_n_9372), .o(n_8673) );
in01m01 g62528_u0 ( .a(FE_OFN1219_n_6886), .o(g62528_sb) );
na02m02 TIMEBOOST_cell_68166 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q), .b(FE_OFN2055_n_8831), .o(TIMEBOOST_net_21291) );
na02f02 TIMEBOOST_cell_39919 ( .a(TIMEBOOST_net_11571), .b(g62468_sb), .o(n_6657) );
in01f02 g62529_u0 ( .a(FE_OFN1231_n_6391), .o(g62529_sb) );
na02f02 TIMEBOOST_cell_70549 ( .a(TIMEBOOST_net_22482), .b(g59380_sb), .o(n_7679) );
in01f01 g62530_u0 ( .a(FE_OFN1250_n_4093), .o(g62530_sb) );
na03f02 TIMEBOOST_cell_68376 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q), .b(TIMEBOOST_net_12328), .c(FE_OFN906_n_4736), .o(TIMEBOOST_net_21396) );
na04f04 TIMEBOOST_cell_24694 ( .a(wishbone_slave_unit_fifos_wbr_be_in_264), .b(g58839_sb), .c(TIMEBOOST_net_13905), .d(FE_OFN1438_n_9372), .o(n_8675) );
na04f04 TIMEBOOST_cell_24626 ( .a(n_9831), .b(g57093_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q), .d(FE_OFN2169_n_8567), .o(n_11648) );
in01f02 g62531_u0 ( .a(FE_OFN1249_n_4093), .o(g62531_sb) );
na03m02 TIMEBOOST_cell_64514 ( .a(n_3749), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q), .c(FE_OFN672_n_4505), .o(TIMEBOOST_net_10335) );
na04f04 TIMEBOOST_cell_24696 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_1__Q), .b(g58837_sb), .c(n_1721), .d(FE_OFN1437_n_9372), .o(n_8677) );
in01f02 g62532_u0 ( .a(FE_OFN1233_n_6391), .o(g62532_sb) );
na03f02 TIMEBOOST_cell_34804 ( .a(TIMEBOOST_net_9553), .b(FE_OFN1409_n_8567), .c(g57417_sb), .o(n_11324) );
na02s01 TIMEBOOST_cell_68214 ( .a(pci_target_unit_del_sync_bc_in), .b(FE_OFN2094_n_2520), .o(TIMEBOOST_net_21315) );
in01f02 g62533_u0 ( .a(FE_OFN1230_n_6391), .o(g62533_sb) );
na02m02 TIMEBOOST_cell_44806 ( .a(TIMEBOOST_net_13297), .b(g60654_sb), .o(n_5669) );
na02f01 TIMEBOOST_cell_3510 ( .a(n_2313), .b(n_2314), .o(TIMEBOOST_net_315) );
in01f02 g62534_u0 ( .a(FE_OFN2064_n_6391), .o(g62534_sb) );
in01m01 TIMEBOOST_cell_31886 ( .a(TIMEBOOST_net_10049), .o(TIMEBOOST_net_10050) );
na02m08 TIMEBOOST_cell_51933 ( .a(pci_target_unit_del_sync_bc_in_202), .b(pci_target_unit_pcit_if_strd_bc_in_718), .o(TIMEBOOST_net_16184) );
na02m06 TIMEBOOST_cell_3512 ( .a(n_2756), .b(n_1229), .o(TIMEBOOST_net_316) );
in01f02 g62535_u0 ( .a(FE_OFN1315_n_6624), .o(g62535_sb) );
na02f02 TIMEBOOST_cell_3785 ( .a(TIMEBOOST_net_452), .b(n_5717), .o(n_7312) );
na02f02 TIMEBOOST_cell_3786 ( .a(n_2839), .b(n_2969), .o(TIMEBOOST_net_453) );
in01f04 g62536_u0 ( .a(FE_OFN1261_n_4143), .o(g62536_sb) );
na04f04 TIMEBOOST_cell_73239 ( .a(TIMEBOOST_net_7208), .b(FE_OFN1143_n_15261), .c(g62033_sb), .d(n_2744), .o(g53935_da) );
na04f04 TIMEBOOST_cell_24606 ( .a(n_9203), .b(g57558_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q), .d(FE_OFN2182_n_8567), .o(n_10803) );
in01f02 g62537_u0 ( .a(FE_OFN1258_n_4143), .o(g62537_sb) );
na02m10 TIMEBOOST_cell_45769 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q), .o(TIMEBOOST_net_13779) );
na04f04 TIMEBOOST_cell_24698 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_8__Q), .b(g58485_sb), .c(FE_OFN252_n_9868), .d(FE_OFN1437_n_9372), .o(n_9350) );
na02m01 TIMEBOOST_cell_63924 ( .a(configuration_pci_err_addr_497), .b(wbm_adr_o_27_), .o(TIMEBOOST_net_20948) );
in01m01 g62538_u0 ( .a(FE_OFN1283_n_4097), .o(g62538_sb) );
na03m02 TIMEBOOST_cell_69962 ( .a(TIMEBOOST_net_20362), .b(FE_OFN1036_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q), .o(TIMEBOOST_net_22189) );
na02s02 TIMEBOOST_cell_38594 ( .a(g58045_sb), .b(FE_OFN215_n_9856), .o(TIMEBOOST_net_10909) );
na03f02 TIMEBOOST_cell_66720 ( .a(TIMEBOOST_net_17374), .b(FE_OFN1268_n_4095), .c(g62678_sb), .o(n_6184) );
in01f01 g62539_u0 ( .a(FE_OFN1284_n_4097), .o(g62539_sb) );
na02m01 TIMEBOOST_cell_30531 ( .a(n_1609), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(TIMEBOOST_net_9370) );
na02f01 TIMEBOOST_cell_37558 ( .a(n_3739), .b(g64819_sb), .o(TIMEBOOST_net_10391) );
in01f02 g62540_u0 ( .a(n_6645), .o(g62540_sb) );
na02s03 TIMEBOOST_cell_68418 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q), .b(TIMEBOOST_net_13879), .o(TIMEBOOST_net_21417) );
in01m02 g62541_u0 ( .a(FE_OFN1219_n_6886), .o(g62541_sb) );
na03f02 TIMEBOOST_cell_72873 ( .a(TIMEBOOST_net_21748), .b(g64143_sb), .c(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_22479) );
na02f02 TIMEBOOST_cell_37559 ( .a(TIMEBOOST_net_10391), .b(g64819_db), .o(n_3740) );
in01s01 TIMEBOOST_cell_17899 ( .a(TIMEBOOST_net_5310), .o(wbs_sel_i_1_) );
in01m01 g62542_u0 ( .a(FE_OFN1242_n_4092), .o(g62542_sb) );
na03s02 TIMEBOOST_cell_33175 ( .a(n_1924), .b(g61777_sb), .c(g61777_db), .o(n_8253) );
in01f01 g62543_u0 ( .a(FE_OFN1284_n_4097), .o(g62543_sb) );
na03f02 TIMEBOOST_cell_34813 ( .a(TIMEBOOST_net_9531), .b(FE_OFN1404_n_8567), .c(g57297_sb), .o(n_11454) );
in01s01 TIMEBOOST_cell_17894 ( .a(TIMEBOOST_net_5305), .o(TIMEBOOST_net_5304) );
na02s01 TIMEBOOST_cell_39741 ( .a(TIMEBOOST_net_11482), .b(g57897_db), .o(n_9227) );
in01f01 g62544_u0 ( .a(FE_OFN1274_n_4096), .o(g62544_sb) );
in01s01 TIMEBOOST_cell_17898 ( .a(TIMEBOOST_net_5309), .o(TIMEBOOST_net_5308) );
in01s01 TIMEBOOST_cell_17888 ( .a(TIMEBOOST_net_5299), .o(TIMEBOOST_net_5298) );
in01m01 g62545_u0 ( .a(FE_OFN1274_n_4096), .o(g62545_sb) );
na02s01 TIMEBOOST_cell_48603 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q), .b(FE_OFN525_n_9899), .o(TIMEBOOST_net_14519) );
in01s01 TIMEBOOST_cell_17893 ( .a(TIMEBOOST_net_5304), .o(wbs_dat_i_6_) );
in01m01 g62546_u0 ( .a(FE_OFN1244_n_4092), .o(g62546_sb) );
na03f02 TIMEBOOST_cell_72551 ( .a(TIMEBOOST_net_23149), .b(FE_OFN916_n_4725), .c(g64335_sb), .o(TIMEBOOST_net_13042) );
na02f02 TIMEBOOST_cell_72213 ( .a(TIMEBOOST_net_23314), .b(g54149_sb), .o(n_13560) );
in01f02 g62547_u0 ( .a(FE_OFN1312_n_6624), .o(g62547_sb) );
na02f02 TIMEBOOST_cell_3787 ( .a(TIMEBOOST_net_453), .b(n_4125), .o(n_4855) );
na02m02 TIMEBOOST_cell_68816 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q), .b(FE_OFN639_n_4669), .o(TIMEBOOST_net_21616) );
in01f02 g62548_u0 ( .a(FE_OFN1243_n_4092), .o(g62548_sb) );
na03f02 TIMEBOOST_cell_72627 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q), .b(g65047_sb), .c(TIMEBOOST_net_10390), .o(TIMEBOOST_net_17083) );
in01s01 TIMEBOOST_cell_17892 ( .a(TIMEBOOST_net_5303), .o(TIMEBOOST_net_5302) );
in01s01 TIMEBOOST_cell_17891 ( .a(TIMEBOOST_net_5302), .o(wbs_dat_i_25_) );
in01m01 g62549_u0 ( .a(FE_OFN1244_n_4092), .o(g62549_sb) );
na03f02 TIMEBOOST_cell_68000 ( .a(TIMEBOOST_net_20954), .b(FE_OFN1212_n_4151), .c(g63190_sb), .o(n_5774) );
in01s01 TIMEBOOST_cell_17885 ( .a(TIMEBOOST_net_5296), .o(wbs_dat_i_24_) );
na02f02 TIMEBOOST_cell_52414 ( .a(TIMEBOOST_net_16424), .b(g63432_sb), .o(n_4627) );
in01f02 g62550_u0 ( .a(FE_OFN2063_n_6391), .o(g62550_sb) );
na04f02 TIMEBOOST_cell_73056 ( .a(n_1955), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q), .c(FE_OFN2081_n_8176), .d(g61786_sb), .o(n_8231) );
na02f08 TIMEBOOST_cell_3513 ( .a(n_2761), .b(TIMEBOOST_net_316), .o(n_3197) );
na03m02 TIMEBOOST_cell_73240 ( .a(TIMEBOOST_net_22160), .b(TIMEBOOST_net_14893), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q), .o(TIMEBOOST_net_13075) );
in01f02 g62551_u0 ( .a(FE_OFN1224_n_6391), .o(g62551_sb) );
na04f06 TIMEBOOST_cell_20898 ( .a(n_1365), .b(n_1350), .c(n_1433), .d(n_1352), .o(n_2400) );
na03s02 TIMEBOOST_cell_33176 ( .a(n_1948), .b(g61772_sb), .c(g61772_db), .o(n_8264) );
in01f02 g62552_u0 ( .a(FE_OFN1224_n_6391), .o(g62552_sb) );
na03f02 TIMEBOOST_cell_66752 ( .a(TIMEBOOST_net_16831), .b(FE_OFN1305_n_13124), .c(g54367_sb), .o(n_13123) );
na02f02 TIMEBOOST_cell_44207 ( .a(TIMEBOOST_net_7359), .b(n_2102), .o(TIMEBOOST_net_12998) );
na02f06 TIMEBOOST_cell_3302 ( .a(n_16474), .b(n_7114), .o(TIMEBOOST_net_211) );
in01f02 g62553_u0 ( .a(FE_OFN1232_n_6391), .o(g62553_sb) );
na02f06 TIMEBOOST_cell_3515 ( .a(TIMEBOOST_net_317), .b(n_2931), .o(n_3324) );
na02m08 TIMEBOOST_cell_45317 ( .a(n_395), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q), .o(TIMEBOOST_net_13553) );
in01f01 g62554_u0 ( .a(FE_OFN1268_n_4095), .o(g62554_sb) );
na02m01 TIMEBOOST_cell_62670 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q), .b(FE_OFN687_n_4417), .o(TIMEBOOST_net_20282) );
na04f04 TIMEBOOST_cell_24178 ( .a(n_9510), .b(g57432_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q), .d(FE_OFN1417_n_8567), .o(n_11302) );
in01m01 g62555_u0 ( .a(FE_OFN1270_n_4095), .o(g62555_sb) );
na02s01 TIMEBOOST_cell_54001 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q), .o(TIMEBOOST_net_17218) );
in01s01 TIMEBOOST_cell_17884 ( .a(TIMEBOOST_net_5295), .o(TIMEBOOST_net_5294) );
in01s01 TIMEBOOST_cell_17883 ( .a(TIMEBOOST_net_5294), .o(wbs_dat_i_3_) );
in01f01 g62556_u0 ( .a(FE_OFN1248_n_4093), .o(g62556_sb) );
na03f04 TIMEBOOST_cell_67002 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_16527), .c(FE_OFN1587_n_13736), .o(g53154_p) );
in01s01 TIMEBOOST_cell_17882 ( .a(TIMEBOOST_net_5293), .o(TIMEBOOST_net_5292) );
in01s01 TIMEBOOST_cell_17881 ( .a(TIMEBOOST_net_5292), .o(wbs_dat_i_7_) );
in01f02 g62557_u0 ( .a(FE_OFN1274_n_4096), .o(g62557_sb) );
na03m02 TIMEBOOST_cell_72246 ( .a(TIMEBOOST_net_20930), .b(FE_OFN1688_n_9528), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q), .o(TIMEBOOST_net_23331) );
in01s01 TIMEBOOST_cell_17890 ( .a(TIMEBOOST_net_5301), .o(TIMEBOOST_net_5300) );
in01s01 TIMEBOOST_cell_17877 ( .a(TIMEBOOST_net_5288), .o(wbs_dat_i_21_) );
in01f02 g62558_u0 ( .a(FE_OFN1323_n_6436), .o(g62558_sb) );
na02f02 TIMEBOOST_cell_3789 ( .a(TIMEBOOST_net_454), .b(n_6983), .o(n_7325) );
na02f04 TIMEBOOST_cell_3790 ( .a(FE_OCP_RBN2018_n_16970), .b(n_16974), .o(TIMEBOOST_net_455) );
in01f02 g62559_u0 ( .a(FE_OFN1212_n_4151), .o(g62559_sb) );
na03f02 TIMEBOOST_cell_34866 ( .a(TIMEBOOST_net_9347), .b(FE_OFN1407_n_8567), .c(g57494_sb), .o(n_10331) );
na03f02 TIMEBOOST_cell_34806 ( .a(TIMEBOOST_net_9441), .b(FE_OFN1401_n_8567), .c(g57334_sb), .o(n_10396) );
in01f02 g62560_u0 ( .a(FE_OFN1323_n_6436), .o(g62560_sb) );
na02m01 TIMEBOOST_cell_53968 ( .a(TIMEBOOST_net_17201), .b(n_4669), .o(TIMEBOOST_net_14117) );
na02f08 TIMEBOOST_cell_3791 ( .a(TIMEBOOST_net_455), .b(n_16967), .o(n_13743) );
na04f04 TIMEBOOST_cell_24813 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q), .b(g58824_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q), .d(FE_OFN2158_n_16439), .o(n_8617) );
in01f02 g62561_u0 ( .a(FE_OFN1323_n_6436), .o(g62561_sb) );
na03f04 TIMEBOOST_cell_73686 ( .a(TIMEBOOST_net_8004), .b(n_3037), .c(n_4641), .o(n_5728) );
na04f04 TIMEBOOST_cell_24804 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q), .b(g58833_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q), .d(FE_OFN2157_n_16439), .o(n_8604) );
na04f04 TIMEBOOST_cell_24805 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__Q), .b(g58832_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q), .d(FE_OFN2153_n_16439), .o(n_8605) );
in01f02 g62562_u0 ( .a(FE_OFN1313_n_6624), .o(g62562_sb) );
na04f04 TIMEBOOST_cell_24806 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q), .b(g58831_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q), .d(FE_OFN2156_n_16439), .o(n_8606) );
na04f04 TIMEBOOST_cell_24807 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q), .b(g58830_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q), .d(FE_OFN2157_n_16439), .o(n_8607) );
in01f02 g62563_u0 ( .a(n_6431), .o(g62563_sb) );
na02f01 TIMEBOOST_cell_49245 ( .a(pci_target_unit_fifos_pcir_data_in_163), .b(FE_OFN1042_n_2037), .o(TIMEBOOST_net_14840) );
in01m01 g62564_u0 ( .a(FE_OFN1193_n_6935), .o(g62564_sb) );
na02s02 TIMEBOOST_cell_49263 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q), .b(FE_OFN588_n_9692), .o(TIMEBOOST_net_14849) );
in01s01 TIMEBOOST_cell_17876 ( .a(TIMEBOOST_net_5287), .o(TIMEBOOST_net_5286) );
in01s01 TIMEBOOST_cell_17887 ( .a(TIMEBOOST_net_5298), .o(wbs_dat_i_4_) );
in01m01 g62565_u0 ( .a(FE_OFN1193_n_6935), .o(g62565_sb) );
na02m01 TIMEBOOST_cell_69766 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q), .o(TIMEBOOST_net_22091) );
in01s01 TIMEBOOST_cell_17875 ( .a(TIMEBOOST_net_5286), .o(wbs_dat_i_28_) );
in01s01 TIMEBOOST_cell_17874 ( .a(TIMEBOOST_net_5285), .o(TIMEBOOST_net_5284) );
in01f02 g62566_u0 ( .a(FE_OFN1285_n_4097), .o(g62566_sb) );
na03f02 TIMEBOOST_cell_34873 ( .a(TIMEBOOST_net_9395), .b(FE_OFN1401_n_8567), .c(g57162_sb), .o(n_11588) );
in01s01 TIMEBOOST_cell_17873 ( .a(TIMEBOOST_net_5284), .o(wbs_dat_i_31_) );
in01s01 TIMEBOOST_cell_17872 ( .a(TIMEBOOST_net_5283), .o(TIMEBOOST_net_5282) );
in01f01 g62567_u0 ( .a(FE_OFN1284_n_4097), .o(g62567_sb) );
na02f02 TIMEBOOST_cell_53079 ( .a(TIMEBOOST_net_13231), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_16757) );
in01s01 TIMEBOOST_cell_17871 ( .a(TIMEBOOST_net_5282), .o(wbs_dat_i_15_) );
na02m02 TIMEBOOST_cell_72123 ( .a(TIMEBOOST_net_23269), .b(g65949_sb), .o(n_1562) );
in01m01 g62568_u0 ( .a(FE_OFN1295_n_4098), .o(g62568_sb) );
na03f02 TIMEBOOST_cell_73720 ( .a(n_12010), .b(TIMEBOOST_net_13554), .c(FE_OFN1748_n_12004), .o(n_12605) );
na03f02 TIMEBOOST_cell_65882 ( .a(n_4009), .b(g62789_sb), .c(g62789_db), .o(n_5412) );
in01f02 g62569_u0 ( .a(FE_OFN1315_n_6624), .o(g62569_sb) );
na02m04 TIMEBOOST_cell_68597 ( .a(TIMEBOOST_net_21506), .b(g64830_sb), .o(TIMEBOOST_net_12823) );
na03f02 TIMEBOOST_cell_73241 ( .a(n_3493), .b(g58605_sb), .c(TIMEBOOST_net_15817), .o(n_13552) );
na02s02 TIMEBOOST_cell_49487 ( .a(FE_OFN1649_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q), .o(TIMEBOOST_net_14961) );
in01f02 g62570_u0 ( .a(FE_OFN1234_n_6391), .o(g62570_sb) );
na03f01 TIMEBOOST_cell_72425 ( .a(TIMEBOOST_net_14006), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q), .c(wbu_addr_in_274), .o(n_9120) );
na03f02 TIMEBOOST_cell_72711 ( .a(g64823_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q), .c(TIMEBOOST_net_10520), .o(TIMEBOOST_net_17401) );
in01s03 TIMEBOOST_cell_45965 ( .a(pci_target_unit_fifos_pcir_data_in_180), .o(TIMEBOOST_net_13926) );
in01f02 g62571_u0 ( .a(FE_OFN1314_n_6624), .o(g62571_sb) );
na02s02 TIMEBOOST_cell_49265 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q), .b(FE_OFN540_n_9690), .o(TIMEBOOST_net_14850) );
in01f01 g62572_u0 ( .a(FE_OFN1200_n_4090), .o(g62572_sb) );
na04m02 TIMEBOOST_cell_72793 ( .a(TIMEBOOST_net_21458), .b(g65784_db), .c(TIMEBOOST_net_17238), .d(g61738_sb), .o(n_8341) );
in01s01 TIMEBOOST_cell_17869 ( .a(TIMEBOOST_net_5280), .o(wbs_dat_i_11_) );
in01f02 g62573_u0 ( .a(FE_OFN1196_n_4090), .o(g62573_sb) );
na02s01 TIMEBOOST_cell_17938 ( .a(TIMEBOOST_net_5332), .b(g67049_sb), .o(n_1428) );
na02s01 TIMEBOOST_cell_17937 ( .a(FE_OFN1778_parchk_pci_ad_reg_in_1222), .b(g67074_db), .o(TIMEBOOST_net_5332) );
in01m01 g62574_u0 ( .a(FE_OFN1193_n_6935), .o(g62574_sb) );
na02f08 TIMEBOOST_cell_47796 ( .a(TIMEBOOST_net_14115), .b(n_16539), .o(n_16540) );
in01f01 g62575_u0 ( .a(FE_OFN1192_n_6935), .o(g62575_sb) );
na02f02 TIMEBOOST_cell_49890 ( .a(TIMEBOOST_net_15162), .b(g63437_sb), .o(n_4928) );
na02f02 TIMEBOOST_cell_43895 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q), .b(g64244_sb), .o(TIMEBOOST_net_12842) );
in01f02 g62576_u0 ( .a(FE_OFN1320_n_6436), .o(g62576_sb) );
na03f02 TIMEBOOST_cell_34817 ( .a(TIMEBOOST_net_9425), .b(FE_OFN1380_n_8567), .c(g57099_sb), .o(n_10481) );
na02f02 TIMEBOOST_cell_3802 ( .a(n_15434), .b(n_3032), .o(TIMEBOOST_net_461) );
in01f02 g62577_u0 ( .a(FE_OFN1246_n_4093), .o(g62577_sb) );
na02f02 TIMEBOOST_cell_72079 ( .a(TIMEBOOST_net_23247), .b(g64248_sb), .o(TIMEBOOST_net_13039) );
in01s01 TIMEBOOST_cell_17867 ( .a(TIMEBOOST_net_5278), .o(wbs_dat_i_14_) );
na02s01 TIMEBOOST_cell_48179 ( .a(pci_target_unit_fifos_pcir_data_in_187), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q), .o(TIMEBOOST_net_14307) );
in01f02 g62578_u0 ( .a(FE_OFN1208_n_6356), .o(g62578_sb) );
na02m01 TIMEBOOST_cell_63664 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q), .b(FE_OFN679_n_4460), .o(TIMEBOOST_net_20818) );
in01s01 TIMEBOOST_cell_17868 ( .a(TIMEBOOST_net_5279), .o(TIMEBOOST_net_5278) );
in01s01 TIMEBOOST_cell_17865 ( .a(TIMEBOOST_net_5276), .o(wbs_dat_i_0_) );
in01m01 g62579_u0 ( .a(FE_OFN1208_n_6356), .o(g62579_sb) );
na02s01 TIMEBOOST_cell_48605 ( .a(g61801_sb), .b(g61801_db), .o(TIMEBOOST_net_14520) );
na02f02 g54317_u2 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q), .b(FE_OFN2127_n_16497), .o(g54317_db) );
in01m01 g62580_u0 ( .a(FE_OFN1222_n_6391), .o(g62580_sb) );
na02f01 g62580_u2 ( .a(n_3697), .b(FE_OFN1222_n_6391), .o(g62580_db) );
in01f01 g62581_u0 ( .a(FE_OFN1250_n_4093), .o(g62581_sb) );
na03m02 TIMEBOOST_cell_64512 ( .a(n_3780), .b(FE_OFN614_n_4501), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q), .o(TIMEBOOST_net_16239) );
na03f01 TIMEBOOST_cell_64511 ( .a(FE_OFN679_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q), .c(n_3764), .o(TIMEBOOST_net_14290) );
na04f04 TIMEBOOST_cell_24608 ( .a(n_9435), .b(g57544_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q), .d(FE_OFN2184_n_8567), .o(n_11200) );
in01f01 g62582_u0 ( .a(FE_OFN1194_n_6935), .o(g62582_sb) );
na02m10 TIMEBOOST_cell_52985 ( .a(wishbone_slave_unit_pcim_sm_data_in_651), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q), .o(TIMEBOOST_net_16710) );
na04f04 TIMEBOOST_cell_24610 ( .a(n_9209), .b(g57541_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q), .d(FE_OFN2177_n_8567), .o(n_10813) );
na04f04 TIMEBOOST_cell_24612 ( .a(n_9439), .b(g57536_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q), .d(FE_OFN2177_n_8567), .o(n_11206) );
in01f02 g62583_u0 ( .a(FE_OFN1224_n_6391), .o(g62583_sb) );
in01f02 g62584_u0 ( .a(FE_OFN1293_n_4098), .o(g62584_sb) );
na02s02 TIMEBOOST_cell_63222 ( .a(g58101_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q), .o(TIMEBOOST_net_20558) );
na04f04 TIMEBOOST_cell_24614 ( .a(n_9444), .b(g57528_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q), .d(FE_OFN2182_n_8567), .o(n_11213) );
na04f04 TIMEBOOST_cell_24616 ( .a(n_9008), .b(g57521_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q), .d(FE_OFN2168_n_8567), .o(n_10316) );
in01f01 g62585_u0 ( .a(FE_OFN1294_n_4098), .o(g62585_sb) );
na04f04 TIMEBOOST_cell_24628 ( .a(n_9125), .b(g57074_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q), .d(FE_OFN2169_n_8567), .o(n_10495) );
na04f04 TIMEBOOST_cell_24630 ( .a(n_9874), .b(g57055_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q), .d(FE_OFN2179_n_8567), .o(n_11681) );
in01m01 g62586_u0 ( .a(FE_OFN1213_n_4151), .o(g62586_sb) );
na04f04 TIMEBOOST_cell_24632 ( .a(n_9881), .b(g57049_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q), .d(FE_OFN2190_n_8567), .o(n_11686) );
na04f04 TIMEBOOST_cell_24634 ( .a(n_9891), .b(g57040_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q), .d(FE_OFN2168_n_8567), .o(n_11694) );
in01f02 g62587_u0 ( .a(FE_OFN1202_n_4090), .o(g62587_sb) );
na04f04 TIMEBOOST_cell_24636 ( .a(n_9061), .b(g57313_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q), .d(FE_OFN2169_n_8567), .o(n_10401) );
na04f04 TIMEBOOST_cell_24638 ( .a(n_9649), .b(g57283_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q), .d(FE_OFN2185_n_8567), .o(n_11472) );
in01f02 g62588_u0 ( .a(n_6431), .o(g62588_sb) );
na02m01 TIMEBOOST_cell_68616 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q), .o(TIMEBOOST_net_21516) );
na02s02 TIMEBOOST_cell_49488 ( .a(TIMEBOOST_net_14961), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_11196) );
in01f01 g62589_u0 ( .a(FE_OFN1194_n_6935), .o(g62589_sb) );
na02s02 TIMEBOOST_cell_38017 ( .a(g58152_sb), .b(TIMEBOOST_net_10620), .o(n_9068) );
na04f04 TIMEBOOST_cell_24640 ( .a(n_9072), .b(g57271_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q), .d(FE_OFN2170_n_8567), .o(n_10416) );
na04f04 TIMEBOOST_cell_24642 ( .a(n_9671), .b(g57259_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q), .d(FE_OFN2187_n_8567), .o(n_11495) );
in01f02 g62590_u0 ( .a(FE_OFN1206_n_6356), .o(g62590_sb) );
na02s01 TIMEBOOST_cell_53969 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_17202) );
na04f02 TIMEBOOST_cell_66469 ( .a(TIMEBOOST_net_15684), .b(g53942_db), .c(n_2692), .d(g63193_sb), .o(n_13503) );
in01f04 TIMEBOOST_cell_17851 ( .a(TIMEBOOST_net_5262), .o(n_2319) );
in01f02 g62591_u0 ( .a(FE_OFN1242_n_4092), .o(g62591_sb) );
in01s01 TIMEBOOST_cell_17880 ( .a(TIMEBOOST_net_5291), .o(TIMEBOOST_net_5290) );
in01s01 TIMEBOOST_cell_17863 ( .a(TIMEBOOST_net_5274), .o(wbs_dat_i_8_) );
in01m01 g62592_u0 ( .a(FE_OFN1283_n_4097), .o(g62592_sb) );
na03f02 TIMEBOOST_cell_34808 ( .a(TIMEBOOST_net_9508), .b(FE_OFN1413_n_8567), .c(g57135_sb), .o(n_10467) );
in01f02 g62593_u0 ( .a(FE_OFN1311_n_6624), .o(g62593_sb) );
na02f02 TIMEBOOST_cell_3803 ( .a(TIMEBOOST_net_461), .b(n_15699), .o(n_4857) );
in01f02 g62594_u0 ( .a(FE_OFN1203_n_4090), .o(g62594_sb) );
in01m01 TIMEBOOST_cell_45987 ( .a(pci_target_unit_fifos_pcir_data_in_163), .o(TIMEBOOST_net_13948) );
na04f04 TIMEBOOST_cell_24560 ( .a(n_9204), .b(g57556_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q), .d(FE_OFN1417_n_8567), .o(n_10804) );
na03s01 TIMEBOOST_cell_72565 ( .a(pci_target_unit_del_sync_addr_in_226), .b(g66402_sb), .c(g66402_db), .o(n_2539) );
no02f04 g62595_u0 ( .a(conf_wb_err_addr_in_968), .b(n_2915), .o(g62595_p) );
ao12f02 g62595_u1 ( .a(g62595_p), .b(conf_wb_err_addr_in_968), .c(n_2915), .o(n_3467) );
in01f01 g62596_u0 ( .a(FE_OFN1294_n_4098), .o(g62596_sb) );
na03f02 TIMEBOOST_cell_47287 ( .a(FE_OFN1734_n_16317), .b(TIMEBOOST_net_13584), .c(FE_OFN1739_n_11019), .o(n_12671) );
na03f02 TIMEBOOST_cell_35056 ( .a(TIMEBOOST_net_9608), .b(FE_OFN1439_n_9372), .c(g58478_sb), .o(n_9361) );
in01f01 g62597_u0 ( .a(FE_OFN1207_n_6356), .o(g62597_sb) );
na03s02 TIMEBOOST_cell_33796 ( .a(n_2195), .b(g61715_sb), .c(g61715_db), .o(n_8395) );
in01s01 TIMEBOOST_cell_17861 ( .a(parchk_pci_ad_out_in_1172), .o(TIMEBOOST_net_5272) );
in01s01 TIMEBOOST_cell_17862 ( .a(TIMEBOOST_net_5272), .o(TIMEBOOST_net_5273) );
in01m01 g62598_u0 ( .a(FE_OFN1207_n_6356), .o(g62598_sb) );
na03f02 TIMEBOOST_cell_67985 ( .a(TIMEBOOST_net_17368), .b(FE_OFN1248_n_4093), .c(g62556_sb), .o(n_6451) );
na02m04 TIMEBOOST_cell_69915 ( .a(TIMEBOOST_net_22165), .b(g64192_sb), .o(n_3976) );
na03f02 TIMEBOOST_cell_35058 ( .a(TIMEBOOST_net_9609), .b(FE_OFN1436_n_9372), .c(g58462_sb), .o(n_9391) );
in01f02 g62599_u0 ( .a(FE_OFN1312_n_6624), .o(g62599_sb) );
na03m02 TIMEBOOST_cell_64727 ( .a(FE_OFN662_n_4392), .b(n_84), .c(n_3770), .o(TIMEBOOST_net_10596) );
in01f04 g62600_u0 ( .a(FE_OFN1314_n_6624), .o(g62600_sb) );
na02m01 TIMEBOOST_cell_38225 ( .a(TIMEBOOST_net_10724), .b(TIMEBOOST_net_5434), .o(n_2649) );
in01f02 g62601_u0 ( .a(FE_OFN1236_n_6391), .o(g62601_sb) );
na02f04 TIMEBOOST_cell_3519 ( .a(TIMEBOOST_net_319), .b(FE_RN_704_0), .o(FE_RN_705_0) );
na02s01 TIMEBOOST_cell_3520 ( .a(n_4869), .b(n_15856), .o(TIMEBOOST_net_320) );
in01m01 g62602_u0 ( .a(FE_OFN1218_n_6886), .o(g62602_sb) );
na03f02 TIMEBOOST_cell_67040 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_16535), .c(FE_OFN1600_n_13995), .o(n_16249) );
na02s02 TIMEBOOST_cell_17932 ( .a(TIMEBOOST_net_5329), .b(n_1989), .o(TIMEBOOST_net_80) );
na02s01 TIMEBOOST_cell_17931 ( .a(pci_target_unit_del_sync_comp_cycle_count_9_), .b(pci_target_unit_del_sync_comp_cycle_count_10_), .o(TIMEBOOST_net_5329) );
in01f02 g62603_u0 ( .a(FE_OFN1218_n_6886), .o(g62603_sb) );
na03f02 TIMEBOOST_cell_73513 ( .a(TIMEBOOST_net_17048), .b(n_6232), .c(g62478_sb), .o(n_6631) );
na02s01 TIMEBOOST_cell_18158 ( .a(TIMEBOOST_net_5442), .b(g65813_sb), .o(n_2571) );
na02f02 TIMEBOOST_cell_17930 ( .a(TIMEBOOST_net_5328), .b(n_937), .o(TIMEBOOST_net_262) );
in01f01 g62604_u0 ( .a(FE_OFN1253_n_4143), .o(g62604_sb) );
in01s01 TIMEBOOST_cell_17860 ( .a(TIMEBOOST_net_5270), .o(TIMEBOOST_net_5271) );
in01s01 TIMEBOOST_cell_17859 ( .a(conf_wb_err_addr_in_944), .o(TIMEBOOST_net_5270) );
in01f02 g62605_u0 ( .a(FE_OFN1223_n_6391), .o(g62605_sb) );
na02f02 TIMEBOOST_cell_3313 ( .a(TIMEBOOST_net_216), .b(FE_RN_356_0), .o(n_5747) );
in01s01 TIMEBOOST_cell_73892 ( .a(n_8229), .o(TIMEBOOST_net_23457) );
in01f02 g62606_u0 ( .a(FE_OFN1233_n_6391), .o(g62606_sb) );
na02s01 TIMEBOOST_cell_51651 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q), .o(TIMEBOOST_net_16043) );
na02f02 TIMEBOOST_cell_3521 ( .a(TIMEBOOST_net_320), .b(n_4818), .o(n_7538) );
in01f01 g62607_u0 ( .a(n_4098), .o(g62607_sb) );
na02f03 TIMEBOOST_cell_72125 ( .a(TIMEBOOST_net_23270), .b(g65900_sb), .o(n_1571) );
na03m02 TIMEBOOST_cell_66082 ( .a(TIMEBOOST_net_20479), .b(FE_OFN1632_n_9531), .c(g58392_sb), .o(n_9006) );
in01f01 g62608_u0 ( .a(FE_OFN1294_n_4098), .o(g62608_sb) );
na02s01 TIMEBOOST_cell_44453 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q), .b(FE_OFN539_n_9690), .o(TIMEBOOST_net_13121) );
in01s01 TIMEBOOST_cell_17858 ( .a(TIMEBOOST_net_5268), .o(TIMEBOOST_net_5269) );
in01s01 TIMEBOOST_cell_17857 ( .a(conf_wb_err_addr_in_954), .o(TIMEBOOST_net_5268) );
in01m01 g62609_u0 ( .a(FE_OFN1241_n_4092), .o(g62609_sb) );
na04f02 TIMEBOOST_cell_73625 ( .a(n_16748), .b(pci_target_unit_pcit_if_strd_addr_in_713), .c(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77), .d(g52642_sb), .o(TIMEBOOST_net_13487) );
na02s04 TIMEBOOST_cell_17929 ( .a(pci_target_unit_del_sync_comp_cycle_count_11_), .b(pci_target_unit_del_sync_comp_cycle_count_10_), .o(TIMEBOOST_net_5328) );
na02m03 TIMEBOOST_cell_17928 ( .a(TIMEBOOST_net_5327), .b(n_929), .o(TIMEBOOST_net_40) );
in01f02 g62610_u0 ( .a(FE_OFN1200_n_4090), .o(g62610_sb) );
na04m02 TIMEBOOST_cell_72794 ( .a(n_4476), .b(g64812_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q), .d(TIMEBOOST_net_20280), .o(TIMEBOOST_net_17096) );
in01f02 TIMEBOOST_cell_17850 ( .a(TIMEBOOST_net_5261), .o(TIMEBOOST_net_5260) );
na03f02 TIMEBOOST_cell_35060 ( .a(TIMEBOOST_net_9590), .b(FE_OFN1440_n_9372), .c(g58471_sb), .o(n_9374) );
in01f01 g62611_u0 ( .a(FE_OFN1222_n_6391), .o(g62611_sb) );
na02f06 TIMEBOOST_cell_3315 ( .a(TIMEBOOST_net_217), .b(n_2485), .o(n_3195) );
na02f02 g62611_u2 ( .a(n_3740), .b(FE_OFN1222_n_6391), .o(g62611_db) );
na03f02 TIMEBOOST_cell_34868 ( .a(TIMEBOOST_net_9343), .b(FE_OFN1420_n_8567), .c(g57338_sb), .o(n_11414) );
in01f02 g62612_u0 ( .a(FE_OFN1315_n_6624), .o(g62612_sb) );
in01f02 g62613_u0 ( .a(FE_OFN1197_n_4090), .o(g62613_sb) );
na03m06 TIMEBOOST_cell_72741 ( .a(n_4498), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q), .c(FE_OFN636_n_4669), .o(TIMEBOOST_net_10617) );
in01f04 TIMEBOOST_cell_17849 ( .a(TIMEBOOST_net_5260), .o(n_2464) );
in01s01 TIMEBOOST_cell_17864 ( .a(TIMEBOOST_net_5275), .o(TIMEBOOST_net_5274) );
in01f02 g62614_u0 ( .a(FE_OFN1233_n_6391), .o(g62614_sb) );
na04m04 TIMEBOOST_cell_67455 ( .a(TIMEBOOST_net_20354), .b(FE_OFN1628_n_4438), .c(g64985_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q), .o(TIMEBOOST_net_13248) );
na02f06 TIMEBOOST_cell_3523 ( .a(n_3107), .b(TIMEBOOST_net_321), .o(n_8476) );
na02m06 TIMEBOOST_cell_3524 ( .a(n_2596), .b(n_2872), .o(TIMEBOOST_net_322) );
in01f01 g62615_u0 ( .a(FE_OFN1272_n_4096), .o(g62615_sb) );
na03f02 TIMEBOOST_cell_65690 ( .a(TIMEBOOST_net_12876), .b(FE_OFN2126_n_16497), .c(g54331_sb), .o(n_12985) );
in01m01 TIMEBOOST_cell_17856 ( .a(TIMEBOOST_net_5266), .o(TIMEBOOST_net_5267) );
na02m02 TIMEBOOST_cell_17927 ( .a(pci_target_unit_wishbone_master_rty_counter_5_), .b(pci_target_unit_wishbone_master_rty_counter_6_), .o(TIMEBOOST_net_5327) );
in01f04 g62616_u0 ( .a(FE_OFN1214_n_4151), .o(g62616_sb) );
na03m02 TIMEBOOST_cell_68894 ( .a(n_4482), .b(g64758_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q), .o(TIMEBOOST_net_21655) );
na02f01 TIMEBOOST_cell_17926 ( .a(TIMEBOOST_net_5326), .b(n_948), .o(TIMEBOOST_net_30) );
in01m02 TIMEBOOST_cell_17855 ( .a(conf_wb_err_addr_in_951), .o(TIMEBOOST_net_5266) );
in01f01 g62617_u0 ( .a(FE_OFN1200_n_4090), .o(g62617_sb) );
na03f02 TIMEBOOST_cell_34951 ( .a(TIMEBOOST_net_9499), .b(FE_OFN1399_n_8567), .c(g57269_sb), .o(n_11483) );
na02s03 TIMEBOOST_cell_17925 ( .a(pci_target_unit_del_sync_comp_cycle_count_5_), .b(pci_target_unit_del_sync_comp_cycle_count_2_), .o(TIMEBOOST_net_5326) );
in01m02 TIMEBOOST_cell_17854 ( .a(TIMEBOOST_net_5265), .o(TIMEBOOST_net_5264) );
in01f02 g62618_u0 ( .a(FE_OFN1320_n_6436), .o(g62618_sb) );
in01s01 TIMEBOOST_cell_67730 ( .a(TIMEBOOST_net_21156), .o(TIMEBOOST_net_21157) );
na04f04 TIMEBOOST_cell_24180 ( .a(n_9197), .b(g57506_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q), .d(FE_OFN1416_n_8567), .o(n_10815) );
in01f02 g62619_u0 ( .a(n_6319), .o(g62619_sb) );
na02s02 TIMEBOOST_cell_39735 ( .a(TIMEBOOST_net_11479), .b(g57892_db), .o(n_9232) );
in01f01 g62620_u0 ( .a(FE_OFN1276_n_4096), .o(g62620_sb) );
na03f02 TIMEBOOST_cell_72795 ( .a(TIMEBOOST_net_23166), .b(g65011_sb), .c(TIMEBOOST_net_22117), .o(TIMEBOOST_net_9947) );
na02s02 TIMEBOOST_cell_17924 ( .a(TIMEBOOST_net_5325), .b(n_1989), .o(TIMEBOOST_net_180) );
na02s01 TIMEBOOST_cell_2892 ( .a(pci_target_unit_wishbone_master_burst_chopped), .b(n_1183), .o(TIMEBOOST_net_6) );
in01f01 g62621_u0 ( .a(FE_OFN1294_n_4098), .o(g62621_sb) );
na02s01 TIMEBOOST_cell_2893 ( .a(TIMEBOOST_net_6), .b(n_898), .o(n_1185) );
na02s01 TIMEBOOST_cell_2894 ( .a(n_705), .b(pci_target_unit_wishbone_master_first_wb_data_access), .o(TIMEBOOST_net_7) );
in01f02 g62622_u0 ( .a(FE_OFN1315_n_6624), .o(g62622_sb) );
na02m01 TIMEBOOST_cell_64138 ( .a(n_8272), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_21055) );
na02m08 TIMEBOOST_cell_70747 ( .a(TIMEBOOST_net_22581), .b(FE_OFN535_n_9823), .o(TIMEBOOST_net_14386) );
na03f02 TIMEBOOST_cell_66742 ( .a(TIMEBOOST_net_17373), .b(FE_OFN1279_n_4097), .c(g63163_sb), .o(n_5810) );
in01f02 g62623_u0 ( .a(FE_OFN1235_n_6391), .o(g62623_sb) );
na03f02 TIMEBOOST_cell_73242 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_788), .b(g54312_sb), .c(TIMEBOOST_net_323), .o(n_13295) );
na02m08 TIMEBOOST_cell_3525 ( .a(n_2873), .b(TIMEBOOST_net_322), .o(n_2874) );
na02s01 TIMEBOOST_cell_38596 ( .a(g58014_sb), .b(FE_OFN215_n_9856), .o(TIMEBOOST_net_10910) );
in01f02 g62624_u0 ( .a(FE_OFN1218_n_6886), .o(g62624_sb) );
na03f02 TIMEBOOST_cell_34963 ( .a(TIMEBOOST_net_9466), .b(FE_OFN1374_n_8567), .c(g57520_sb), .o(n_11220) );
na02f01 TIMEBOOST_cell_68497 ( .a(TIMEBOOST_net_21456), .b(g66397_sb), .o(n_2546) );
na03m04 TIMEBOOST_cell_73168 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q), .b(g64312_sb), .c(g64312_db), .o(n_3863) );
in01f02 g62625_u0 ( .a(FE_OFN1234_n_6391), .o(g62625_sb) );
na04f04 TIMEBOOST_cell_73006 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q), .b(TIMEBOOST_net_12695), .c(g65966_sb), .d(FE_OFN713_n_8140), .o(TIMEBOOST_net_16951) );
in01f02 g62626_u0 ( .a(FE_OFN1232_n_6391), .o(g62626_sb) );
na03f02 TIMEBOOST_cell_73687 ( .a(n_14661), .b(n_8757), .c(g52443_da), .o(n_14808) );
in01f02 g62627_u0 ( .a(FE_OFN1236_n_6391), .o(g62627_sb) );
na02m02 TIMEBOOST_cell_49209 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q), .b(g65815_sb), .o(TIMEBOOST_net_14822) );
na03f02 TIMEBOOST_cell_34810 ( .a(TIMEBOOST_net_9393), .b(FE_OFN1374_n_8567), .c(g57254_sb), .o(n_11500) );
in01m01 g62628_u0 ( .a(FE_OFN1283_n_4097), .o(g62628_sb) );
na02s01 TIMEBOOST_cell_64194 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q), .o(TIMEBOOST_net_21083) );
in01f02 g62629_u0 ( .a(FE_OFN1213_n_4151), .o(g62629_sb) );
na03m02 TIMEBOOST_cell_69628 ( .a(FE_OFN1643_n_4671), .b(n_3777), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q), .o(TIMEBOOST_net_22022) );
in01f02 g62630_u0 ( .a(n_6232), .o(g62630_sb) );
in01f02 g62631_u0 ( .a(FE_OFN1253_n_4143), .o(g62631_sb) );
na03m02 TIMEBOOST_cell_69770 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(FE_OFN927_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_22093) );
na02s01 TIMEBOOST_cell_2895 ( .a(TIMEBOOST_net_7), .b(n_1183), .o(n_2027) );
na03m04 TIMEBOOST_cell_73126 ( .a(FE_OFN1077_n_4740), .b(TIMEBOOST_net_17273), .c(g64211_sb), .o(n_3958) );
in01f02 g62632_u0 ( .a(n_6287), .o(g62632_sb) );
na02s02 TIMEBOOST_cell_43626 ( .a(TIMEBOOST_net_12707), .b(TIMEBOOST_net_10528), .o(TIMEBOOST_net_9384) );
na02s01 TIMEBOOST_cell_42883 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q), .o(TIMEBOOST_net_12336) );
in01f02 g62633_u0 ( .a(FE_OFN1323_n_6436), .o(g62633_sb) );
na03f02 TIMEBOOST_cell_73243 ( .a(n_2770), .b(g59121_sb), .c(TIMEBOOST_net_16463), .o(n_13504) );
in01f02 g62634_u0 ( .a(FE_OFN1223_n_6391), .o(g62634_sb) );
in01s01 TIMEBOOST_cell_63574 ( .a(pci_target_unit_fifos_pcir_data_in_172), .o(TIMEBOOST_net_20754) );
na02m02 TIMEBOOST_cell_49247 ( .a(g58406_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q), .o(TIMEBOOST_net_14841) );
in01f02 g62635_u0 ( .a(FE_OFN1315_n_6624), .o(g62635_sb) );
na03s02 TIMEBOOST_cell_66582 ( .a(TIMEBOOST_net_20604), .b(g58487_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q), .o(TIMEBOOST_net_9565) );
na03f02 TIMEBOOST_cell_67988 ( .a(TIMEBOOST_net_21033), .b(FE_OFN1293_n_4098), .c(g62584_sb), .o(n_6384) );
in01f02 g62636_u0 ( .a(FE_OFN1322_n_6436), .o(g62636_sb) );
na04f02 TIMEBOOST_cell_73391 ( .a(configuration_pci_err_addr_480), .b(FE_OFN1186_n_3476), .c(wbm_adr_o_10_), .d(g60605_sb), .o(n_4849) );
na02m10 TIMEBOOST_cell_54513 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_9__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_392), .o(TIMEBOOST_net_17474) );
in01s01 TIMEBOOST_cell_67779 ( .a(TIMEBOOST_net_21206), .o(pci_target_unit_fifos_pcir_data_in_182) );
in01m02 g62637_u0 ( .a(FE_OFN1289_n_4098), .o(g62637_sb) );
na02f04 TIMEBOOST_cell_69583 ( .a(TIMEBOOST_net_21999), .b(g63530_sb), .o(n_3429) );
na02m01 TIMEBOOST_cell_3233 ( .a(TIMEBOOST_net_176), .b(g60688_sb), .o(n_3524) );
in01f01 g62638_u0 ( .a(FE_OFN1248_n_4093), .o(g62638_sb) );
na02f01 TIMEBOOST_cell_54181 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q), .b(FE_OFN1074_n_4740), .o(TIMEBOOST_net_17308) );
in01f02 g62639_u0 ( .a(FE_OFN1293_n_4098), .o(g62639_sb) );
na03f02 TIMEBOOST_cell_68356 ( .a(FE_OFN905_n_4736), .b(TIMEBOOST_net_20175), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q), .o(TIMEBOOST_net_21386) );
na02m01 TIMEBOOST_cell_47818 ( .a(TIMEBOOST_net_14126), .b(g60688_sb), .o(TIMEBOOST_net_13043) );
na03m01 TIMEBOOST_cell_64415 ( .a(TIMEBOOST_net_20793), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_411), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q), .o(TIMEBOOST_net_16796) );
in01m01 g62640_u0 ( .a(FE_OFN1225_n_6391), .o(g62640_sb) );
na02f02 g59230_u2 ( .a(n_3350), .b(FE_OFN1699_n_5751), .o(g59230_db) );
in01f01 g62641_u0 ( .a(FE_OFN1276_n_4096), .o(g62641_sb) );
na04m02 TIMEBOOST_cell_72746 ( .a(n_4498), .b(FE_OFN1644_n_4671), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q), .d(g65370_sb), .o(n_4519) );
na02f02 TIMEBOOST_cell_50520 ( .a(TIMEBOOST_net_15477), .b(g62891_sb), .o(n_6095) );
no02s01 TIMEBOOST_cell_2898 ( .a(n_23), .b(wbs_bte_i_1_), .o(TIMEBOOST_net_9) );
in01m01 g62642_u0 ( .a(FE_OFN1241_n_4092), .o(g62642_sb) );
na02f02 TIMEBOOST_cell_71617 ( .a(TIMEBOOST_net_23016), .b(FE_OFN1757_n_12681), .o(n_12481) );
in01f01 g62643_u0 ( .a(FE_OFN1243_n_4092), .o(g62643_sb) );
na03f02 TIMEBOOST_cell_34949 ( .a(TIMEBOOST_net_9541), .b(FE_OFN1420_n_8567), .c(g57306_sb), .o(n_11445) );
na03f02 TIMEBOOST_cell_73688 ( .a(TIMEBOOST_net_22948), .b(TIMEBOOST_net_8580), .c(TIMEBOOST_net_22956), .o(n_14826) );
na02m02 TIMEBOOST_cell_68604 ( .a(g65083_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q), .o(TIMEBOOST_net_21510) );
in01f02 g62644_u0 ( .a(FE_OFN1233_n_6391), .o(g62644_sb) );
na02f02 TIMEBOOST_cell_72239 ( .a(TIMEBOOST_net_23327), .b(g63170_sb), .o(n_4953) );
na02f04 TIMEBOOST_cell_3532 ( .a(FE_OCP_RBN2231_FE_RN_390_0), .b(n_15914), .o(TIMEBOOST_net_326) );
in01f02 g62645_u0 ( .a(FE_OFN1284_n_4097), .o(g62645_sb) );
na02m02 TIMEBOOST_cell_3241 ( .a(n_2420), .b(TIMEBOOST_net_180), .o(n_2491) );
na02m10 TIMEBOOST_cell_47953 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q), .o(TIMEBOOST_net_14194) );
in01f02 g62646_u0 ( .a(FE_OFN1234_n_6391), .o(g62646_sb) );
na03f02 TIMEBOOST_cell_67986 ( .a(TIMEBOOST_net_20524), .b(FE_OFN1293_n_4098), .c(g62483_sb), .o(n_6621) );
na02f08 TIMEBOOST_cell_3533 ( .a(n_15910), .b(TIMEBOOST_net_326), .o(n_15915) );
na02s01 TIMEBOOST_cell_3534 ( .a(n_5757), .b(n_15741), .o(TIMEBOOST_net_327) );
in01f02 g62647_u0 ( .a(n_6431), .o(g62647_sb) );
na02m06 TIMEBOOST_cell_45605 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q), .o(TIMEBOOST_net_13697) );
in01m01 g62648_u0 ( .a(FE_OFN1224_n_6391), .o(g62648_sb) );
na03f02 TIMEBOOST_cell_73721 ( .a(TIMEBOOST_net_11884), .b(g52650_db), .c(TIMEBOOST_net_22988), .o(n_14838) );
na04f04 TIMEBOOST_cell_67434 ( .a(n_3598), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q), .c(FE_OFN1232_n_6391), .d(g62626_sb), .o(n_6303) );
na02s01 TIMEBOOST_cell_43079 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_12434) );
in01f02 g62649_u0 ( .a(FE_OFN1223_n_6391), .o(g62649_sb) );
na03f02 TIMEBOOST_cell_67043 ( .a(FE_OFN1605_n_13997), .b(TIMEBOOST_net_8615), .c(FE_OFN1601_n_13995), .o(FE_RN_893_0) );
in01f01 g62650_u0 ( .a(FE_OFN1272_n_4096), .o(g62650_sb) );
na02s02 TIMEBOOST_cell_50058 ( .a(TIMEBOOST_net_15246), .b(TIMEBOOST_net_10348), .o(TIMEBOOST_net_9433) );
na02f02 TIMEBOOST_cell_54358 ( .a(TIMEBOOST_net_17396), .b(FE_OFN1203_n_4090), .o(TIMEBOOST_net_15718) );
in01f02 g62651_u0 ( .a(FE_OFN1200_n_4090), .o(g62651_sb) );
in01s01 TIMEBOOST_cell_73846 ( .a(n_7400), .o(TIMEBOOST_net_23411) );
na02s01 TIMEBOOST_cell_2904 ( .a(n_705), .b(pci_target_unit_wishbone_master_rty_counter_0_), .o(TIMEBOOST_net_12) );
in01f01 g62652_u0 ( .a(FE_OFN1242_n_4092), .o(g62652_sb) );
na02f02 TIMEBOOST_cell_53645 ( .a(TIMEBOOST_net_13246), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_17040) );
in01f01 g62653_u0 ( .a(FE_OFN1193_n_6935), .o(g62653_sb) );
na03f02 TIMEBOOST_cell_70298 ( .a(TIMEBOOST_net_17285), .b(FE_OFN1148_n_13249), .c(n_2121), .o(TIMEBOOST_net_22357) );
na02f01 TIMEBOOST_cell_2906 ( .a(n_707), .b(wishbone_slave_unit_pci_initiator_sm_transfer), .o(TIMEBOOST_net_13) );
na02s01 TIMEBOOST_cell_45447 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q), .o(TIMEBOOST_net_13618) );
in01f02 g62654_u0 ( .a(n_6645), .o(g62654_sb) );
in01f02 g62655_u0 ( .a(n_6232), .o(g62655_sb) );
na03m02 TIMEBOOST_cell_71298 ( .a(g58368_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q), .c(FE_OFN1668_n_9477), .o(TIMEBOOST_net_22857) );
na02s02 TIMEBOOST_cell_48718 ( .a(TIMEBOOST_net_14576), .b(TIMEBOOST_net_10442), .o(TIMEBOOST_net_9389) );
in01f02 g62656_u0 ( .a(FE_OFN1235_n_6391), .o(g62656_sb) );
na02f04 TIMEBOOST_cell_3535 ( .a(TIMEBOOST_net_327), .b(n_4809), .o(n_5758) );
na02m02 g64912_u2 ( .a(n_4399), .b(FE_OFN623_n_4409), .o(g64912_db) );
in01f01 g62657_u0 ( .a(FE_OFN1247_n_4093), .o(g62657_sb) );
na02s01 TIMEBOOST_cell_71428 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q), .o(TIMEBOOST_net_22922) );
in01m01 g62658_u0 ( .a(FE_OFN1249_n_4093), .o(g62658_sb) );
na02m08 TIMEBOOST_cell_45399 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q), .o(TIMEBOOST_net_13594) );
na02m02 TIMEBOOST_cell_71299 ( .a(TIMEBOOST_net_22857), .b(FE_OFN272_n_9828), .o(n_9458) );
na02f01 TIMEBOOST_cell_71967 ( .a(TIMEBOOST_net_23191), .b(FE_OFN643_n_4677), .o(TIMEBOOST_net_14513) );
in01f01 g62659_u0 ( .a(FE_OFN1212_n_4151), .o(g62659_sb) );
na03s01 TIMEBOOST_cell_20866 ( .a(n_8876), .b(g56933_sb), .c(pci_target_unit_fifos_pcir_flush_in), .o(TIMEBOOST_net_418) );
na03f02 TIMEBOOST_cell_70420 ( .a(n_4010), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q), .c(FE_OFN1138_g64577_p), .o(TIMEBOOST_net_22418) );
in01f04 g62660_u0 ( .a(FE_OFN1311_n_6624), .o(g62660_sb) );
na02s01 TIMEBOOST_cell_53011 ( .a(configuration_pci_err_data_531), .b(wbm_dat_o_30_), .o(TIMEBOOST_net_16723) );
na03m02 TIMEBOOST_cell_72482 ( .a(TIMEBOOST_net_23130), .b(FE_OFN903_n_4736), .c(g64196_sb), .o(TIMEBOOST_net_13104) );
in01m01 g62661_u0 ( .a(FE_OFN1283_n_4097), .o(g62661_sb) );
na02s01 g65775_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q), .b(FE_OFN937_n_2292), .o(g65775_db) );
in01m10 TIMEBOOST_cell_45929 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .o(TIMEBOOST_net_13890) );
in01f02 g62662_u0 ( .a(FE_OFN1231_n_6391), .o(g62662_sb) );
na02s02 TIMEBOOST_cell_48315 ( .a(FE_OFN572_n_9502), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q), .o(TIMEBOOST_net_14375) );
na02f01 TIMEBOOST_cell_3538 ( .a(g64835_db), .b(n_6935), .o(TIMEBOOST_net_329) );
in01f04 g62663_u0 ( .a(FE_OFN1311_n_6624), .o(g62663_sb) );
in01f02 g62664_u0 ( .a(n_6287), .o(g62664_sb) );
na03s02 TIMEBOOST_cell_72585 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q), .b(TIMEBOOST_net_20576), .c(FE_OFN231_n_9839), .o(TIMEBOOST_net_16454) );
na02f04 TIMEBOOST_cell_69919 ( .a(TIMEBOOST_net_22167), .b(n_16543), .o(TIMEBOOST_net_11894) );
in01f01 g62665_u0 ( .a(FE_OFN1269_n_4095), .o(g62665_sb) );
in01f02 g62666_u0 ( .a(FE_OFN1314_n_6624), .o(g62666_sb) );
na02s02 TIMEBOOST_cell_52472 ( .a(TIMEBOOST_net_16453), .b(TIMEBOOST_net_12817), .o(TIMEBOOST_net_9426) );
na03m02 TIMEBOOST_cell_69154 ( .a(TIMEBOOST_net_20263), .b(FE_OFN928_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q), .o(TIMEBOOST_net_21785) );
in01f02 g62667_u0 ( .a(FE_OFN1293_n_4098), .o(g62667_sb) );
na03f02 TIMEBOOST_cell_73669 ( .a(TIMEBOOST_net_17159), .b(FE_OFN1248_n_4093), .c(g62893_sb), .o(n_6091) );
in01f01 g62668_u0 ( .a(FE_OFN1285_n_4097), .o(g62668_sb) );
no04f80 TIMEBOOST_cell_20870 ( .a(FE_RN_57_0), .b(FE_RN_58_0), .c(wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_), .d(wishbone_slave_unit_fifos_outGreyCount_2_), .o(n_15735) );
in01f01 g62669_u0 ( .a(FE_OFN1202_n_4090), .o(g62669_sb) );
na03f80 TIMEBOOST_cell_20871 ( .a(n_15314), .b(n_16818), .c(n_15317), .o(n_15414) );
na03f02 TIMEBOOST_cell_73689 ( .a(TIMEBOOST_net_22949), .b(TIMEBOOST_net_13489), .c(TIMEBOOST_net_22955), .o(n_14841) );
na02f04 TIMEBOOST_cell_2922 ( .a(conf_wb_err_addr_in_954), .b(conf_wb_err_addr_in_955), .o(TIMEBOOST_net_21) );
in01f01 g62670_u0 ( .a(FE_OFN1247_n_4093), .o(g62670_sb) );
na03f02 TIMEBOOST_cell_34947 ( .a(TIMEBOOST_net_9501), .b(FE_OFN1368_n_8567), .c(g57091_sb), .o(n_10489) );
na02f20 TIMEBOOST_cell_2923 ( .a(TIMEBOOST_net_21), .b(n_913), .o(n_2750) );
na02m01 TIMEBOOST_cell_2924 ( .a(wbm_adr_o_29_), .b(wbm_adr_o_30_), .o(TIMEBOOST_net_22) );
in01m01 g62671_u0 ( .a(FE_OFN1270_n_4095), .o(g62671_sb) );
na03f02 TIMEBOOST_cell_34803 ( .a(TIMEBOOST_net_9552), .b(FE_OFN1411_n_8567), .c(g57419_sb), .o(n_11320) );
na02f02 TIMEBOOST_cell_2925 ( .a(n_879), .b(TIMEBOOST_net_22), .o(n_880) );
na02m01 TIMEBOOST_cell_2926 ( .a(wbm_adr_o_28_), .b(wbm_adr_o_29_), .o(TIMEBOOST_net_23) );
in01f01 g62672_u0 ( .a(FE_OFN1261_n_4143), .o(g62672_sb) );
na02m02 TIMEBOOST_cell_2927 ( .a(n_875), .b(TIMEBOOST_net_23), .o(n_876) );
na03m02 TIMEBOOST_cell_64509 ( .a(n_3752), .b(FE_OFN644_n_4677), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q), .o(TIMEBOOST_net_14514) );
in01f02 g62673_u0 ( .a(FE_OFN1312_n_6624), .o(g62673_sb) );
na03f20 TIMEBOOST_cell_31950 ( .a(TIMEBOOST_net_8634), .b(n_8511), .c(n_1074), .o(n_2440) );
na02m02 TIMEBOOST_cell_37572 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q), .b(FE_OFN622_n_4409), .o(TIMEBOOST_net_10398) );
na02m06 TIMEBOOST_cell_68738 ( .a(FE_OFN682_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_21577) );
in01m01 g62674_u0 ( .a(FE_OFN1249_n_4093), .o(g62674_sb) );
na03f02 TIMEBOOST_cell_66471 ( .a(TIMEBOOST_net_16785), .b(FE_OFN1311_n_6624), .c(g62593_sb), .o(n_6366) );
na02m04 TIMEBOOST_cell_68389 ( .a(TIMEBOOST_net_21402), .b(g65291_sb), .o(TIMEBOOST_net_16156) );
na03f02 TIMEBOOST_cell_73751 ( .a(TIMEBOOST_net_16039), .b(n_12099), .c(FE_OFN1756_n_12681), .o(n_12496) );
in01f02 g62675_u0 ( .a(FE_OFN1202_n_4090), .o(g62675_sb) );
na02m10 TIMEBOOST_cell_45607 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q), .o(TIMEBOOST_net_13698) );
in01f02 g62676_u0 ( .a(FE_OFN365_n_4093), .o(g62676_sb) );
na02s01 TIMEBOOST_cell_38211 ( .a(TIMEBOOST_net_10717), .b(TIMEBOOST_net_8732), .o(n_9491) );
in01f02 g62677_u0 ( .a(n_6554), .o(g62677_sb) );
na02f20 TIMEBOOST_cell_49371 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_782), .o(TIMEBOOST_net_14903) );
in01s01 TIMEBOOST_cell_67744 ( .a(TIMEBOOST_net_21170), .o(TIMEBOOST_net_21171) );
in01f02 g62678_u0 ( .a(FE_OFN1268_n_4095), .o(g62678_sb) );
na03f02 TIMEBOOST_cell_73019 ( .a(TIMEBOOST_net_12716), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .c(g52652_sb), .o(n_14734) );
na02m06 TIMEBOOST_cell_3223 ( .a(n_2473), .b(TIMEBOOST_net_171), .o(n_2474) );
na03f02 TIMEBOOST_cell_73752 ( .a(TIMEBOOST_net_13594), .b(FE_OCPN1827_n_14995), .c(FE_OFN1553_n_12104), .o(n_12746) );
in01f02 g62679_u0 ( .a(FE_OFN1230_n_6391), .o(g62679_sb) );
na02s02 TIMEBOOST_cell_68347 ( .a(TIMEBOOST_net_21381), .b(g65806_sb), .o(n_1589) );
na02f01 TIMEBOOST_cell_3540 ( .a(g65019_db), .b(n_6935), .o(TIMEBOOST_net_330) );
in01f01 g62680_u0 ( .a(FE_OFN1268_n_4095), .o(g62680_sb) );
na03f02 TIMEBOOST_cell_67047 ( .a(FE_OFN1606_n_13997), .b(TIMEBOOST_net_13748), .c(FE_OFN1599_n_13995), .o(n_14476) );
na03f02 TIMEBOOST_cell_66903 ( .a(FE_OFN1747_n_12004), .b(TIMEBOOST_net_16000), .c(n_11977), .o(n_12612) );
na02f06 TIMEBOOST_cell_2934 ( .a(n_550), .b(n_875), .o(TIMEBOOST_net_27) );
in01f01 g62681_u0 ( .a(FE_OFN1268_n_4095), .o(g62681_sb) );
na02f04 TIMEBOOST_cell_2935 ( .a(TIMEBOOST_net_27), .b(n_2235), .o(n_1382) );
na02m04 TIMEBOOST_cell_2936 ( .a(n_879), .b(n_519), .o(TIMEBOOST_net_28) );
in01f01 g62682_u0 ( .a(FE_OFN1208_n_6356), .o(g62682_sb) );
na03s01 TIMEBOOST_cell_35789 ( .a(g58399_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q), .c(g58399_db), .o(n_9209) );
na02m02 TIMEBOOST_cell_2937 ( .a(TIMEBOOST_net_28), .b(n_1968), .o(n_1353) );
na02f20 TIMEBOOST_cell_2938 ( .a(conf_wb_err_addr_in_953), .b(conf_wb_err_addr_in_950), .o(TIMEBOOST_net_29) );
in01f01 g62683_u0 ( .a(FE_OFN1250_n_4093), .o(g62683_sb) );
na03f02 TIMEBOOST_cell_72797 ( .a(TIMEBOOST_net_21609), .b(g64362_sb), .c(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_22457) );
na02f40 TIMEBOOST_cell_2939 ( .a(TIMEBOOST_net_29), .b(n_521), .o(n_1639) );
na02f01 TIMEBOOST_cell_39627 ( .a(TIMEBOOST_net_11425), .b(g62841_sb), .o(n_5290) );
in01f01 g62684_u0 ( .a(FE_OFN1264_n_4095), .o(g62684_sb) );
na02f03 TIMEBOOST_cell_2941 ( .a(TIMEBOOST_net_30), .b(n_1187), .o(n_2009) );
in01m02 g62685_u0 ( .a(FE_OFN1269_n_4095), .o(g62685_sb) );
na02m02 TIMEBOOST_cell_68895 ( .a(TIMEBOOST_net_21655), .b(g64758_db), .o(TIMEBOOST_net_17547) );
na02m04 TIMEBOOST_cell_2943 ( .a(TIMEBOOST_net_31), .b(n_1186), .o(n_2007) );
na03s02 TIMEBOOST_cell_72969 ( .a(n_1915), .b(g61783_sb), .c(g61783_db), .o(n_8239) );
oa12f04 g62686_u0 ( .a(n_2955), .b(n_2954), .c(wbu_addr_in_273), .o(n_3332) );
oa12f02 g62687_u0 ( .a(n_3148), .b(n_3147), .c(wbu_addr_in_276), .o(n_3465) );
in01f02 g62688_u0 ( .a(FE_OFN1231_n_6391), .o(g62688_sb) );
na02f02 TIMEBOOST_cell_40305 ( .a(TIMEBOOST_net_11764), .b(g54175_da), .o(g53935_db) );
na03f02 TIMEBOOST_cell_73339 ( .a(TIMEBOOST_net_13135), .b(n_7618), .c(g59806_sb), .o(n_7617) );
in01f01 g62689_u0 ( .a(FE_OFN1243_n_4092), .o(g62689_sb) );
na02m02 TIMEBOOST_cell_69027 ( .a(TIMEBOOST_net_21721), .b(FE_OFN640_n_4669), .o(TIMEBOOST_net_16265) );
na02f02 TIMEBOOST_cell_2945 ( .a(TIMEBOOST_net_32), .b(n_1186), .o(n_1426) );
na04m02 TIMEBOOST_cell_64658 ( .a(n_3741), .b(g64776_sb), .c(g64776_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q), .o(TIMEBOOST_net_17075) );
in01f01 g62690_u0 ( .a(FE_OFN1243_n_4092), .o(g62690_sb) );
na03m02 TIMEBOOST_cell_72799 ( .a(n_4442), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q), .c(TIMEBOOST_net_12542), .o(TIMEBOOST_net_20968) );
na02f01 TIMEBOOST_cell_70749 ( .a(TIMEBOOST_net_22582), .b(TIMEBOOST_net_16994), .o(n_5513) );
na04f08 TIMEBOOST_cell_73244 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .c(pci_target_unit_pcit_if_strd_addr_in_708), .d(g52637_sb), .o(TIMEBOOST_net_7473) );
in01m01 g62691_u0 ( .a(FE_OFN1241_n_4092), .o(g62691_sb) );
na02m10 TIMEBOOST_cell_53049 ( .a(configuration_pci_err_data_517), .b(wbm_dat_o_16_), .o(TIMEBOOST_net_16742) );
na02f02 TIMEBOOST_cell_3244 ( .a(n_1269), .b(n_3007), .o(TIMEBOOST_net_182) );
oa12s01 g62692_u0 ( .a(pci_target_unit_pcit_if_comp_flush_in), .b(FE_OFN781_n_2746), .c(n_15397), .o(n_4667) );
in01f02 g62693_u0 ( .a(FE_OFN1270_n_4095), .o(g62693_sb) );
na02s01 TIMEBOOST_cell_3175 ( .a(TIMEBOOST_net_147), .b(g65850_sb), .o(n_1585) );
na02m02 TIMEBOOST_cell_49210 ( .a(TIMEBOOST_net_14822), .b(g65815_db), .o(n_1901) );
in01s01 g62695_u0 ( .a(n_15788), .o(n_4666) );
in01f02 g62697_u0 ( .a(FE_OFN1232_n_6391), .o(g62697_sb) );
na02s01 TIMEBOOST_cell_28003 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q), .o(TIMEBOOST_net_8106) );
na02f10 TIMEBOOST_cell_3543 ( .a(TIMEBOOST_net_331), .b(n_3379), .o(n_7618) );
na02s01 TIMEBOOST_cell_48579 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q), .o(TIMEBOOST_net_14507) );
in01m01 g62698_u0 ( .a(FE_OFN1270_n_4095), .o(g62698_sb) );
na02m02 TIMEBOOST_cell_68388 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q), .b(n_4677), .o(TIMEBOOST_net_21402) );
na02f40 TIMEBOOST_cell_3213 ( .a(TIMEBOOST_net_166), .b(n_4743), .o(n_7498) );
na02f02 TIMEBOOST_cell_71010 ( .a(TIMEBOOST_net_17031), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_22713) );
no02f04 g62699_u0 ( .a(conf_wb_err_addr_in_965), .b(n_2429), .o(g62699_p) );
ao12f02 g62699_u1 ( .a(g62699_p), .b(conf_wb_err_addr_in_965), .c(n_2429), .o(n_3154) );
oa12f02 g62700_u0 ( .a(n_3325), .b(n_3324), .c(wbm_adr_o_27_), .o(n_4160) );
in01f02 g62701_u0 ( .a(FE_OFN1234_n_6391), .o(g62701_sb) );
na02m06 TIMEBOOST_cell_45319 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q), .o(TIMEBOOST_net_13554) );
na03m02 TIMEBOOST_cell_70366 ( .a(FE_OFN2021_n_4778), .b(TIMEBOOST_net_16647), .c(TIMEBOOST_net_634), .o(TIMEBOOST_net_22391) );
oa12f02 g62702_u0 ( .a(n_3446), .b(n_1098), .c(n_4662), .o(n_4664) );
oa12f02 g62703_u0 ( .a(n_3444), .b(n_1658), .c(n_4662), .o(n_4663) );
oa12f02 g62704_u0 ( .a(n_3445), .b(n_1688), .c(n_4662), .o(n_4661) );
oa12f02 g62705_u0 ( .a(n_3443), .b(n_2262), .c(n_4662), .o(n_4660) );
in01f01 g62706_u0 ( .a(FE_OFN1268_n_4095), .o(g62706_sb) );
na02s02 TIMEBOOST_cell_30759 ( .a(n_9099), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q), .o(TIMEBOOST_net_9484) );
na02s01 TIMEBOOST_cell_2948 ( .a(n_261), .b(wbu_addr_in_277), .o(TIMEBOOST_net_34) );
in01f02 g62707_u0 ( .a(FE_OFN1250_n_4093), .o(g62707_sb) );
na03f02 TIMEBOOST_cell_66905 ( .a(FE_OFN1748_n_12004), .b(n_12010), .c(TIMEBOOST_net_13549), .o(n_12669) );
na02s01 TIMEBOOST_cell_2949 ( .a(TIMEBOOST_net_34), .b(n_1285), .o(n_1286) );
na02s06 TIMEBOOST_cell_2950 ( .a(pci_target_unit_del_sync_comp_cycle_count_7_), .b(pci_target_unit_del_sync_comp_cycle_count_8_), .o(TIMEBOOST_net_35) );
oa12f02 g62708_u0 ( .a(n_2019), .b(n_2018), .c(pci_target_unit_wishbone_master_rty_counter_7_), .o(n_2451) );
oa12f02 g62709_u0 ( .a(n_2949), .b(n_2948), .c(wbm_adr_o_24_), .o(n_3331) );
in01f01 g62710_u0 ( .a(FE_OFN1244_n_4092), .o(g62710_sb) );
na03s01 TIMEBOOST_cell_72411 ( .a(wbs_dat_i_8_), .b(g61885_sb), .c(TIMEBOOST_net_9648), .o(TIMEBOOST_net_12837) );
na02m04 TIMEBOOST_cell_2951 ( .a(TIMEBOOST_net_35), .b(n_1690), .o(n_878) );
in01s01 TIMEBOOST_cell_45980 ( .a(TIMEBOOST_net_13941), .o(TIMEBOOST_net_13940) );
in01f02 g62711_u0 ( .a(FE_OFN1241_n_4092), .o(g62711_sb) );
na03f02 TIMEBOOST_cell_73697 ( .a(TIMEBOOST_net_13510), .b(n_12004), .c(n_12010), .o(n_12652) );
in01s01 TIMEBOOST_cell_45981 ( .a(conf_wb_err_addr_in_949), .o(TIMEBOOST_net_13942) );
na02f01 TIMEBOOST_cell_2954 ( .a(n_2629), .b(n_2311), .o(TIMEBOOST_net_37) );
in01f02 g62712_u0 ( .a(FE_OFN1206_n_6356), .o(g62712_sb) );
na02f01 TIMEBOOST_cell_2955 ( .a(TIMEBOOST_net_37), .b(n_15407), .o(n_2616) );
in01f02 g62713_u0 ( .a(FE_OFN1246_n_4093), .o(g62713_sb) );
na02f02 TIMEBOOST_cell_52502 ( .a(TIMEBOOST_net_16468), .b(g61867_sb), .o(n_8102) );
in01f02 g62714_u0 ( .a(FE_OFN1288_n_4098), .o(g62714_sb) );
na02s01 TIMEBOOST_cell_38628 ( .a(n_3749), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q), .o(TIMEBOOST_net_10926) );
na02m02 g52461_u1 ( .a(wbs_adr_i_14_), .b(g52461_sb), .o(g52461_da) );
in01f02 g62715_u0 ( .a(FE_OFN1207_n_6356), .o(g62715_sb) );
na02f06 TIMEBOOST_cell_2961 ( .a(TIMEBOOST_net_40), .b(n_1437), .o(n_2018) );
na02f01 TIMEBOOST_cell_2962 ( .a(pci_target_unit_wishbone_master_rty_counter_5_), .b(pci_target_unit_wishbone_master_rty_counter_4_), .o(TIMEBOOST_net_41) );
in01f01 g62716_u0 ( .a(n_4662), .o(g62716_sb) );
in01s01 TIMEBOOST_cell_45886 ( .a(TIMEBOOST_net_13846), .o(TIMEBOOST_net_13847) );
na03s02 TIMEBOOST_cell_65873 ( .a(n_1879), .b(TIMEBOOST_net_21055), .c(g61909_sb), .o(n_8003) );
na02s01 TIMEBOOST_cell_30977 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_13__Q), .b(FE_OFN211_n_9858), .o(TIMEBOOST_net_9593) );
ao12f02 g62717_u0 ( .a(n_3326), .b(conf_wb_err_addr_in_945), .c(FE_OFN1142_n_15261), .o(n_4158) );
ao12f02 g62718_u0 ( .a(n_3323), .b(conf_wb_err_addr_in_948), .c(FE_OFN1142_n_15261), .o(n_4157) );
in01f01 g62719_u0 ( .a(FE_OFN1192_n_6935), .o(g62719_sb) );
na03f02 TIMEBOOST_cell_73626 ( .a(TIMEBOOST_net_16814), .b(n_16748), .c(g52633_sb), .o(n_14674) );
na03f02 TIMEBOOST_cell_65922 ( .a(TIMEBOOST_net_20444), .b(FE_OFN1170_n_5592), .c(g62120_sb), .o(n_5576) );
in01m01 g62720_u0 ( .a(FE_OFN881_g64577_p), .o(g62720_sb) );
na03m02 TIMEBOOST_cell_72521 ( .a(TIMEBOOST_net_21403), .b(g65272_sb), .c(TIMEBOOST_net_21615), .o(TIMEBOOST_net_17028) );
na04f04 TIMEBOOST_cell_73392 ( .a(wbm_dat_o_13_), .b(configuration_pci_err_data_514), .c(FE_OFN1184_n_3476), .d(g60644_sb), .o(n_5684) );
na02s02 TIMEBOOST_cell_49440 ( .a(TIMEBOOST_net_14937), .b(g57988_sb), .o(TIMEBOOST_net_9482) );
in01f01 g62721_u0 ( .a(FE_OFN1130_g64577_p), .o(g62721_sb) );
na02f02 TIMEBOOST_cell_69365 ( .a(TIMEBOOST_net_21890), .b(g60690_sb), .o(TIMEBOOST_net_5476) );
na03f02 TIMEBOOST_cell_67053 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_16542), .c(FE_OFN1600_n_13995), .o(n_16242) );
na02s01 TIMEBOOST_cell_52579 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q), .o(TIMEBOOST_net_16507) );
in01f02 g62722_u0 ( .a(FE_OFN2105_g64577_p), .o(g62722_sb) );
in01m01 TIMEBOOST_cell_64263 ( .a(TIMEBOOST_net_21119), .o(TIMEBOOST_net_21118) );
na02s01 TIMEBOOST_cell_52581 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q), .o(TIMEBOOST_net_16508) );
in01m02 g62723_u0 ( .a(FE_OFN1132_g64577_p), .o(g62723_sb) );
na02s01 TIMEBOOST_cell_52583 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q), .o(TIMEBOOST_net_16509) );
na02m02 TIMEBOOST_cell_68755 ( .a(TIMEBOOST_net_21585), .b(g65012_sb), .o(TIMEBOOST_net_12508) );
na02f02 TIMEBOOST_cell_54271 ( .a(n_4399), .b(g62607_sb), .o(TIMEBOOST_net_17353) );
na02f01 g62724_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q), .b(FE_OFN1106_g64577_p), .o(g62724_db) );
in01f02 g62725_u0 ( .a(FE_OFN2106_g64577_p), .o(g62725_sb) );
na04f04 TIMEBOOST_cell_42512 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_778), .c(FE_OFN2134_n_13124), .d(g54342_sb), .o(n_12972) );
na02s01 TIMEBOOST_cell_38410 ( .a(FE_OFN221_n_9846), .b(g58020_sb), .o(TIMEBOOST_net_10817) );
in01f02 g62726_u0 ( .a(FE_OFN877_g64577_p), .o(g62726_sb) );
na03f02 TIMEBOOST_cell_34812 ( .a(TIMEBOOST_net_9411), .b(FE_OFN1383_n_8567), .c(g57122_sb), .o(n_11624) );
na03f02 TIMEBOOST_cell_65957 ( .a(TIMEBOOST_net_20437), .b(FE_OFN1171_n_5592), .c(g62139_sb), .o(n_5554) );
na02m02 TIMEBOOST_cell_68708 ( .a(g64883_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q), .o(TIMEBOOST_net_21562) );
in01f01 g62727_u0 ( .a(FE_OFN1118_g64577_p), .o(g62727_sb) );
na02s01 TIMEBOOST_cell_71968 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q), .b(FE_OFN1631_n_9531), .o(TIMEBOOST_net_23192) );
na02f02 TIMEBOOST_cell_71315 ( .a(TIMEBOOST_net_22865), .b(FE_OFN714_n_8140), .o(TIMEBOOST_net_16371) );
in01f01 g62728_u0 ( .a(FE_OFN1129_g64577_p), .o(g62728_sb) );
na04f04 TIMEBOOST_cell_42514 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_790), .c(FE_OFN2136_n_13124), .d(g54355_sb), .o(n_13125) );
na02f01 TIMEBOOST_cell_52925 ( .a(TIMEBOOST_net_13064), .b(FE_OFN1134_g64577_p), .o(TIMEBOOST_net_16680) );
in01m01 g62729_u0 ( .a(FE_OFN1106_g64577_p), .o(g62729_sb) );
na02s01 TIMEBOOST_cell_38412 ( .a(FE_OFN221_n_9846), .b(g57958_sb), .o(TIMEBOOST_net_10818) );
na02s01 TIMEBOOST_cell_52585 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q), .o(TIMEBOOST_net_16510) );
in01m01 g62730_u0 ( .a(FE_OFN1115_g64577_p), .o(g62730_sb) );
na02m02 TIMEBOOST_cell_30477 ( .a(n_9590), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q), .o(TIMEBOOST_net_9343) );
na03m02 TIMEBOOST_cell_46926 ( .a(TIMEBOOST_net_12747), .b(g58301_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q), .o(TIMEBOOST_net_9376) );
in01f01 g62731_u0 ( .a(FE_OFN1120_g64577_p), .o(g62731_sb) );
na03f02 TIMEBOOST_cell_73722 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_16873), .c(FE_OFN1577_n_12028), .o(n_12599) );
na02s01 TIMEBOOST_cell_45571 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q), .o(TIMEBOOST_net_13680) );
in01m02 g62732_u0 ( .a(FE_OFN1118_g64577_p), .o(g62732_sb) );
na02f02 TIMEBOOST_cell_54462 ( .a(TIMEBOOST_net_17448), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_15494) );
na04f04 TIMEBOOST_cell_42516 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_783), .c(FE_OFN2134_n_13124), .d(g54347_sb), .o(n_13095) );
na02s01 TIMEBOOST_cell_45579 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q), .o(TIMEBOOST_net_13684) );
in01f01 g62733_u0 ( .a(FE_OFN1125_g64577_p), .o(g62733_sb) );
na04s03 TIMEBOOST_cell_72912 ( .a(g61918_sb), .b(TIMEBOOST_net_152), .c(g65850_sb), .d(g61935_db), .o(n_7953) );
na02m02 TIMEBOOST_cell_42820 ( .a(TIMEBOOST_net_12304), .b(g58785_sb), .o(n_9839) );
in01m01 g62734_u0 ( .a(FE_OFN881_g64577_p), .o(g62734_sb) );
na02f01 g62734_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN881_g64577_p), .o(g62734_db) );
in01f02 g62735_u0 ( .a(FE_OFN1137_g64577_p), .o(g62735_sb) );
na02s01 TIMEBOOST_cell_45401 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_13595) );
na03f02 TIMEBOOST_cell_34744 ( .a(TIMEBOOST_net_9399), .b(FE_OFN1387_n_8567), .c(g57192_sb), .o(n_11561) );
na04f04 TIMEBOOST_cell_42518 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_791), .c(FE_OFN2136_n_13124), .d(g54356_sb), .o(n_13086) );
in01f01 g62736_u0 ( .a(FE_OFN1132_g64577_p), .o(g62736_sb) );
na02m02 TIMEBOOST_cell_54484 ( .a(TIMEBOOST_net_17459), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_15338) );
na04f04 TIMEBOOST_cell_47198 ( .a(n_2917), .b(n_2860), .c(n_3048), .d(n_2829), .o(n_4169) );
na04f04 TIMEBOOST_cell_42520 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_777), .c(FE_OFN2134_n_13124), .d(g54341_sb), .o(n_12974) );
in01f01 g62737_u0 ( .a(FE_OFN1125_g64577_p), .o(g62737_sb) );
na02m02 TIMEBOOST_cell_63935 ( .a(TIMEBOOST_net_20953), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_15815) );
na04f04 TIMEBOOST_cell_42522 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_785), .c(FE_OFN2134_n_13124), .d(g54350_sb), .o(n_13091) );
in01f02 g62738_u0 ( .a(FE_OFN1097_g64577_p), .o(g62738_sb) );
na04f04 TIMEBOOST_cell_42138 ( .a(configuration_wb_err_data_583), .b(FE_OFN1173_n_5592), .c(parchk_pci_ad_out_in_1180), .d(g62083_sb), .o(n_5626) );
na03m02 TIMEBOOST_cell_68868 ( .a(g65090_sb), .b(n_4442), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q), .o(TIMEBOOST_net_21642) );
na03f02 TIMEBOOST_cell_70618 ( .a(n_3991), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q), .c(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_22517) );
in01f01 g62739_u0 ( .a(FE_OFN1120_g64577_p), .o(g62739_sb) );
na02f10 TIMEBOOST_cell_42720 ( .a(n_235), .b(TIMEBOOST_net_12254), .o(n_5641) );
na03f02 TIMEBOOST_cell_73169 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q), .b(g64235_sb), .c(TIMEBOOST_net_20414), .o(TIMEBOOST_net_13110) );
in01f02 g62740_u0 ( .a(FE_OFN1112_g64577_p), .o(g62740_sb) );
na04f04 TIMEBOOST_cell_42524 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_781), .c(FE_OFN2134_n_13124), .d(g54345_sb), .o(n_12968) );
in01m01 g62741_u0 ( .a(FE_OFN1116_g64577_p), .o(g62741_sb) );
na03f02 TIMEBOOST_cell_68646 ( .a(FE_OFN664_n_4495), .b(g64799_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q), .o(TIMEBOOST_net_21531) );
na02s01 TIMEBOOST_cell_38416 ( .a(FE_OFN213_n_9124), .b(g57951_sb), .o(TIMEBOOST_net_10820) );
na02s02 TIMEBOOST_cell_68292 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q), .b(wbu_addr_in_269), .o(TIMEBOOST_net_21354) );
in01f02 g62742_u0 ( .a(FE_OFN2105_g64577_p), .o(g62742_sb) );
na03m02 TIMEBOOST_cell_68744 ( .a(FE_OFN661_n_4392), .b(g64923_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q), .o(TIMEBOOST_net_21580) );
na03m04 TIMEBOOST_cell_73020 ( .a(TIMEBOOST_net_17256), .b(FE_OFN1036_n_4732), .c(g64267_sb), .o(n_3906) );
na02m10 TIMEBOOST_cell_45581 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q), .o(TIMEBOOST_net_13685) );
in01f02 g62743_u0 ( .a(FE_OFN1119_g64577_p), .o(g62743_sb) );
na03f02 TIMEBOOST_cell_73627 ( .a(TIMEBOOST_net_13447), .b(n_16748), .c(g52644_sb), .o(n_14746) );
na04f04 TIMEBOOST_cell_42526 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_779), .c(FE_OFN2135_n_13124), .d(g54343_sb), .o(n_12970) );
na03f02 TIMEBOOST_cell_72524 ( .a(TIMEBOOST_net_21389), .b(g64191_sb), .c(FE_OFN2105_g64577_p), .o(TIMEBOOST_net_22470) );
in01f02 g62744_u0 ( .a(FE_OFN1127_g64577_p), .o(g62744_sb) );
na02f02 TIMEBOOST_cell_54430 ( .a(TIMEBOOST_net_17432), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_15330) );
na02f02 TIMEBOOST_cell_53080 ( .a(TIMEBOOST_net_16757), .b(g62419_sb), .o(n_6759) );
na02m02 TIMEBOOST_cell_49792 ( .a(TIMEBOOST_net_15113), .b(FE_OFN1691_n_9528), .o(TIMEBOOST_net_12747) );
in01f01 g62745_u0 ( .a(FE_OFN1118_g64577_p), .o(g62745_sb) );
na03f02 TIMEBOOST_cell_67998 ( .a(TIMEBOOST_net_21032), .b(FE_OFN1293_n_4098), .c(g62449_sb), .o(n_6699) );
in01f01 g62746_u0 ( .a(FE_OFN1094_g64577_p), .o(g62746_sb) );
na03m02 TIMEBOOST_cell_72858 ( .a(g65405_sb), .b(TIMEBOOST_net_16623), .c(TIMEBOOST_net_16922), .o(TIMEBOOST_net_13246) );
na02m10 TIMEBOOST_cell_52587 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q), .o(TIMEBOOST_net_16511) );
in01f02 g62747_u0 ( .a(FE_OFN1139_g64577_p), .o(g62747_sb) );
na02m01 TIMEBOOST_cell_69260 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q), .b(n_4470), .o(TIMEBOOST_net_21838) );
na03f02 TIMEBOOST_cell_34745 ( .a(TIMEBOOST_net_9562), .b(FE_OFN1370_n_8567), .c(g57401_sb), .o(n_11342) );
in01f02 g62748_u0 ( .a(FE_OFN1139_g64577_p), .o(g62748_sb) );
na02s02 TIMEBOOST_cell_71857 ( .a(TIMEBOOST_net_23136), .b(g65778_sb), .o(n_1600) );
na04f04 TIMEBOOST_cell_73315 ( .a(n_3976), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q), .c(FE_OFN1135_g64577_p), .d(g62839_sb), .o(n_5296) );
in01f01 g62749_u0 ( .a(FE_OFN1125_g64577_p), .o(g62749_sb) );
na02f02 TIMEBOOST_cell_44302 ( .a(TIMEBOOST_net_13045), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_11399) );
in01f06 g62750_u0 ( .a(FE_OFN1133_g64577_p), .o(g62750_sb) );
na03m02 TIMEBOOST_cell_73170 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q), .b(g64283_sb), .c(g64283_db), .o(n_3890) );
na04f04 TIMEBOOST_cell_73139 ( .a(pci_target_unit_fifos_pciw_addr_data_in_151), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q), .c(FE_OFN1077_n_4740), .d(g64082_sb), .o(n_4073) );
in01s01 TIMEBOOST_cell_73917 ( .a(TIMEBOOST_net_23481), .o(TIMEBOOST_net_23482) );
in01f04 g62751_u0 ( .a(FE_OFN1124_g64577_p), .o(g62751_sb) );
na02m02 TIMEBOOST_cell_68709 ( .a(TIMEBOOST_net_21562), .b(TIMEBOOST_net_10506), .o(TIMEBOOST_net_17114) );
na02f02 TIMEBOOST_cell_26206 ( .a(TIMEBOOST_net_7207), .b(FE_OFN1144_n_15261), .o(TIMEBOOST_net_660) );
na04m02 TIMEBOOST_cell_72827 ( .a(n_4473), .b(g64968_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q), .d(TIMEBOOST_net_10587), .o(TIMEBOOST_net_16789) );
in01m01 g62752_u0 ( .a(FE_OFN1120_g64577_p), .o(g62752_sb) );
na03f04 TIMEBOOST_cell_73393 ( .a(TIMEBOOST_net_8387), .b(FE_OFN1182_n_3476), .c(g60629_sb), .o(n_5708) );
na02m08 TIMEBOOST_cell_69550 ( .a(g64946_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q), .o(TIMEBOOST_net_21983) );
na03m02 TIMEBOOST_cell_68966 ( .a(n_3777), .b(g65079_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q), .o(TIMEBOOST_net_21691) );
in01f02 g62753_u0 ( .a(FE_OFN1119_g64577_p), .o(g62753_sb) );
na02s01 TIMEBOOST_cell_47952 ( .a(TIMEBOOST_net_14193), .b(FE_OFN950_n_2055), .o(TIMEBOOST_net_12497) );
na02m01 TIMEBOOST_cell_37404 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q), .b(n_4677), .o(TIMEBOOST_net_10314) );
na03m02 TIMEBOOST_cell_72499 ( .a(TIMEBOOST_net_23132), .b(FE_OFN672_n_4505), .c(g65668_sb), .o(n_1960) );
in01f02 g62754_u0 ( .a(FE_OFN1265_n_4095), .o(g62754_sb) );
na02m04 TIMEBOOST_cell_2963 ( .a(TIMEBOOST_net_41), .b(n_907), .o(n_2001) );
na03f02 TIMEBOOST_cell_66962 ( .a(FE_OCPN1866_n_12377), .b(FE_OFN1756_n_12681), .c(TIMEBOOST_net_13666), .o(n_12673) );
in01f02 g62755_u0 ( .a(FE_OFN1233_n_6391), .o(g62755_sb) );
na02f01 TIMEBOOST_cell_69364 ( .a(wbu_latency_tim_val_in), .b(n_6986), .o(TIMEBOOST_net_21890) );
in01m02 TIMEBOOST_cell_63585 ( .a(TIMEBOOST_net_20764), .o(TIMEBOOST_net_20765) );
na02s02 TIMEBOOST_cell_48580 ( .a(TIMEBOOST_net_14507), .b(FE_OFN1689_n_9528), .o(TIMEBOOST_net_11081) );
in01f01 g62756_u0 ( .a(FE_OFN1128_g64577_p), .o(g62756_sb) );
na02s01 TIMEBOOST_cell_47615 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_75), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_14025) );
in01s01 g62757_u0 ( .a(FE_OFN1092_g64577_p), .o(g62757_sb) );
na04f04 TIMEBOOST_cell_73316 ( .a(n_3875), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q), .c(FE_OFN1119_g64577_p), .d(g63093_sb), .o(n_5066) );
na02f01 TIMEBOOST_cell_70962 ( .a(TIMEBOOST_net_20587), .b(FE_OFN1208_n_6356), .o(TIMEBOOST_net_22689) );
in01f02 g62758_u0 ( .a(FE_OFN1320_n_6436), .o(g62758_sb) );
na02f02 TIMEBOOST_cell_70309 ( .a(TIMEBOOST_net_22362), .b(TIMEBOOST_net_350), .o(n_13664) );
na03f02 TIMEBOOST_cell_73340 ( .a(TIMEBOOST_net_13136), .b(n_7618), .c(g59807_sb), .o(n_7616) );
na02f01 TIMEBOOST_cell_69812 ( .a(FE_OFN1810_n_4454), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q), .o(TIMEBOOST_net_22114) );
in01m01 g62759_u0 ( .a(FE_OFN1116_g64577_p), .o(g62759_sb) );
na02s01 TIMEBOOST_cell_70871 ( .a(TIMEBOOST_net_22643), .b(FE_OFN1657_n_9502), .o(TIMEBOOST_net_16812) );
in01f01 g62760_u0 ( .a(FE_OFN1252_n_4143), .o(g62760_sb) );
na02s02 TIMEBOOST_cell_48846 ( .a(TIMEBOOST_net_14640), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_9508) );
na02f04 TIMEBOOST_cell_2966 ( .a(n_1998), .b(n_2215), .o(TIMEBOOST_net_43) );
in01f01 g62761_u0 ( .a(FE_OFN1265_n_4095), .o(g62761_sb) );
na02s02 TIMEBOOST_cell_25975 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q), .b(FE_OFN952_n_2055), .o(TIMEBOOST_net_7092) );
na02f04 TIMEBOOST_cell_2967 ( .a(TIMEBOOST_net_43), .b(n_2214), .o(n_2701) );
na02m01 TIMEBOOST_cell_2968 ( .a(n_561), .b(n_1416), .o(TIMEBOOST_net_44) );
in01f01 g62762_u0 ( .a(FE_OFN1121_g64577_p), .o(g62762_sb) );
na02m01 TIMEBOOST_cell_62666 ( .a(FE_OFN681_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q), .o(TIMEBOOST_net_20280) );
in01f02 g62763_u0 ( .a(n_6554), .o(g62763_sb) );
na03f02 TIMEBOOST_cell_73806 ( .a(TIMEBOOST_net_13785), .b(FE_OFN1775_n_13800), .c(FE_OFN1769_n_14054), .o(n_14445) );
na02m02 TIMEBOOST_cell_48852 ( .a(TIMEBOOST_net_14643), .b(g58069_sb), .o(TIMEBOOST_net_10855) );
na02f02 TIMEBOOST_cell_44582 ( .a(TIMEBOOST_net_13185), .b(g63012_sb), .o(n_5225) );
in01f01 g62764_u0 ( .a(FE_OFN1130_g64577_p), .o(g62764_sb) );
na04f04 TIMEBOOST_cell_20964 ( .a(FE_RN_613_0), .b(FE_RN_615_0), .c(FE_RN_618_0), .d(FE_RN_611_0), .o(FE_RN_619_0) );
na02m01 TIMEBOOST_cell_48073 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_128), .o(TIMEBOOST_net_14254) );
in01s01 TIMEBOOST_cell_73893 ( .a(TIMEBOOST_net_23457), .o(TIMEBOOST_net_23458) );
in01f01 g62765_u0 ( .a(FE_OFN1132_g64577_p), .o(g62765_sb) );
na03m04 TIMEBOOST_cell_72651 ( .a(TIMEBOOST_net_21493), .b(g64908_sb), .c(TIMEBOOST_net_21677), .o(TIMEBOOST_net_17513) );
na02f02 TIMEBOOST_cell_50270 ( .a(TIMEBOOST_net_15352), .b(g62394_sb), .o(n_6809) );
na02m02 TIMEBOOST_cell_68594 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q), .b(g65021_sb), .o(TIMEBOOST_net_21505) );
in01m02 g62766_u0 ( .a(FE_OFN1130_g64577_p), .o(g62766_sb) );
na03f02 TIMEBOOST_cell_34815 ( .a(TIMEBOOST_net_9341), .b(FE_OFN1413_n_8567), .c(g57440_sb), .o(n_10351) );
na03f02 TIMEBOOST_cell_73781 ( .a(n_13993), .b(TIMEBOOST_net_13714), .c(FE_OFN1588_n_13736), .o(n_14285) );
in01f01 g62767_u0 ( .a(FE_OFN1119_g64577_p), .o(g62767_sb) );
na02m10 TIMEBOOST_cell_70746 ( .a(FE_OFN225_n_9122), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q), .o(TIMEBOOST_net_22581) );
na03f02 TIMEBOOST_cell_65034 ( .a(TIMEBOOST_net_10448), .b(g64254_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q), .o(TIMEBOOST_net_17319) );
in01f06 g62768_u0 ( .a(FE_OFN1136_g64577_p), .o(g62768_sb) );
na03m04 TIMEBOOST_cell_72772 ( .a(n_4493), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q), .c(TIMEBOOST_net_12597), .o(TIMEBOOST_net_17054) );
in01f02 g62769_u0 ( .a(FE_OFN1137_g64577_p), .o(g62769_sb) );
na03m02 TIMEBOOST_cell_65523 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q), .b(g65839_sb), .c(g65839_db), .o(n_1880) );
in01f02 g62770_u0 ( .a(FE_OFN1135_g64577_p), .o(g62770_sb) );
na03f02 TIMEBOOST_cell_66738 ( .a(TIMEBOOST_net_16826), .b(FE_OFN1305_n_13124), .c(g54358_sb), .o(n_13084) );
na02m02 TIMEBOOST_cell_64100 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q), .b(n_4918), .o(TIMEBOOST_net_21036) );
in01f01 g62771_u0 ( .a(FE_OFN1131_g64577_p), .o(g62771_sb) );
na03f02 TIMEBOOST_cell_73394 ( .a(TIMEBOOST_net_16728), .b(FE_OFN1184_n_3476), .c(g60652_sb), .o(n_5672) );
in01s01 TIMEBOOST_cell_73982 ( .a(n_14623), .o(TIMEBOOST_net_23547) );
in01f02 g62772_u0 ( .a(FE_OFN1116_g64577_p), .o(g62772_sb) );
na02f01 TIMEBOOST_cell_43914 ( .a(TIMEBOOST_net_12851), .b(FE_OFN2127_n_16497), .o(TIMEBOOST_net_11378) );
na02f02 TIMEBOOST_cell_27998 ( .a(n_13901), .b(TIMEBOOST_net_8103), .o(TIMEBOOST_net_764) );
in01m01 g62773_u0 ( .a(FE_OFN881_g64577_p), .o(g62773_sb) );
na02f01 g62773_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q), .b(FE_OFN881_g64577_p), .o(g62773_db) );
na02m01 TIMEBOOST_cell_52589 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q), .o(TIMEBOOST_net_16512) );
in01m01 g62774_u0 ( .a(FE_OFN1120_g64577_p), .o(g62774_sb) );
na02m01 TIMEBOOST_cell_43915 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q), .o(TIMEBOOST_net_12852) );
na03f06 TIMEBOOST_cell_73075 ( .a(TIMEBOOST_net_22049), .b(FE_OFN2251_n_2101), .c(g54236_sb), .o(TIMEBOOST_net_23315) );
na02m06 TIMEBOOST_cell_51935 ( .a(pci_target_unit_del_sync_bc_in_201), .b(pci_target_unit_pcit_if_strd_bc_in_717), .o(TIMEBOOST_net_16185) );
in01f01 g62775_u0 ( .a(FE_OFN1136_g64577_p), .o(g62775_sb) );
na03f01 TIMEBOOST_cell_64504 ( .a(n_3741), .b(FE_OFN1679_n_4655), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q), .o(TIMEBOOST_net_14604) );
na02s02 TIMEBOOST_cell_48913 ( .a(FE_OFN254_n_9825), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q), .o(TIMEBOOST_net_14674) );
in01f01 g62776_u0 ( .a(FE_OFN1112_g64577_p), .o(g62776_sb) );
na03m02 TIMEBOOST_cell_66094 ( .a(pci_target_unit_wishbone_master_bc_register_reg_1__Q), .b(g52591_sb), .c(TIMEBOOST_net_5512), .o(n_14686) );
na03f02 TIMEBOOST_cell_73829 ( .a(TIMEBOOST_net_13787), .b(n_13903), .c(FE_OFN1596_n_13741), .o(n_14252) );
in01f02 g62777_u0 ( .a(FE_OFN1106_g64577_p), .o(g62777_sb) );
na02m02 TIMEBOOST_cell_69608 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q), .o(TIMEBOOST_net_22012) );
na02f02 g62777_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q), .b(FE_OFN1106_g64577_p), .o(g62777_db) );
na02s01 TIMEBOOST_cell_69607 ( .a(TIMEBOOST_net_22011), .b(FE_OFN1800_n_9690), .o(TIMEBOOST_net_16948) );
in01m01 g62778_u0 ( .a(FE_OFN882_g64577_p), .o(g62778_sb) );
na02s03 TIMEBOOST_cell_43101 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q), .o(TIMEBOOST_net_12445) );
na03m02 TIMEBOOST_cell_65110 ( .a(n_3777), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q), .c(FE_OFN671_n_4505), .o(TIMEBOOST_net_14464) );
in01m01 g62779_u0 ( .a(FE_OFN1115_g64577_p), .o(g62779_sb) );
na02f01 TIMEBOOST_cell_51318 ( .a(TIMEBOOST_net_15876), .b(FE_OFN1100_g64577_p), .o(TIMEBOOST_net_11369) );
na02m02 TIMEBOOST_cell_69414 ( .a(g64941_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q), .o(TIMEBOOST_net_21915) );
in01f01 g62780_u0 ( .a(FE_OFN1100_g64577_p), .o(g62780_sb) );
na02s01 TIMEBOOST_cell_52591 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q), .o(TIMEBOOST_net_16513) );
in01f01 g62781_u0 ( .a(FE_OFN1123_g64577_p), .o(g62781_sb) );
na03m04 TIMEBOOST_cell_73021 ( .a(FE_OFN1031_n_4732), .b(TIMEBOOST_net_17257), .c(g64300_sb), .o(n_3875) );
na03f02 TIMEBOOST_cell_72984 ( .a(TIMEBOOST_net_16308), .b(FE_OFN948_n_2248), .c(g65914_sb), .o(n_1568) );
in01f01 g62782_u0 ( .a(FE_OFN1130_g64577_p), .o(g62782_sb) );
na02s01 TIMEBOOST_cell_47935 ( .a(FE_OFN527_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q), .o(TIMEBOOST_net_14185) );
na02f01 TIMEBOOST_cell_49389 ( .a(TIMEBOOST_net_8316), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q), .o(TIMEBOOST_net_14912) );
na02f02 TIMEBOOST_cell_69029 ( .a(TIMEBOOST_net_21722), .b(g65094_sb), .o(TIMEBOOST_net_15243) );
in01s01 g62783_u0 ( .a(FE_OFN1097_g64577_p), .o(g62783_sb) );
na02f02 TIMEBOOST_cell_64052 ( .a(n_14618), .b(FE_OFN1189_n_5742), .o(TIMEBOOST_net_21012) );
na02m01 g62783_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q), .b(FE_OFN1097_g64577_p), .o(g62783_db) );
na02m10 TIMEBOOST_cell_52593 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q), .o(TIMEBOOST_net_16514) );
in01f01 g62784_u0 ( .a(FE_OFN1124_g64577_p), .o(g62784_sb) );
na03s01 TIMEBOOST_cell_41921 ( .a(g58349_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q), .c(g58349_db), .o(n_9472) );
in01s01 TIMEBOOST_cell_73970 ( .a(wbm_dat_i_5_), .o(TIMEBOOST_net_23535) );
na02s01 TIMEBOOST_cell_38498 ( .a(FE_OFN241_n_9830), .b(g57970_sb), .o(TIMEBOOST_net_10861) );
in01f02 g62785_u0 ( .a(FE_OFN1119_g64577_p), .o(g62785_sb) );
na04f04 TIMEBOOST_cell_73628 ( .a(pci_target_unit_pcit_if_strd_addr_in_700), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64), .c(n_16748), .d(g52629_sb), .o(n_14661) );
na03s02 TIMEBOOST_cell_52423 ( .a(TIMEBOOST_net_12435), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q), .c(FE_OFN574_n_9902), .o(TIMEBOOST_net_16429) );
na03m02 TIMEBOOST_cell_65960 ( .a(n_3830), .b(g63013_sb), .c(g63013_db), .o(n_5223) );
in01f01 g62786_u0 ( .a(FE_OFN1132_g64577_p), .o(g62786_sb) );
na04f08 TIMEBOOST_cell_20982 ( .a(FE_OFN1026_n_16760), .b(FE_RN_882_0), .c(n_16507), .d(FE_RN_836_0), .o(FE_RN_838_0) );
in01s01 TIMEBOOST_cell_45880 ( .a(TIMEBOOST_net_13840), .o(TIMEBOOST_net_13841) );
na02s03 TIMEBOOST_cell_69156 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q), .o(TIMEBOOST_net_21786) );
in01m01 g62787_u0 ( .a(FE_OFN1124_g64577_p), .o(g62787_sb) );
na02s02 TIMEBOOST_cell_52424 ( .a(TIMEBOOST_net_16429), .b(g58072_sb), .o(TIMEBOOST_net_9506) );
in01m01 g62788_u0 ( .a(FE_OFN1121_g64577_p), .o(g62788_sb) );
na03m02 TIMEBOOST_cell_65961 ( .a(n_3912), .b(g63047_sb), .c(g63047_db), .o(n_5158) );
na02s01 TIMEBOOST_cell_45449 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q), .o(TIMEBOOST_net_13619) );
na03s02 TIMEBOOST_cell_33795 ( .a(n_2202), .b(g61710_sb), .c(g61710_db), .o(n_8406) );
in01f01 g62789_u0 ( .a(FE_OFN1094_g64577_p), .o(g62789_sb) );
na02s01 TIMEBOOST_cell_38598 ( .a(g58013_sb), .b(FE_OFN213_n_9124), .o(TIMEBOOST_net_10911) );
na02m10 TIMEBOOST_cell_52595 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q), .o(TIMEBOOST_net_16515) );
in01m01 g62790_u0 ( .a(FE_OFN1123_g64577_p), .o(g62790_sb) );
na02m02 TIMEBOOST_cell_62456 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_144), .o(TIMEBOOST_net_20175) );
in01f02 g62791_u0 ( .a(FE_OFN877_g64577_p), .o(g62791_sb) );
na02s02 TIMEBOOST_cell_39178 ( .a(FE_OFN270_n_9836), .b(g58217_sb), .o(TIMEBOOST_net_11201) );
na02s01 TIMEBOOST_cell_28867 ( .a(n_741), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .o(TIMEBOOST_net_8538) );
in01m01 g62792_u0 ( .a(FE_OFN1112_g64577_p), .o(g62792_sb) );
na02f10 TIMEBOOST_cell_62884 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_786), .o(TIMEBOOST_net_20389) );
in01f01 g62793_u0 ( .a(FE_OFN1123_g64577_p), .o(g62793_sb) );
na03f02 TIMEBOOST_cell_72962 ( .a(pci_target_unit_del_sync_addr_in_225), .b(g65228_sb), .c(TIMEBOOST_net_7151), .o(n_2659) );
na03f02 TIMEBOOST_cell_72908 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q), .b(g63567_sb), .c(g63567_db), .o(TIMEBOOST_net_12968) );
in01f01 g62794_u0 ( .a(FE_OFN1112_g64577_p), .o(g62794_sb) );
na03s02 TIMEBOOST_cell_72553 ( .a(g58222_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q), .c(g58222_sb), .o(TIMEBOOST_net_12993) );
na02f02 TIMEBOOST_cell_68959 ( .a(TIMEBOOST_net_21687), .b(TIMEBOOST_net_20322), .o(TIMEBOOST_net_17052) );
in01m01 g62795_u0 ( .a(FE_OFN1130_g64577_p), .o(g62795_sb) );
na02s01 TIMEBOOST_cell_68429 ( .a(TIMEBOOST_net_21422), .b(g58151_db), .o(TIMEBOOST_net_14261) );
in01f01 g62796_u0 ( .a(FE_OFN1136_g64577_p), .o(g62796_sb) );
na02m10 TIMEBOOST_cell_45321 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q), .o(TIMEBOOST_net_13555) );
na03m02 TIMEBOOST_cell_72555 ( .a(TIMEBOOST_net_20209), .b(FE_OFN917_n_4725), .c(g64278_sb), .o(TIMEBOOST_net_13053) );
na03m02 TIMEBOOST_cell_72875 ( .a(TIMEBOOST_net_21750), .b(g65752_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q), .o(TIMEBOOST_net_13089) );
in01f01 g62797_u0 ( .a(FE_OFN1132_g64577_p), .o(g62797_sb) );
na04f02 TIMEBOOST_cell_67233 ( .a(n_4479), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q), .c(g64784_sb), .d(FE_OFN1660_n_4490), .o(n_4480) );
in01s01 TIMEBOOST_cell_63584 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_), .o(TIMEBOOST_net_20764) );
na02f02 TIMEBOOST_cell_28000 ( .a(n_13901), .b(TIMEBOOST_net_8104), .o(TIMEBOOST_net_763) );
na02m10 TIMEBOOST_cell_45775 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q), .o(TIMEBOOST_net_13782) );
na03f02 TIMEBOOST_cell_73245 ( .a(n_3856), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q), .c(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_15182) );
na04f02 TIMEBOOST_cell_67990 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q), .b(n_4913), .c(FE_OFN1274_n_4096), .d(g62544_sb), .o(n_7379) );
in01f01 g62799_u0 ( .a(FE_OFN1100_g64577_p), .o(g62799_sb) );
na02s01 TIMEBOOST_cell_52597 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q), .o(TIMEBOOST_net_16516) );
na02m10 TIMEBOOST_cell_45101 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56), .b(pci_target_unit_pcit_if_strd_addr_in_692), .o(TIMEBOOST_net_13445) );
na02m04 TIMEBOOST_cell_69453 ( .a(TIMEBOOST_net_21934), .b(TIMEBOOST_net_14397), .o(TIMEBOOST_net_13359) );
in01m01 g62800_u0 ( .a(FE_OFN1115_g64577_p), .o(g62800_sb) );
na02m06 TIMEBOOST_cell_71987 ( .a(TIMEBOOST_net_23201), .b(g65306_sb), .o(TIMEBOOST_net_12593) );
na02f02 TIMEBOOST_cell_51661 ( .a(FE_OFN1735_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q), .o(TIMEBOOST_net_16048) );
in01f01 g62801_u0 ( .a(FE_OFN2104_g64577_p), .o(g62801_sb) );
na02s02 TIMEBOOST_cell_47739 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q), .b(g65847_sb), .o(TIMEBOOST_net_14087) );
na02m01 TIMEBOOST_cell_37416 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(g65782_sb), .o(TIMEBOOST_net_10320) );
na02s02 TIMEBOOST_cell_70431 ( .a(TIMEBOOST_net_22423), .b(TIMEBOOST_net_20508), .o(TIMEBOOST_net_14471) );
in01m01 g62802_u0 ( .a(FE_OFN2105_g64577_p), .o(g62802_sb) );
na02f02 TIMEBOOST_cell_69923 ( .a(TIMEBOOST_net_22169), .b(n_16000), .o(TIMEBOOST_net_14908) );
na02m01 TIMEBOOST_cell_42903 ( .a(TIMEBOOST_net_9654), .b(n_4725), .o(TIMEBOOST_net_12346) );
na02s01 TIMEBOOST_cell_68168 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_392), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q), .o(TIMEBOOST_net_21292) );
in01f01 g62803_u0 ( .a(FE_OFN1134_g64577_p), .o(g62803_sb) );
na02f01 TIMEBOOST_cell_62547 ( .a(TIMEBOOST_net_20220), .b(FE_OFN918_n_4725), .o(TIMEBOOST_net_14349) );
na03m02 TIMEBOOST_cell_67911 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q), .b(g65872_sb), .c(TIMEBOOST_net_12903), .o(n_1870) );
na03f02 TIMEBOOST_cell_73514 ( .a(TIMEBOOST_net_13362), .b(n_6645), .c(g62654_sb), .o(n_6235) );
in01f02 g62805_u0 ( .a(FE_OFN1100_g64577_p), .o(g62805_sb) );
na02f02 TIMEBOOST_cell_63969 ( .a(TIMEBOOST_net_20970), .b(FE_OFN1214_n_4151), .o(TIMEBOOST_net_15863) );
in01m01 g62806_u0 ( .a(FE_OFN1122_g64577_p), .o(g62806_sb) );
na02f02 TIMEBOOST_cell_70680 ( .a(TIMEBOOST_net_20466), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_22548) );
in01s01 TIMEBOOST_cell_72358 ( .a(pci_target_unit_fifos_pcir_data_in_159), .o(TIMEBOOST_net_23391) );
na03f02 TIMEBOOST_cell_72840 ( .a(g65883_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q), .c(TIMEBOOST_net_14442), .o(TIMEBOOST_net_17013) );
in01f01 g62807_u0 ( .a(FE_OFN1100_g64577_p), .o(g62807_sb) );
na02m02 TIMEBOOST_cell_69724 ( .a(FE_OFN1680_n_4655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q), .o(TIMEBOOST_net_22070) );
na02m08 TIMEBOOST_cell_52733 ( .a(pci_target_unit_pcit_if_strd_addr_in_689), .b(n_2526), .o(TIMEBOOST_net_16584) );
na02f02 TIMEBOOST_cell_69719 ( .a(TIMEBOOST_net_22067), .b(g65347_sb), .o(TIMEBOOST_net_10801) );
in01f01 g62808_u0 ( .a(FE_OFN1106_g64577_p), .o(g62808_sb) );
na02f02 TIMEBOOST_cell_64000 ( .a(wbm_adr_o_11_), .b(g63204_sb), .o(TIMEBOOST_net_20986) );
na02f01 g62808_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q), .b(FE_OFN1106_g64577_p), .o(g62808_db) );
na02m20 TIMEBOOST_cell_52795 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q), .b(pci_target_unit_fifos_pciw_cbe_in_153), .o(TIMEBOOST_net_16615) );
in01f01 g62809_u0 ( .a(FE_OFN2105_g64577_p), .o(g62809_sb) );
in01s01 TIMEBOOST_cell_45881 ( .a(TIMEBOOST_net_13945), .o(TIMEBOOST_net_13842) );
na02s02 TIMEBOOST_cell_39725 ( .a(TIMEBOOST_net_11474), .b(g57906_db), .o(n_9221) );
in01f01 g62810_u0 ( .a(FE_OFN1129_g64577_p), .o(g62810_sb) );
na04m02 TIMEBOOST_cell_67913 ( .a(TIMEBOOST_net_16295), .b(TIMEBOOST_net_12796), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q), .d(FE_OFN702_n_7845), .o(TIMEBOOST_net_14807) );
na02m02 TIMEBOOST_cell_69455 ( .a(TIMEBOOST_net_21935), .b(TIMEBOOST_net_16274), .o(TIMEBOOST_net_17559) );
in01m01 g62811_u0 ( .a(FE_OFN1104_g64577_p), .o(g62811_sb) );
na03f02 TIMEBOOST_cell_66739 ( .a(TIMEBOOST_net_16833), .b(FE_OFN1305_n_13124), .c(g54354_sb), .o(n_13087) );
na03f02 TIMEBOOST_cell_35005 ( .a(TIMEBOOST_net_9573), .b(g57323_sb), .c(FE_OFN2191_n_8567), .o(n_11427) );
in01f01 g62812_u0 ( .a(FE_OFN1112_g64577_p), .o(g62812_sb) );
na03f80 TIMEBOOST_cell_41297 ( .a(n_978), .b(n_16496), .c(n_2887), .o(n_15929) );
na02m02 TIMEBOOST_cell_68279 ( .a(TIMEBOOST_net_21347), .b(TIMEBOOST_net_14165), .o(n_2061) );
in01f02 g62813_u0 ( .a(FE_OFN1135_g64577_p), .o(g62813_sb) );
na02f02 TIMEBOOST_cell_71011 ( .a(TIMEBOOST_net_22713), .b(g63192_sb), .o(n_5772) );
in01s01 TIMEBOOST_cell_73847 ( .a(TIMEBOOST_net_23411), .o(TIMEBOOST_net_23412) );
na02s02 TIMEBOOST_cell_70719 ( .a(TIMEBOOST_net_22567), .b(TIMEBOOST_net_20458), .o(TIMEBOOST_net_17315) );
in01m01 g62814_u0 ( .a(FE_OFN877_g64577_p), .o(g62814_sb) );
na02f01 TIMEBOOST_cell_63947 ( .a(TIMEBOOST_net_20959), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_15692) );
na03f02 TIMEBOOST_cell_73796 ( .a(TIMEBOOST_net_16538), .b(FE_OFN1601_n_13995), .c(FE_OFN1605_n_13997), .o(g53275_p) );
na03f02 TIMEBOOST_cell_65680 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q), .b(g64309_sb), .c(TIMEBOOST_net_14919), .o(TIMEBOOST_net_13078) );
in01m01 g62815_u0 ( .a(FE_OFN882_g64577_p), .o(g62815_sb) );
na03m02 TIMEBOOST_cell_65103 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q), .c(FE_OFN615_n_4501), .o(TIMEBOOST_net_17233) );
na02f01 TIMEBOOST_cell_70192 ( .a(TIMEBOOST_net_12871), .b(FE_OFN2125_n_16497), .o(TIMEBOOST_net_22304) );
in01s01 TIMEBOOST_cell_73918 ( .a(wbm_dat_i_10_), .o(TIMEBOOST_net_23483) );
in01f02 g62816_u0 ( .a(FE_OFN1122_g64577_p), .o(g62816_sb) );
na03f06 TIMEBOOST_cell_65990 ( .a(TIMEBOOST_net_16975), .b(FE_OFN2105_g64577_p), .c(g62842_sb), .o(n_5288) );
na03f02 TIMEBOOST_cell_66209 ( .a(TIMEBOOST_net_20975), .b(FE_OFN1252_n_4143), .c(g62424_sb), .o(n_7387) );
in01f02 g62817_u0 ( .a(FE_OFN2105_g64577_p), .o(g62817_sb) );
na03f02 TIMEBOOST_cell_73782 ( .a(n_13993), .b(TIMEBOOST_net_13718), .c(FE_OFN1588_n_13736), .o(n_14270) );
in01f01 g62818_u0 ( .a(FE_OFN882_g64577_p), .o(g62818_sb) );
na02f02 TIMEBOOST_cell_28002 ( .a(n_13901), .b(TIMEBOOST_net_8105), .o(TIMEBOOST_net_761) );
in01s02 TIMEBOOST_cell_64262 ( .a(TIMEBOOST_net_21118), .o(pci_target_unit_fifos_pcir_data_in_186) );
in01m01 g62819_u0 ( .a(FE_OFN2105_g64577_p), .o(g62819_sb) );
na03f02 TIMEBOOST_cell_67987 ( .a(TIMEBOOST_net_17430), .b(FE_OFN1208_n_6356), .c(g62392_sb), .o(n_6814) );
na02m02 TIMEBOOST_cell_63129 ( .a(TIMEBOOST_net_20511), .b(g58397_db), .o(n_9437) );
in01m02 TIMEBOOST_cell_67738 ( .a(TIMEBOOST_net_21164), .o(TIMEBOOST_net_21165) );
in01f01 g62820_u0 ( .a(FE_OFN1125_g64577_p), .o(g62820_sb) );
na02f02 TIMEBOOST_cell_71013 ( .a(TIMEBOOST_net_22714), .b(g62883_sb), .o(n_6111) );
na02s06 TIMEBOOST_cell_68250 ( .a(n_8884), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q), .o(TIMEBOOST_net_21333) );
in01f02 g62821_u0 ( .a(FE_OFN1097_g64577_p), .o(g62821_sb) );
na02s01 TIMEBOOST_cell_42795 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q), .o(TIMEBOOST_net_12292) );
na03m02 TIMEBOOST_cell_68922 ( .a(g64787_sb), .b(n_4645), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q), .o(TIMEBOOST_net_21669) );
na02s02 TIMEBOOST_cell_42783 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__Q), .b(FE_OFN2054_n_8831), .o(TIMEBOOST_net_12286) );
in01f01 g62822_u0 ( .a(FE_OFN1133_g64577_p), .o(g62822_sb) );
in01s01 TIMEBOOST_cell_63583 ( .a(TIMEBOOST_net_20762), .o(TIMEBOOST_net_20763) );
na03f02 TIMEBOOST_cell_67960 ( .a(n_3957), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q), .c(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_15184) );
in01f01 g62823_u0 ( .a(FE_OFN1112_g64577_p), .o(g62823_sb) );
na02s01 TIMEBOOST_cell_70718 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q), .b(FE_OFN601_n_9687), .o(TIMEBOOST_net_22567) );
in01f02 g62824_u0 ( .a(FE_OFN1116_g64577_p), .o(g62824_sb) );
na02s02 TIMEBOOST_cell_37285 ( .a(TIMEBOOST_net_10254), .b(g65706_sb), .o(n_2200) );
na03f04 TIMEBOOST_cell_66706 ( .a(TIMEBOOST_net_14762), .b(n_8750), .c(n_7543), .o(n_8749) );
na02f02 TIMEBOOST_cell_52276 ( .a(TIMEBOOST_net_16355), .b(g64098_sb), .o(n_4057) );
in01f01 g62825_u0 ( .a(FE_OFN1124_g64577_p), .o(g62825_sb) );
na03f02 TIMEBOOST_cell_73822 ( .a(TIMEBOOST_net_13804), .b(n_13903), .c(FE_OCP_RBN1962_FE_OFN1591_n_13741), .o(n_16250) );
na02f02 TIMEBOOST_cell_68070 ( .a(n_513), .b(n_1285), .o(TIMEBOOST_net_21243) );
na03f02 TIMEBOOST_cell_73662 ( .a(TIMEBOOST_net_20581), .b(FE_OFN1236_n_6391), .c(g62981_sb), .o(n_5920) );
in01f01 g62826_u0 ( .a(FE_OFN2106_g64577_p), .o(g62826_sb) );
na02s01 TIMEBOOST_cell_45103 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79), .b(pci_target_unit_pcit_if_strd_addr_in_715), .o(TIMEBOOST_net_13446) );
na03m02 TIMEBOOST_cell_68610 ( .a(n_3764), .b(g65016_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q), .o(TIMEBOOST_net_21513) );
na02f02 TIMEBOOST_cell_69197 ( .a(TIMEBOOST_net_21806), .b(g64287_sb), .o(n_3886) );
in01f01 g62827_u0 ( .a(FE_OFN1120_g64577_p), .o(g62827_sb) );
na02m01 TIMEBOOST_cell_29257 ( .a(n_7835), .b(n_1117), .o(TIMEBOOST_net_8733) );
na02m08 TIMEBOOST_cell_51937 ( .a(pci_target_unit_pcit_if_strd_bc_in_719), .b(pci_target_unit_del_sync_bc_in_203), .o(TIMEBOOST_net_16186) );
na02m02 TIMEBOOST_cell_68605 ( .a(TIMEBOOST_net_21510), .b(TIMEBOOST_net_10386), .o(TIMEBOOST_net_17023) );
in01f01 g62828_u0 ( .a(FE_OFN2106_g64577_p), .o(g62828_sb) );
na02m04 TIMEBOOST_cell_53241 ( .a(n_9627), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q), .o(TIMEBOOST_net_16838) );
na03f02 TIMEBOOST_cell_72713 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q), .b(g65942_sb), .c(g65942_db), .o(n_1563) );
in01m01 g62829_u0 ( .a(FE_OFN1124_g64577_p), .o(g62829_sb) );
in01f01 g62830_u0 ( .a(FE_OFN1120_g64577_p), .o(g62830_sb) );
na02s01 TIMEBOOST_cell_43743 ( .a(g58057_sb), .b(FE_OFN235_n_9834), .o(TIMEBOOST_net_12766) );
in01s01 TIMEBOOST_cell_46003 ( .a(TIMEBOOST_net_13964), .o(TIMEBOOST_net_13861) );
na02f02 TIMEBOOST_cell_48131 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q), .b(g65854_sb), .o(TIMEBOOST_net_14283) );
in01f02 g62831_u0 ( .a(FE_OFN877_g64577_p), .o(g62831_sb) );
na03f02 TIMEBOOST_cell_34746 ( .a(TIMEBOOST_net_9400), .b(FE_OFN1389_n_8567), .c(g57349_sb), .o(n_11401) );
na03m02 TIMEBOOST_cell_66098 ( .a(pci_target_unit_wishbone_master_bc_register_reg_0__Q), .b(g52590_sb), .c(TIMEBOOST_net_5513), .o(n_14687) );
na02f02 TIMEBOOST_cell_49674 ( .a(TIMEBOOST_net_15054), .b(g62026_sb), .o(n_7844) );
in01f01 g62832_u0 ( .a(FE_OFN1136_g64577_p), .o(g62832_sb) );
na03f02 TIMEBOOST_cell_34748 ( .a(TIMEBOOST_net_9440), .b(FE_OFN1412_n_8567), .c(g57583_sb), .o(n_10291) );
na02m10 TIMEBOOST_cell_53051 ( .a(configuration_pci_err_data_525), .b(wbm_dat_o_24_), .o(TIMEBOOST_net_16743) );
in01f01 g62833_u0 ( .a(FE_OFN1134_g64577_p), .o(g62833_sb) );
na03f02 TIMEBOOST_cell_67989 ( .a(TIMEBOOST_net_13250), .b(FE_OFN1193_n_6935), .c(g62653_sb), .o(n_6238) );
na03s02 TIMEBOOST_cell_41900 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q), .b(g58355_sb), .c(g58355_db), .o(n_9467) );
in01m02 g62834_u0 ( .a(FE_OFN1118_g64577_p), .o(g62834_sb) );
na03f02 TIMEBOOST_cell_73556 ( .a(TIMEBOOST_net_17512), .b(FE_OFN1234_n_6391), .c(g62701_sb), .o(n_6156) );
na02f02 TIMEBOOST_cell_69840 ( .a(n_1906), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q), .o(TIMEBOOST_net_22128) );
in01f02 g62835_u0 ( .a(FE_OFN1106_g64577_p), .o(g62835_sb) );
na02m02 TIMEBOOST_cell_69567 ( .a(TIMEBOOST_net_21991), .b(TIMEBOOST_net_16918), .o(n_1937) );
na02f01 g62835_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN1106_g64577_p), .o(g62835_db) );
na02m08 TIMEBOOST_cell_52599 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q), .o(TIMEBOOST_net_16517) );
in01f01 g62836_u0 ( .a(FE_OFN2105_g64577_p), .o(g62836_sb) );
na03f02 TIMEBOOST_cell_34750 ( .a(TIMEBOOST_net_9335), .b(FE_OFN1400_n_8567), .c(g57549_sb), .o(n_11196) );
na02m02 TIMEBOOST_cell_51454 ( .a(TIMEBOOST_net_15944), .b(g52646_sb), .o(TIMEBOOST_net_5666) );
in01m02 g62837_u0 ( .a(FE_OFN1119_g64577_p), .o(g62837_sb) );
na02s01 TIMEBOOST_cell_29273 ( .a(FE_OFN1651_n_9428), .b(n_8892), .o(TIMEBOOST_net_8741) );
na02f02 TIMEBOOST_cell_45104 ( .a(TIMEBOOST_net_13446), .b(n_16748), .o(TIMEBOOST_net_11886) );
na03m04 TIMEBOOST_cell_72743 ( .a(n_4482), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q), .c(TIMEBOOST_net_12513), .o(TIMEBOOST_net_17508) );
in01m01 g62838_u0 ( .a(FE_OFN1122_g64577_p), .o(g62838_sb) );
na02f01 TIMEBOOST_cell_51467 ( .a(n_2768), .b(n_3593), .o(TIMEBOOST_net_15951) );
na03f02 TIMEBOOST_cell_73246 ( .a(TIMEBOOST_net_23305), .b(g64089_sb), .c(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_22460) );
in01f02 g62839_u0 ( .a(FE_OFN1135_g64577_p), .o(g62839_sb) );
na02m02 TIMEBOOST_cell_68897 ( .a(TIMEBOOST_net_21656), .b(g64933_sb), .o(TIMEBOOST_net_21037) );
na04f04 TIMEBOOST_cell_68018 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_412), .b(g54193_sb), .c(TIMEBOOST_net_7615), .d(FE_OFN1085_n_13221), .o(n_13424) );
na02s02 TIMEBOOST_cell_17969 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q), .b(n_8831), .o(TIMEBOOST_net_5348) );
in01f02 g62840_u0 ( .a(FE_OFN1135_g64577_p), .o(g62840_sb) );
na02f02 TIMEBOOST_cell_49796 ( .a(TIMEBOOST_net_15115), .b(g54139_da), .o(n_13562) );
na03f02 TIMEBOOST_cell_73557 ( .a(TIMEBOOST_net_8877), .b(g54184_sb), .c(g54184_db), .o(n_13359) );
na04m08 TIMEBOOST_cell_72745 ( .a(FE_OFN614_n_4501), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q), .c(n_4479), .d(g64807_sb), .o(TIMEBOOST_net_7584) );
in01m01 g62841_u0 ( .a(FE_OFN1115_g64577_p), .o(g62841_sb) );
na02m02 TIMEBOOST_cell_54274 ( .a(TIMEBOOST_net_17354), .b(g58371_db), .o(TIMEBOOST_net_9545) );
na02s01 TIMEBOOST_cell_48097 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q), .b(pci_target_unit_fifos_pcir_data_in_173), .o(TIMEBOOST_net_14266) );
na03f02 TIMEBOOST_cell_66938 ( .a(FE_OFN1753_n_12086), .b(FE_OFN2210_n_11027), .c(TIMEBOOST_net_13616), .o(n_12711) );
in01f08 g62842_u0 ( .a(FE_OFN2106_g64577_p), .o(g62842_sb) );
na02m02 TIMEBOOST_cell_69536 ( .a(g64859_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q), .o(TIMEBOOST_net_21976) );
in01m01 g62843_u0 ( .a(FE_OFN1104_g64577_p), .o(g62843_sb) );
na02s01 TIMEBOOST_cell_52601 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q), .o(TIMEBOOST_net_16518) );
na02m10 TIMEBOOST_cell_28999 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q), .o(TIMEBOOST_net_8604) );
na03f02 TIMEBOOST_cell_73515 ( .a(TIMEBOOST_net_17054), .b(n_6431), .c(g62939_sb), .o(n_6003) );
in01m01 g62844_u0 ( .a(FE_OFN881_g64577_p), .o(g62844_sb) );
na02m02 TIMEBOOST_cell_68632 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q), .b(FE_OFN679_n_4460), .o(TIMEBOOST_net_21524) );
na02f01 g62844_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q), .b(FE_OFN881_g64577_p), .o(g62844_db) );
na02m02 TIMEBOOST_cell_50019 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q), .b(g58296_sb), .o(TIMEBOOST_net_15227) );
in01f02 g62845_u0 ( .a(FE_OFN1135_g64577_p), .o(g62845_sb) );
na02m02 TIMEBOOST_cell_69231 ( .a(TIMEBOOST_net_21823), .b(n_4470), .o(TIMEBOOST_net_16329) );
na02m02 TIMEBOOST_cell_69630 ( .a(g65298_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q), .o(TIMEBOOST_net_22023) );
na03f02 TIMEBOOST_cell_67991 ( .a(TIMEBOOST_net_13247), .b(FE_OFN1242_n_4092), .c(g62652_sb), .o(n_6240) );
in01f01 g62846_u0 ( .a(FE_OFN1136_g64577_p), .o(g62846_sb) );
na02m06 TIMEBOOST_cell_69246 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_21831) );
na02s01 TIMEBOOST_cell_48101 ( .a(pci_target_unit_pcit_if_strd_addr_in_686), .b(n_2598), .o(TIMEBOOST_net_14268) );
na02m02 g64948_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q), .b(FE_OFN649_n_4497), .o(g64948_db) );
in01m01 g62847_u0 ( .a(FE_OFN1121_g64577_p), .o(g62847_sb) );
no02f10 TIMEBOOST_cell_44073 ( .a(FE_RN_66_0), .b(n_15402), .o(TIMEBOOST_net_12931) );
in01m01 g62848_u0 ( .a(FE_OFN1106_g64577_p), .o(g62848_sb) );
na02f01 g62848_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN1106_g64577_p), .o(g62848_db) );
na02m06 TIMEBOOST_cell_68596 ( .a(FE_OFN631_n_4454), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_21506) );
in01m01 g62849_u0 ( .a(FE_OFN877_g64577_p), .o(g62849_sb) );
na02s02 TIMEBOOST_cell_43655 ( .a(FE_OFN223_n_9844), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q), .o(TIMEBOOST_net_12722) );
na03f02 TIMEBOOST_cell_70012 ( .a(n_1909), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q), .c(FE_OFN714_n_8140), .o(TIMEBOOST_net_22214) );
in01f01 g62850_u0 ( .a(FE_OFN1129_g64577_p), .o(g62850_sb) );
na03f02 TIMEBOOST_cell_66936 ( .a(FE_OFN1753_n_12086), .b(FE_OFN1568_n_11027), .c(TIMEBOOST_net_13618), .o(n_12650) );
na02f02 TIMEBOOST_cell_70311 ( .a(TIMEBOOST_net_22363), .b(g54154_sb), .o(n_13657) );
na03f02 TIMEBOOST_cell_35062 ( .a(TIMEBOOST_net_9600), .b(FE_OFN1439_n_9372), .c(g58476_sb), .o(n_9363) );
in01m01 g62851_u0 ( .a(FE_OFN881_g64577_p), .o(g62851_sb) );
na02f02 TIMEBOOST_cell_49154 ( .a(TIMEBOOST_net_14794), .b(g61770_sb), .o(n_8269) );
na03f02 TIMEBOOST_cell_47334 ( .a(FE_OFN1558_n_12042), .b(TIMEBOOST_net_13625), .c(FE_OFN1574_n_12028), .o(n_12656) );
in01m01 g62852_u0 ( .a(FE_OFN1104_g64577_p), .o(g62852_sb) );
na04f04 TIMEBOOST_cell_67692 ( .a(TIMEBOOST_net_16867), .b(FE_OFN2200_n_10256), .c(g52603_sb), .d(TIMEBOOST_net_696), .o(n_11868) );
na02m10 TIMEBOOST_cell_52789 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_150), .o(TIMEBOOST_net_16612) );
in01f01 g62853_u0 ( .a(FE_OFN1120_g64577_p), .o(g62853_sb) );
na02s01 TIMEBOOST_cell_43065 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q), .o(TIMEBOOST_net_12427) );
na03f02 TIMEBOOST_cell_34871 ( .a(TIMEBOOST_net_9415), .b(FE_OFN1396_n_8567), .c(g57219_sb), .o(n_11536) );
na03s02 TIMEBOOST_cell_63054 ( .a(FE_OFN250_n_9789), .b(FE_OFN593_n_9694), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q), .o(TIMEBOOST_net_20474) );
in01m02 g62854_u0 ( .a(FE_OFN1118_g64577_p), .o(g62854_sb) );
na02m06 TIMEBOOST_cell_68516 ( .a(g65286_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q), .o(TIMEBOOST_net_21466) );
na03m02 TIMEBOOST_cell_73107 ( .a(g64827_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q), .c(TIMEBOOST_net_14682), .o(TIMEBOOST_net_20525) );
in01f02 g62855_u0 ( .a(FE_OFN1112_g64577_p), .o(g62855_sb) );
na02m01 TIMEBOOST_cell_29299 ( .a(n_3747), .b(FE_OFN643_n_4677), .o(TIMEBOOST_net_8754) );
na02m02 TIMEBOOST_cell_69384 ( .a(FE_OFN646_n_4497), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q), .o(TIMEBOOST_net_21900) );
in01f02 g62856_u0 ( .a(FE_OFN1135_g64577_p), .o(g62856_sb) );
na03m04 TIMEBOOST_cell_72841 ( .a(g65305_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q), .c(TIMEBOOST_net_23229), .o(TIMEBOOST_net_17499) );
na02f02 TIMEBOOST_cell_38755 ( .a(TIMEBOOST_net_10989), .b(g65920_db), .o(n_1566) );
na02s02 TIMEBOOST_cell_38500 ( .a(FE_OFN254_n_9825), .b(g58228_sb), .o(TIMEBOOST_net_10862) );
in01f01 g62857_u0 ( .a(FE_OFN1137_g64577_p), .o(g62857_sb) );
na03s02 TIMEBOOST_cell_72533 ( .a(TIMEBOOST_net_21149), .b(g65714_sb), .c(g65714_db), .o(n_1944) );
na02m02 TIMEBOOST_cell_68862 ( .a(n_4498), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q), .o(TIMEBOOST_net_21639) );
na03f02 TIMEBOOST_cell_73395 ( .a(TIMEBOOST_net_16735), .b(FE_OFN1184_n_3476), .c(g60613_sb), .o(n_4841) );
in01s01 g62858_u0 ( .a(FE_OFN1097_g64577_p), .o(g62858_sb) );
na02s01 TIMEBOOST_cell_38422 ( .a(FE_OFN211_n_9858), .b(g57981_sb), .o(TIMEBOOST_net_10823) );
na02m01 g62858_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q), .b(FE_OFN1097_g64577_p), .o(g62858_db) );
na03f06 TIMEBOOST_cell_71440 ( .a(configuration_wb_err_addr_556), .b(n_15444), .c(FE_RN_566_0), .o(TIMEBOOST_net_22928) );
in01f01 g62859_u0 ( .a(FE_OFN1100_g64577_p), .o(g62859_sb) );
na02s02 TIMEBOOST_cell_63128 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q), .b(g58397_sb), .o(TIMEBOOST_net_20511) );
in01f02 g62860_u0 ( .a(FE_OFN2104_g64577_p), .o(g62860_sb) );
na03f02 TIMEBOOST_cell_34743 ( .a(TIMEBOOST_net_9398), .b(FE_OFN1387_n_8567), .c(g57535_sb), .o(n_11207) );
in01f06 g62861_u0 ( .a(FE_OFN2104_g64577_p), .o(g62861_sb) );
na03f02 TIMEBOOST_cell_47376 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_13684), .c(FE_OFN1581_n_12306), .o(n_12490) );
na03f02 TIMEBOOST_cell_73463 ( .a(TIMEBOOST_net_17472), .b(FE_OFN1269_n_4095), .c(g63189_sb), .o(n_5776) );
in01s01 TIMEBOOST_cell_64261 ( .a(TIMEBOOST_net_21117), .o(TIMEBOOST_net_21116) );
in01f01 g62862_u0 ( .a(FE_OFN1136_g64577_p), .o(g62862_sb) );
na02s02 TIMEBOOST_cell_63325 ( .a(TIMEBOOST_net_20609), .b(g58260_sb), .o(TIMEBOOST_net_9573) );
na02s01 g65698_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q), .b(FE_OFN937_n_2292), .o(g65698_db) );
in01f01 g62863_u0 ( .a(FE_OFN1131_g64577_p), .o(g62863_sb) );
na02s02 TIMEBOOST_cell_72162 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q), .b(FE_OFN702_n_7845), .o(TIMEBOOST_net_23289) );
na02m02 TIMEBOOST_cell_54682 ( .a(TIMEBOOST_net_17558), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_15342) );
in01f04 g62864_u0 ( .a(FE_OFN1123_g64577_p), .o(g62864_sb) );
na03s02 TIMEBOOST_cell_41744 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q), .b(g58449_sb), .c(g58449_db), .o(n_9407) );
in01m01 g62865_u0 ( .a(FE_OFN882_g64577_p), .o(g62865_sb) );
na03s01 TIMEBOOST_cell_64501 ( .a(TIMEBOOST_net_14048), .b(g65964_sb), .c(TIMEBOOST_net_20848), .o(n_7911) );
na02f01 TIMEBOOST_cell_54232 ( .a(TIMEBOOST_net_17333), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_15166) );
na03f02 TIMEBOOST_cell_34904 ( .a(TIMEBOOST_net_9449), .b(FE_OFN1391_n_8567), .c(g57572_sb), .o(n_11179) );
na02f01 TIMEBOOST_cell_26105 ( .a(pci_target_unit_pcit_if_strd_addr_in_696), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7157) );
ao22f06 g62868_u0 ( .a(n_4642), .b(n_16160), .c(n_1447), .d(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_17030) );
ao12f02 g62869_u0 ( .a(n_3321), .b(n_16000), .c(n_2833), .o(n_4155) );
ao12f02 g62870_u0 ( .a(n_4136), .b(FE_OFN1066_n_15808), .c(configuration_pci_err_data_504), .o(n_4803) );
ao12f02 g62871_u0 ( .a(n_4135), .b(FE_OFN1066_n_15808), .c(configuration_pci_err_data_506), .o(n_4802) );
oa12f02 g62872_u0 ( .a(n_3327), .b(conf_wb_err_addr_in_943), .c(FE_OFN1142_n_15261), .o(n_4154) );
no02f01 g62873_u0 ( .a(n_1419), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_), .o(g62873_p) );
ao12f01 g62873_u1 ( .a(g62873_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_), .c(n_1419), .o(n_2274) );
no02s01 g62874_u0 ( .a(n_2013), .b(wbu_addr_in_254), .o(g62874_p) );
ao12s01 g62874_u1 ( .a(g62874_p), .b(wbu_addr_in_254), .c(n_2013), .o(n_2273) );
no02f04 g62875_u0 ( .a(conf_wb_err_addr_in_957), .b(n_2436), .o(g62875_p) );
ao12f02 g62875_u1 ( .a(g62875_p), .b(conf_wb_err_addr_in_957), .c(n_2436), .o(n_3153) );
no02f01 g62876_u0 ( .a(conf_wb_err_addr_in_946), .b(n_1463), .o(g62876_p) );
ao12f01 g62876_u1 ( .a(g62876_p), .b(conf_wb_err_addr_in_946), .c(n_1463), .o(n_2272) );
no02s02 g62877_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_3_), .b(n_1190), .o(g62877_p) );
ao12s01 g62877_u1 ( .a(g62877_p), .b(pci_target_unit_del_sync_comp_cycle_count_3_), .c(n_1190), .o(n_2024) );
oa12f02 g62878_u0 ( .a(n_3447), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_), .c(n_4662), .o(n_4659) );
no02f04 g62879_u0 ( .a(n_2012), .b(wbm_adr_o_5_), .o(g62879_p) );
ao12f02 g62879_u1 ( .a(g62879_p), .b(wbm_adr_o_5_), .c(n_2012), .o(n_2271) );
no02m01 g62880_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_3_), .b(n_1213), .o(g62880_p) );
ao12m01 g62880_u1 ( .a(g62880_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_3_), .c(n_1213), .o(n_2023) );
no02f01 g62881_u0 ( .a(n_1216), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_), .o(g62881_p) );
ao12f01 g62881_u1 ( .a(g62881_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_), .c(n_1216), .o(n_2022) );
no02f02 g62882_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(FE_OFN1192_n_6935), .o(g62882_p) );
ao12f02 g62882_u1 ( .a(g62882_p), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .c(FE_OFN1192_n_6935), .o(n_6112) );
in01f01 g62883_u0 ( .a(FE_OFN1202_n_4090), .o(g62883_sb) );
na03f02 TIMEBOOST_cell_66785 ( .a(TIMEBOOST_net_17063), .b(n_6319), .c(g62990_sb), .o(n_5902) );
na02f01 TIMEBOOST_cell_2969 ( .a(TIMEBOOST_net_44), .b(n_1175), .o(n_1417) );
na02m02 TIMEBOOST_cell_44390 ( .a(TIMEBOOST_net_13089), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_11424) );
in01f02 g62884_u0 ( .a(FE_OFN1288_n_4098), .o(g62884_sb) );
na03f02 TIMEBOOST_cell_73247 ( .a(TIMEBOOST_net_22283), .b(g64092_sb), .c(FE_OFN1116_g64577_p), .o(TIMEBOOST_net_22463) );
na03m02 TIMEBOOST_cell_64842 ( .a(TIMEBOOST_net_16902), .b(g64902_sb), .c(TIMEBOOST_net_20336), .o(TIMEBOOST_net_13226) );
in01f02 g62885_u0 ( .a(FE_OFN1310_n_6624), .o(g62885_sb) );
na02f04 TIMEBOOST_cell_71906 ( .a(g63548_db), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q), .o(TIMEBOOST_net_23161) );
na04m04 TIMEBOOST_cell_72544 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(g65764_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q), .d(g65764_db), .o(TIMEBOOST_net_22039) );
na02m01 TIMEBOOST_cell_68172 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_400), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q), .o(TIMEBOOST_net_21294) );
in01m02 g62886_u0 ( .a(FE_OFN1289_n_4098), .o(g62886_sb) );
na02s02 TIMEBOOST_cell_54170 ( .a(TIMEBOOST_net_17302), .b(g58170_sb), .o(TIMEBOOST_net_16400) );
no02f10 TIMEBOOST_cell_2973 ( .a(TIMEBOOST_net_46), .b(n_15999), .o(n_16000) );
no02s02 TIMEBOOST_cell_2974 ( .a(n_382), .b(wbs_adr_i_5_), .o(TIMEBOOST_net_47) );
in01m01 g62887_u0 ( .a(FE_OFN1249_n_4093), .o(g62887_sb) );
na02f01 TIMEBOOST_cell_70630 ( .a(TIMEBOOST_net_13041), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_22523) );
na02s01 TIMEBOOST_cell_47740 ( .a(TIMEBOOST_net_14087), .b(g65847_db), .o(n_1655) );
in01f02 g62888_u0 ( .a(FE_OFN1258_n_4143), .o(g62888_sb) );
no03f02 TIMEBOOST_cell_35109 ( .a(n_15769), .b(n_2416), .c(FE_OFN1506_n_15768), .o(n_11448) );
na02f02 TIMEBOOST_cell_70347 ( .a(TIMEBOOST_net_22381), .b(g63595_sb), .o(n_7161) );
na02f02 TIMEBOOST_cell_51468 ( .a(TIMEBOOST_net_15951), .b(n_3454), .o(TIMEBOOST_net_452) );
in01f02 g62889_u0 ( .a(FE_OFN1253_n_4143), .o(g62889_sb) );
na03f02 TIMEBOOST_cell_33479 ( .a(TIMEBOOST_net_8789), .b(FE_OFN1168_n_5592), .c(g62098_sb), .o(n_5606) );
na03f04 TIMEBOOST_cell_68606 ( .a(n_2078), .b(n_1742), .c(n_2778), .o(TIMEBOOST_net_21511) );
in01f01 g62890_u0 ( .a(FE_OFN1265_n_4095), .o(g62890_sb) );
na03f02 TIMEBOOST_cell_73558 ( .a(TIMEBOOST_net_17509), .b(FE_OFN1234_n_6391), .c(g62646_sb), .o(n_6257) );
na02m02 TIMEBOOST_cell_68452 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q), .b(FE_OFN670_n_4505), .o(TIMEBOOST_net_21434) );
na02f01 TIMEBOOST_cell_2982 ( .a(pci_target_unit_pci_target_if_target_rd_completed), .b(n_12595), .o(TIMEBOOST_net_51) );
in01f01 g62891_u0 ( .a(FE_OFN1272_n_4096), .o(g62891_sb) );
na02f02 TIMEBOOST_cell_2983 ( .a(TIMEBOOST_net_51), .b(n_2287), .o(n_2746) );
na02f02 TIMEBOOST_cell_54470 ( .a(TIMEBOOST_net_17452), .b(FE_OFN1214_n_4151), .o(TIMEBOOST_net_15869) );
in01m01 g62892_u0 ( .a(FE_OFN1219_n_6886), .o(g62892_sb) );
na02f01 TIMEBOOST_cell_27219 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_7714) );
na02f01 TIMEBOOST_cell_49704 ( .a(TIMEBOOST_net_15069), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_13439) );
na03f02 TIMEBOOST_cell_73248 ( .a(TIMEBOOST_net_23307), .b(g54326_sb), .c(g54040_sb), .o(TIMEBOOST_net_22888) );
in01f01 g62893_u0 ( .a(FE_OFN1248_n_4093), .o(g62893_sb) );
na02m02 TIMEBOOST_cell_54294 ( .a(TIMEBOOST_net_17364), .b(FE_OFN1203_n_4090), .o(TIMEBOOST_net_15419) );
na02f02 TIMEBOOST_cell_71479 ( .a(TIMEBOOST_net_22947), .b(TIMEBOOST_net_16007), .o(n_14815) );
na03f02 TIMEBOOST_cell_41993 ( .a(TIMEBOOST_net_10976), .b(g64204_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q), .o(TIMEBOOST_net_9309) );
in01f02 g62894_u0 ( .a(FE_OFN1202_n_4090), .o(g62894_sb) );
na02m02 TIMEBOOST_cell_43703 ( .a(FE_OFN1807_n_4501), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q), .o(TIMEBOOST_net_12746) );
in01f02 g62895_u0 ( .a(FE_OFN1260_n_4143), .o(g62895_sb) );
na04f02 TIMEBOOST_cell_25260 ( .a(n_14454), .b(n_13972), .c(n_14556), .d(n_13857), .o(n_14601) );
in01s01 TIMEBOOST_cell_73919 ( .a(TIMEBOOST_net_23483), .o(TIMEBOOST_net_23484) );
in01f01 g62896_u0 ( .a(FE_OFN1284_n_4097), .o(g62896_sb) );
na04f02 TIMEBOOST_cell_25261 ( .a(n_16244), .b(n_14000), .c(n_13999), .d(n_16241), .o(n_16247) );
na03m02 TIMEBOOST_cell_71970 ( .a(n_4470), .b(g64962_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q), .o(TIMEBOOST_net_23193) );
na02f04 TIMEBOOST_cell_39763 ( .a(TIMEBOOST_net_11493), .b(g54152_sb), .o(n_13448) );
in01m02 g62897_u0 ( .a(FE_OFN1294_n_4098), .o(g62897_sb) );
na02m02 TIMEBOOST_cell_43563 ( .a(pci_target_unit_fifos_pciw_addr_data_in_147), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_12676) );
na03f02 TIMEBOOST_cell_66377 ( .a(TIMEBOOST_net_17066), .b(FE_OFN1225_n_6391), .c(g62460_sb), .o(n_6676) );
na03m02 TIMEBOOST_cell_72846 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q), .b(g65330_sb), .c(TIMEBOOST_net_22016), .o(TIMEBOOST_net_17425) );
in01f02 g62898_u0 ( .a(FE_OFN1310_n_6624), .o(g62898_sb) );
na04f02 TIMEBOOST_cell_35121 ( .a(wbs_dat_o_15_), .b(g52509_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_114), .d(FE_OFN1472_g52675_p), .o(n_13744) );
na02f02 TIMEBOOST_cell_3833 ( .a(FE_RN_26_0), .b(TIMEBOOST_net_476), .o(n_12817) );
na02m02 g54194_u2 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_30__Q), .b(FE_OFN1085_n_13221), .o(g54194_db) );
in01f01 g62899_u0 ( .a(FE_OFN1214_n_4151), .o(g62899_sb) );
na02m02 TIMEBOOST_cell_25987 ( .a(g65375_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q), .o(TIMEBOOST_net_7098) );
na02f02 TIMEBOOST_cell_38753 ( .a(TIMEBOOST_net_10988), .b(g65856_db), .o(n_1582) );
na02m02 TIMEBOOST_cell_68107 ( .a(TIMEBOOST_net_21261), .b(g61880_sb), .o(TIMEBOOST_net_17293) );
in01f02 g62900_u0 ( .a(FE_OFN1284_n_4097), .o(g62900_sb) );
na03m02 TIMEBOOST_cell_65611 ( .a(TIMEBOOST_net_12839), .b(g64228_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q), .o(TIMEBOOST_net_15071) );
na02s01 TIMEBOOST_cell_48641 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q), .b(g58453_sb), .o(TIMEBOOST_net_14538) );
na04f02 TIMEBOOST_cell_67235 ( .a(g64967_sb), .b(FE_OFN619_n_4490), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q), .d(n_4444), .o(n_4374) );
in01f04 g62901_u0 ( .a(FE_OFN1322_n_6436), .o(g62901_sb) );
no02f04 TIMEBOOST_cell_3835 ( .a(TIMEBOOST_net_477), .b(n_13340), .o(n_13907) );
na02f08 TIMEBOOST_cell_71837 ( .a(TIMEBOOST_net_23126), .b(parchk_pci_cbe_out_in), .o(n_2376) );
in01f02 g62902_u0 ( .a(FE_OFN1316_n_6624), .o(g62902_sb) );
na03f02 TIMEBOOST_cell_65362 ( .a(TIMEBOOST_net_16312), .b(n_5633), .c(g62133_sb), .o(n_5561) );
na02f02 TIMEBOOST_cell_3837 ( .a(n_12714), .b(TIMEBOOST_net_478), .o(n_15937) );
in01f02 g62903_u0 ( .a(FE_OFN1264_n_4095), .o(g62903_sb) );
na03f02 TIMEBOOST_cell_73396 ( .a(TIMEBOOST_net_16722), .b(FE_OFN1180_n_3476), .c(g60631_sb), .o(n_5705) );
in01f01 g62904_u0 ( .a(FE_OFN1250_n_4093), .o(g62904_sb) );
na02s02 TIMEBOOST_cell_49211 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q), .b(g65820_sb), .o(TIMEBOOST_net_14823) );
na02s02 TIMEBOOST_cell_68281 ( .a(TIMEBOOST_net_21348), .b(TIMEBOOST_net_14162), .o(n_2189) );
no02s01 TIMEBOOST_cell_44973 ( .a(FE_RN_284_0), .b(parchk_pci_cbe_out_in), .o(TIMEBOOST_net_13381) );
in01f02 g62905_u0 ( .a(n_6287), .o(g62905_sb) );
na02s02 TIMEBOOST_cell_48853 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q), .b(FE_OFN221_n_9846), .o(TIMEBOOST_net_14644) );
na02f01 TIMEBOOST_cell_3402 ( .a(n_4718), .b(n_2087), .o(TIMEBOOST_net_261) );
in01f02 g62906_u0 ( .a(FE_OFN1315_n_6624), .o(g62906_sb) );
na03s01 TIMEBOOST_cell_64500 ( .a(TIMEBOOST_net_14055), .b(g65861_sb), .c(TIMEBOOST_net_20847), .o(n_7915) );
in01s01 TIMEBOOST_cell_73964 ( .a(wbm_dat_i_31_), .o(TIMEBOOST_net_23529) );
na02m02 TIMEBOOST_cell_72124 ( .a(TIMEBOOST_net_20351), .b(FE_OFN948_n_2248), .o(TIMEBOOST_net_23270) );
in01f01 g62907_u0 ( .a(FE_OFN1248_n_4093), .o(g62907_sb) );
in01s01 TIMEBOOST_cell_73971 ( .a(TIMEBOOST_net_23535), .o(TIMEBOOST_net_23536) );
na03f02 TIMEBOOST_cell_66907 ( .a(FE_OFN1733_n_16317), .b(TIMEBOOST_net_16487), .c(FE_OFN1738_n_11019), .o(n_12639) );
na02m02 TIMEBOOST_cell_43166 ( .a(TIMEBOOST_net_12477), .b(FE_OFN1797_n_2299), .o(TIMEBOOST_net_10746) );
in01f02 g62908_u0 ( .a(FE_OFN1258_n_4143), .o(g62908_sb) );
in01s01 TIMEBOOST_cell_45887 ( .a(parchk_pci_ad_out_in_1170), .o(TIMEBOOST_net_13848) );
na02m06 TIMEBOOST_cell_69058 ( .a(FE_OFN615_n_4501), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q), .o(TIMEBOOST_net_21737) );
in01f02 g62909_u0 ( .a(FE_OFN1231_n_6391), .o(g62909_sb) );
na02s01 TIMEBOOST_cell_27997 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q), .o(TIMEBOOST_net_8103) );
na03f02 TIMEBOOST_cell_73559 ( .a(TIMEBOOST_net_17080), .b(FE_OFN1230_n_6391), .c(g62975_sb), .o(n_5932) );
in01m01 g62910_u0 ( .a(FE_OFN1278_n_4097), .o(g62910_sb) );
in01s01 TIMEBOOST_cell_45888 ( .a(TIMEBOOST_net_13848), .o(TIMEBOOST_net_13849) );
na02m04 TIMEBOOST_cell_48645 ( .a(n_3744), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q), .o(TIMEBOOST_net_14540) );
in01f02 g62911_u0 ( .a(n_6287), .o(g62911_sb) );
na02f01 TIMEBOOST_cell_3403 ( .a(TIMEBOOST_net_261), .b(n_3314), .o(n_3402) );
na02f02 TIMEBOOST_cell_68229 ( .a(TIMEBOOST_net_21322), .b(n_3123), .o(TIMEBOOST_net_7213) );
in01f02 g62912_u0 ( .a(FE_OFN1312_n_6624), .o(g62912_sb) );
na03m02 TIMEBOOST_cell_72924 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q), .b(g65289_sb), .c(TIMEBOOST_net_22122), .o(TIMEBOOST_net_20539) );
in01f01 g62913_u0 ( .a(FE_OFN1212_n_4151), .o(g62913_sb) );
in01s01 TIMEBOOST_cell_45889 ( .a(TIMEBOOST_net_13850), .o(wbs_adr_i_30_) );
na02f02 TIMEBOOST_cell_3217 ( .a(TIMEBOOST_net_168), .b(n_2477), .o(n_2478) );
na03f02 TIMEBOOST_cell_66754 ( .a(TIMEBOOST_net_17393), .b(FE_OFN1213_n_4151), .c(g62464_sb), .o(n_6668) );
in01f02 g62914_u0 ( .a(FE_OFN1276_n_4096), .o(g62914_sb) );
in01s01 TIMEBOOST_cell_45890 ( .a(TIMEBOOST_net_13851), .o(TIMEBOOST_net_13850) );
na03m02 TIMEBOOST_cell_72801 ( .a(TIMEBOOST_net_21550), .b(g65744_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q), .o(TIMEBOOST_net_22865) );
na03s02 TIMEBOOST_cell_41947 ( .a(FE_OFN215_n_9856), .b(g58234_sb), .c(g58234_db), .o(n_9557) );
in01f01 g62915_u0 ( .a(FE_OFN1204_n_4090), .o(g62915_sb) );
na02s01 TIMEBOOST_cell_25993 ( .a(pci_target_unit_del_sync_addr_in_215), .b(parchk_pci_ad_reg_in_1216), .o(TIMEBOOST_net_7101) );
na03m02 TIMEBOOST_cell_72639 ( .a(g65025_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q), .c(TIMEBOOST_net_10637), .o(TIMEBOOST_net_20520) );
na04f04 TIMEBOOST_cell_42139 ( .a(configuration_wb_err_data_586), .b(FE_OFN1173_n_5592), .c(parchk_pci_ad_out_in_1183), .d(g62086_sb), .o(n_5622) );
in01f02 g62916_u0 ( .a(FE_OFN1193_n_6935), .o(g62916_sb) );
na02s01 TIMEBOOST_cell_25994 ( .a(TIMEBOOST_net_7101), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_5440) );
na02m02 TIMEBOOST_cell_70106 ( .a(g65332_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q), .o(TIMEBOOST_net_22261) );
na04f02 TIMEBOOST_cell_73057 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q), .b(FE_OFN2081_n_8176), .c(n_2061), .d(g61718_sb), .o(n_8389) );
in01f04 g62917_u0 ( .a(FE_OFN1248_n_4093), .o(g62917_sb) );
na02s01 TIMEBOOST_cell_25995 ( .a(pci_target_unit_del_sync_addr_in_234), .b(parchk_pci_ad_reg_in_1235), .o(TIMEBOOST_net_7102) );
na02m06 TIMEBOOST_cell_48649 ( .a(n_3774), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q), .o(TIMEBOOST_net_14542) );
na02s02 TIMEBOOST_cell_30593 ( .a(n_9735), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q), .o(TIMEBOOST_net_9401) );
in01f04 g62918_u0 ( .a(FE_OFN1248_n_4093), .o(g62918_sb) );
na03s02 TIMEBOOST_cell_65187 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q), .b(g65809_sb), .c(g65809_db), .o(n_1904) );
in01f02 g62919_u0 ( .a(n_6554), .o(g62919_sb) );
na02m02 TIMEBOOST_cell_70019 ( .a(TIMEBOOST_net_22217), .b(g61753_sb), .o(n_8309) );
na02f08 TIMEBOOST_cell_3405 ( .a(n_2180), .b(TIMEBOOST_net_262), .o(n_3024) );
na02f02 TIMEBOOST_cell_71610 ( .a(TIMEBOOST_net_16041), .b(n_12099), .o(TIMEBOOST_net_23013) );
in01f01 g62920_u0 ( .a(FE_OFN1226_n_6391), .o(g62920_sb) );
na02s01 TIMEBOOST_cell_25997 ( .a(pci_target_unit_del_sync_addr_in_231), .b(parchk_pci_ad_reg_in_1232), .o(TIMEBOOST_net_7103) );
na02s01 TIMEBOOST_cell_62648 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q), .o(TIMEBOOST_net_20271) );
na03m02 TIMEBOOST_cell_65134 ( .a(n_3774), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q), .c(FE_OFN618_n_4490), .o(TIMEBOOST_net_16238) );
in01f02 g62921_u0 ( .a(n_6232), .o(g62921_sb) );
na02m06 TIMEBOOST_cell_68664 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q), .b(FE_OFN686_n_4417), .o(TIMEBOOST_net_21540) );
na02f10 TIMEBOOST_cell_3407 ( .a(TIMEBOOST_net_263), .b(n_2176), .o(n_3073) );
na02m02 TIMEBOOST_cell_3408 ( .a(n_2463), .b(n_2596), .o(TIMEBOOST_net_264) );
in01f01 g62922_u0 ( .a(FE_OFN1244_n_4092), .o(g62922_sb) );
na03m02 TIMEBOOST_cell_72623 ( .a(n_4473), .b(FE_OFN640_n_4669), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q), .o(TIMEBOOST_net_23238) );
na02f02 TIMEBOOST_cell_69033 ( .a(TIMEBOOST_net_21724), .b(g65262_sb), .o(TIMEBOOST_net_20917) );
in01f01 g62923_u0 ( .a(FE_OFN1272_n_4096), .o(g62923_sb) );
na02s01 TIMEBOOST_cell_25999 ( .a(pci_target_unit_del_sync_addr_in_225), .b(parchk_pci_ad_reg_in_1226), .o(TIMEBOOST_net_7104) );
na02f04 TIMEBOOST_cell_3023 ( .a(TIMEBOOST_net_71), .b(n_1168), .o(n_3080) );
na03s02 TIMEBOOST_cell_41995 ( .a(g58405_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q), .c(g58405_db), .o(n_9002) );
in01f02 g62924_u0 ( .a(n_6645), .o(g62924_sb) );
na02s01 TIMEBOOST_cell_27999 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q), .o(TIMEBOOST_net_8104) );
na02f02 TIMEBOOST_cell_3409 ( .a(n_2738), .b(TIMEBOOST_net_264), .o(n_2989) );
in01f01 g62925_u0 ( .a(FE_OFN1192_n_6935), .o(g62925_sb) );
na03f02 TIMEBOOST_cell_73723 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13603), .c(FE_OFN1577_n_12028), .o(n_12749) );
na02f02 g62925_u2 ( .a(n_4261), .b(FE_OFN1192_n_6935), .o(g62925_db) );
in01f02 g62926_u0 ( .a(n_6232), .o(g62926_sb) );
na03m02 TIMEBOOST_cell_73038 ( .a(TIMEBOOST_net_21822), .b(FE_OFN1679_n_4655), .c(TIMEBOOST_net_22069), .o(TIMEBOOST_net_17420) );
na02f04 TIMEBOOST_cell_3411 ( .a(TIMEBOOST_net_265), .b(n_2738), .o(n_3174) );
in01m01 g62927_u0 ( .a(FE_OFN1244_n_4092), .o(g62927_sb) );
na02s01 TIMEBOOST_cell_26000 ( .a(TIMEBOOST_net_7104), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_5449) );
na03f02 TIMEBOOST_cell_73397 ( .a(TIMEBOOST_net_16441), .b(FE_OFN1184_n_3476), .c(g60612_sb), .o(n_4842) );
in01f01 g62928_u0 ( .a(FE_OFN1202_n_4090), .o(g62928_sb) );
na02s01 TIMEBOOST_cell_26001 ( .a(pci_target_unit_del_sync_addr_in_230), .b(parchk_pci_ad_reg_in_1231), .o(TIMEBOOST_net_7105) );
na02m02 TIMEBOOST_cell_69099 ( .a(TIMEBOOST_net_21757), .b(g65274_sb), .o(TIMEBOOST_net_12550) );
na03f02 TIMEBOOST_cell_66744 ( .a(TIMEBOOST_net_16825), .b(FE_OFN1306_n_13124), .c(g54365_sb), .o(n_13077) );
in01f01 g62929_u0 ( .a(FE_OFN1248_n_4093), .o(g62929_sb) );
na03m02 TIMEBOOST_cell_72625 ( .a(g65039_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q), .c(TIMEBOOST_net_16232), .o(TIMEBOOST_net_17539) );
na03f02 TIMEBOOST_cell_72669 ( .a(TIMEBOOST_net_16584), .b(FE_OFN784_n_2678), .c(g65243_sb), .o(n_2639) );
na04f04 TIMEBOOST_cell_67604 ( .a(TIMEBOOST_net_16415), .b(TIMEBOOST_net_10435), .c(TIMEBOOST_net_6860), .d(g63438_sb), .o(n_4621) );
in01f01 g62930_u0 ( .a(FE_OFN1264_n_4095), .o(g62930_sb) );
na02s01 TIMEBOOST_cell_26003 ( .a(pci_target_unit_del_sync_addr_in_214), .b(parchk_pci_ad_reg_in_1215), .o(TIMEBOOST_net_7106) );
in01f02 g62931_u0 ( .a(FE_OFN1235_n_6391), .o(g62931_sb) );
na02f02 TIMEBOOST_cell_49553 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_400), .b(n_1786), .o(TIMEBOOST_net_14994) );
na03f02 TIMEBOOST_cell_73753 ( .a(TIMEBOOST_net_23382), .b(n_12099), .c(FE_OFN1757_n_12681), .o(n_12526) );
in01m01 g62932_u0 ( .a(FE_OFN1283_n_4097), .o(g62932_sb) );
na03f02 TIMEBOOST_cell_73398 ( .a(TIMEBOOST_net_16742), .b(FE_OFN1184_n_3476), .c(g60647_sb), .o(n_5679) );
na02f04 TIMEBOOST_cell_68607 ( .a(TIMEBOOST_net_21511), .b(n_2795), .o(n_3281) );
na02s01 TIMEBOOST_cell_43067 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_12428) );
in01f01 g62933_u0 ( .a(FE_OFN1276_n_4096), .o(g62933_sb) );
na02s01 TIMEBOOST_cell_26005 ( .a(pci_target_unit_del_sync_addr_in_223), .b(parchk_pci_ad_reg_in_1224), .o(TIMEBOOST_net_7107) );
na02f01 TIMEBOOST_cell_3035 ( .a(TIMEBOOST_net_77), .b(n_9175), .o(n_2276) );
na02f02 TIMEBOOST_cell_54390 ( .a(TIMEBOOST_net_17412), .b(FE_OFN1243_n_4092), .o(TIMEBOOST_net_15807) );
in01f01 g62934_u0 ( .a(FE_OFN1275_n_4096), .o(g62934_sb) );
na02s01 TIMEBOOST_cell_26006 ( .a(TIMEBOOST_net_7107), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_5442) );
na03f02 TIMEBOOST_cell_68550 ( .a(FE_OFN1001_n_15978), .b(conf_wb_err_bc_in_847), .c(n_213), .o(TIMEBOOST_net_21483) );
na03f02 TIMEBOOST_cell_73783 ( .a(TIMEBOOST_net_16517), .b(FE_OCP_RBN1996_n_13971), .c(FE_OFN1588_n_13736), .o(g53250_p) );
in01f01 g62935_u0 ( .a(FE_OFN1276_n_4096), .o(g62935_sb) );
na02s01 TIMEBOOST_cell_26007 ( .a(pci_target_unit_del_sync_addr_in_218), .b(parchk_pci_ad_reg_in_1219), .o(TIMEBOOST_net_7108) );
na03f02 TIMEBOOST_cell_73754 ( .a(n_13901), .b(TIMEBOOST_net_13694), .c(FE_OFN1593_n_13741), .o(g53243_p) );
na03f02 TIMEBOOST_cell_72629 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q), .c(TIMEBOOST_net_12821), .o(TIMEBOOST_net_20543) );
in01f02 g62936_u0 ( .a(FE_OFN1234_n_6391), .o(g62936_sb) );
na02m01 TIMEBOOST_cell_43783 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(FE_OFN928_n_4730), .o(TIMEBOOST_net_12786) );
na03f02 TIMEBOOST_cell_67993 ( .a(TIMEBOOST_net_17548), .b(FE_OFN1248_n_4093), .c(g62638_sb), .o(n_6273) );
na02m01 TIMEBOOST_cell_48485 ( .a(n_4394), .b(FE_OFN618_n_4490), .o(TIMEBOOST_net_14460) );
in01f01 g62937_u0 ( .a(FE_OFN1194_n_6935), .o(g62937_sb) );
na02m01 TIMEBOOST_cell_49337 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_134), .o(TIMEBOOST_net_14886) );
na02m02 TIMEBOOST_cell_3041 ( .a(TIMEBOOST_net_80), .b(n_1632), .o(n_1990) );
na03f02 TIMEBOOST_cell_67995 ( .a(TIMEBOOST_net_20528), .b(FE_OFN1283_n_4097), .c(g62896_sb), .o(n_6085) );
in01f02 g62938_u0 ( .a(FE_OFN1236_n_6391), .o(g62938_sb) );
na02m01 TIMEBOOST_cell_48405 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q), .o(TIMEBOOST_net_14420) );
na04s04 TIMEBOOST_cell_46769 ( .a(g58208_sb), .b(FE_OFN266_n_9884), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q), .d(g58208_db), .o(TIMEBOOST_net_9429) );
na03s02 TIMEBOOST_cell_72539 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q), .b(FE_OFN560_n_9895), .c(TIMEBOOST_net_12457), .o(TIMEBOOST_net_16997) );
in01f02 g62939_u0 ( .a(n_6431), .o(g62939_sb) );
in01s01 TIMEBOOST_cell_73848 ( .a(n_8530), .o(TIMEBOOST_net_23413) );
na02f02 TIMEBOOST_cell_71519 ( .a(TIMEBOOST_net_22967), .b(FE_OFN1566_n_12502), .o(n_12630) );
in01m02 g62940_u0 ( .a(FE_OFN1289_n_4098), .o(g62940_sb) );
na02s01 TIMEBOOST_cell_26009 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_145), .o(TIMEBOOST_net_7109) );
in01s01 TIMEBOOST_cell_73983 ( .a(TIMEBOOST_net_23547), .o(TIMEBOOST_net_23548) );
na02f02 TIMEBOOST_cell_50950 ( .a(TIMEBOOST_net_15692), .b(g62356_sb), .o(n_6887) );
in01f02 g62941_u0 ( .a(FE_OFN1233_n_6391), .o(g62941_sb) );
na02f02 TIMEBOOST_cell_69459 ( .a(TIMEBOOST_net_21937), .b(TIMEBOOST_net_14512), .o(TIMEBOOST_net_17106) );
na02f08 TIMEBOOST_cell_3557 ( .a(TIMEBOOST_net_338), .b(n_7216), .o(n_7704) );
na02f01 TIMEBOOST_cell_18026 ( .a(TIMEBOOST_net_5376), .b(FE_OCPN1832_n_16949), .o(n_1827) );
in01m01 g62942_u0 ( .a(FE_OFN1222_n_6391), .o(g62942_sb) );
na03s03 TIMEBOOST_cell_72362 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q), .b(pci_target_unit_fifos_pcir_data_in_183), .c(FE_OFN1784_n_1699), .o(TIMEBOOST_net_23136) );
na02f02 TIMEBOOST_cell_3247 ( .a(TIMEBOOST_net_183), .b(n_2754), .o(n_3200) );
na02f04 TIMEBOOST_cell_3248 ( .a(n_1436), .b(wishbone_slave_unit_pcim_if_del_burst_in), .o(TIMEBOOST_net_184) );
in01m01 g62943_u0 ( .a(FE_OFN1283_n_4097), .o(g62943_sb) );
na03f02 TIMEBOOST_cell_73698 ( .a(TIMEBOOST_net_13512), .b(FE_OFN1762_n_10780), .c(FE_OFN1583_n_12306), .o(n_12628) );
na02m02 TIMEBOOST_cell_71931 ( .a(TIMEBOOST_net_23173), .b(n_4470), .o(TIMEBOOST_net_15240) );
in01f02 g62944_u0 ( .a(FE_OFN1264_n_4095), .o(g62944_sb) );
na03m02 TIMEBOOST_cell_68482 ( .a(n_3780), .b(g65099_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q), .o(TIMEBOOST_net_21449) );
in01f02 g62945_u0 ( .a(FE_OFN1234_n_6391), .o(g62945_sb) );
na03f02 TIMEBOOST_cell_73341 ( .a(n_17039), .b(n_2768), .c(n_17027), .o(TIMEBOOST_net_431) );
na04f04 TIMEBOOST_cell_34995 ( .a(n_9591), .b(g57337_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q), .d(FE_OFN1370_n_8567), .o(n_11415) );
in01f01 g62946_u0 ( .a(FE_OFN1243_n_4092), .o(g62946_sb) );
na02f01 TIMEBOOST_cell_3048 ( .a(FE_RN_264_0), .b(n_16496), .o(TIMEBOOST_net_84) );
na02m10 TIMEBOOST_cell_45105 ( .a(pci_target_unit_pcit_if_strd_addr_in_687), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51), .o(TIMEBOOST_net_13447) );
in01f02 g62947_u0 ( .a(FE_OFN1315_n_6624), .o(g62947_sb) );
na02m02 TIMEBOOST_cell_49959 ( .a(TIMEBOOST_net_10926), .b(g64835_sb), .o(TIMEBOOST_net_15197) );
in01f02 g62948_u0 ( .a(FE_OFN1312_n_6624), .o(g62948_sb) );
na03m02 TIMEBOOST_cell_65902 ( .a(n_3869), .b(g63089_sb), .c(g63089_db), .o(n_5076) );
na03f02 TIMEBOOST_cell_66695 ( .a(TIMEBOOST_net_17135), .b(FE_OFN1310_n_6624), .c(g63178_sb), .o(n_5792) );
in01f02 g62949_u0 ( .a(FE_OFN1293_n_4098), .o(g62949_sb) );
na03m02 TIMEBOOST_cell_72367 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_1_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_0_), .c(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .o(TIMEBOOST_net_32) );
na02f04 TIMEBOOST_cell_3051 ( .a(TIMEBOOST_net_85), .b(n_2701), .o(n_2702) );
in01f01 g62950_u0 ( .a(FE_OFN1243_n_4092), .o(g62950_sb) );
na03f02 TIMEBOOST_cell_34839 ( .a(TIMEBOOST_net_9439), .b(FE_OFN1380_n_8567), .c(g57336_sb), .o(n_10393) );
in01s01 TIMEBOOST_cell_63563 ( .a(TIMEBOOST_net_20743), .o(TIMEBOOST_net_20742) );
in01f01 g62951_u0 ( .a(FE_OFN1272_n_4096), .o(g62951_sb) );
na03f02 TIMEBOOST_cell_70208 ( .a(n_13745), .b(n_15405), .c(n_2276), .o(TIMEBOOST_net_22312) );
na02f08 TIMEBOOST_cell_3055 ( .a(TIMEBOOST_net_87), .b(n_2236), .o(n_2706) );
na02m02 TIMEBOOST_cell_63740 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q), .b(FE_OFN2256_n_8060), .o(TIMEBOOST_net_20856) );
in01f02 g62952_u0 ( .a(FE_OFN1260_n_4143), .o(g62952_sb) );
na03m02 TIMEBOOST_cell_68322 ( .a(TIMEBOOST_net_21173), .b(g65873_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q), .o(TIMEBOOST_net_21369) );
na02f04 TIMEBOOST_cell_3057 ( .a(TIMEBOOST_net_88), .b(n_2229), .o(n_2230) );
na02f08 TIMEBOOST_cell_3058 ( .a(n_1824), .b(n_373), .o(TIMEBOOST_net_89) );
in01f02 g62953_u0 ( .a(FE_OFN2063_n_6391), .o(g62953_sb) );
na02s02 TIMEBOOST_cell_52422 ( .a(TIMEBOOST_net_16428), .b(g57949_sb), .o(TIMEBOOST_net_9463) );
na02f02 TIMEBOOST_cell_3561 ( .a(TIMEBOOST_net_340), .b(n_3202), .o(n_3491) );
na02f04 TIMEBOOST_cell_3562 ( .a(n_2754), .b(n_3192), .o(TIMEBOOST_net_341) );
in01m01 g62954_u0 ( .a(FE_OFN1295_n_4098), .o(g62954_sb) );
na02m01 TIMEBOOST_cell_53375 ( .a(n_2512), .b(pci_target_unit_pcit_if_strd_addr_in_691), .o(TIMEBOOST_net_16905) );
na02f08 TIMEBOOST_cell_3059 ( .a(TIMEBOOST_net_89), .b(n_8498), .o(n_2678) );
na03f02 TIMEBOOST_cell_33361 ( .a(TIMEBOOST_net_7309), .b(g54317_sb), .c(g54317_db), .o(n_13291) );
in01f02 g62955_u0 ( .a(FE_OFN1312_n_6624), .o(g62955_sb) );
na02m08 TIMEBOOST_cell_68454 ( .a(FE_OFN669_n_4505), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q), .o(TIMEBOOST_net_21435) );
na02s02 TIMEBOOST_cell_43507 ( .a(TIMEBOOST_net_21153), .b(g65724_sb), .o(TIMEBOOST_net_12648) );
na04m04 TIMEBOOST_cell_73058 ( .a(n_1648), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q), .c(FE_OFN710_n_8232), .d(g61951_sb), .o(n_7923) );
in01f02 g62956_u0 ( .a(FE_OFN1313_n_6624), .o(g62956_sb) );
na03f04 TIMEBOOST_cell_73489 ( .a(n_3290), .b(pciu_bar0_in_378), .c(n_3057), .o(TIMEBOOST_net_9576) );
na03m02 TIMEBOOST_cell_69018 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q), .b(FE_OFN1625_n_4438), .c(n_3774), .o(TIMEBOOST_net_21717) );
na02m02 TIMEBOOST_cell_69985 ( .a(TIMEBOOST_net_22200), .b(g61757_sb), .o(n_8299) );
in01f01 g62957_u0 ( .a(FE_OFN1250_n_4093), .o(g62957_sb) );
na02m06 TIMEBOOST_cell_52735 ( .a(pci_target_unit_pcit_if_strd_addr_in_695), .b(pci_target_unit_del_sync_addr_in_213), .o(TIMEBOOST_net_16585) );
na02f06 TIMEBOOST_cell_3062 ( .a(n_2411), .b(wbm_adr_o_2_), .o(TIMEBOOST_net_91) );
in01f01 g62958_u0 ( .a(FE_OFN1294_n_4098), .o(g62958_sb) );
na02s02 TIMEBOOST_cell_43803 ( .a(TIMEBOOST_net_23390), .b(FE_OFN1015_n_2053), .o(TIMEBOOST_net_12796) );
na02f06 TIMEBOOST_cell_3063 ( .a(TIMEBOOST_net_91), .b(n_1975), .o(n_2934) );
na02s01 TIMEBOOST_cell_53013 ( .a(configuration_pci_err_data), .b(wbm_dat_o_0_), .o(TIMEBOOST_net_16724) );
in01f01 g62959_u0 ( .a(FE_OFN1294_n_4098), .o(g62959_sb) );
na02m06 TIMEBOOST_cell_69721 ( .a(TIMEBOOST_net_22068), .b(g65351_sb), .o(TIMEBOOST_net_12742) );
na02s01 TIMEBOOST_cell_3066 ( .a(g65390_sb), .b(g65390_db), .o(TIMEBOOST_net_93) );
in01f02 g62960_u0 ( .a(FE_OFN1323_n_6436), .o(g62960_sb) );
na03m02 TIMEBOOST_cell_72598 ( .a(FE_OFN580_n_9531), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q), .c(FE_OFN268_n_9880), .o(TIMEBOOST_net_22867) );
na02f02 TIMEBOOST_cell_38067 ( .a(g58401_db), .b(TIMEBOOST_net_10645), .o(n_9004) );
in01f02 g62961_u0 ( .a(FE_OFN1312_n_6624), .o(g62961_sb) );
na02f02 TIMEBOOST_cell_50158 ( .a(TIMEBOOST_net_15296), .b(g60662_sb), .o(n_5657) );
in01f02 g62962_u0 ( .a(FE_OFN1293_n_4098), .o(g62962_sb) );
na02m01 TIMEBOOST_cell_26018 ( .a(TIMEBOOST_net_7113), .b(FE_OFN2256_n_8060), .o(TIMEBOOST_net_5468) );
na02s01 TIMEBOOST_cell_3067 ( .a(TIMEBOOST_net_93), .b(n_2675), .o(n_2630) );
in01f02 g62963_u0 ( .a(FE_OFN1223_n_6391), .o(g62963_sb) );
na02m02 TIMEBOOST_cell_68899 ( .a(TIMEBOOST_net_21657), .b(g65888_db), .o(TIMEBOOST_net_17456) );
na03f02 TIMEBOOST_cell_73823 ( .a(TIMEBOOST_net_13790), .b(n_13873), .c(FE_OFN1593_n_13741), .o(n_16211) );
in01f02 g62964_u0 ( .a(n_6287), .o(g62964_sb) );
na02f02 TIMEBOOST_cell_53470 ( .a(TIMEBOOST_net_16952), .b(g61758_sb), .o(n_8297) );
na02m04 TIMEBOOST_cell_48769 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q), .b(n_3752), .o(TIMEBOOST_net_14602) );
na03f02 TIMEBOOST_cell_73784 ( .a(TIMEBOOST_net_16521), .b(FE_OCP_RBN1996_n_13971), .c(FE_OFN1588_n_13736), .o(g53235_p) );
in01f02 g62965_u0 ( .a(FE_OFN1270_n_4095), .o(g62965_sb) );
no02f06 TIMEBOOST_cell_3069 ( .a(TIMEBOOST_net_94), .b(n_16286), .o(n_16288) );
na03f02 TIMEBOOST_cell_34757 ( .a(TIMEBOOST_net_9409), .b(FE_OFN1392_n_8567), .c(g57363_sb), .o(n_11384) );
in01f01 g62966_u0 ( .a(FE_OFN1226_n_6391), .o(g62966_sb) );
na02m02 TIMEBOOST_cell_69016 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q), .o(TIMEBOOST_net_21716) );
na02f03 TIMEBOOST_cell_50105 ( .a(pciu_bar0_in_371), .b(n_4806), .o(TIMEBOOST_net_15270) );
in01f02 g62967_u0 ( .a(FE_OFN1323_n_6436), .o(g62967_sb) );
na03f02 TIMEBOOST_cell_66804 ( .a(n_4617), .b(g61698_sb), .c(g61698_db), .o(n_5716) );
na03s02 TIMEBOOST_cell_46600 ( .a(TIMEBOOST_net_12834), .b(g63605_sb), .c(g63605_db), .o(n_7165) );
na02s02 TIMEBOOST_cell_68776 ( .a(TIMEBOOST_net_20210), .b(FE_OFN953_n_2055), .o(TIMEBOOST_net_21596) );
in01f02 g62968_u0 ( .a(FE_OFN1317_n_6624), .o(g62968_sb) );
na02s01 TIMEBOOST_cell_48152 ( .a(TIMEBOOST_net_14293), .b(FE_OFN223_n_9844), .o(TIMEBOOST_net_10500) );
na04f04 TIMEBOOST_cell_73059 ( .a(n_1599), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q), .c(FE_OFN712_n_8140), .d(g61824_sb), .o(n_8139) );
in01f02 g62969_u0 ( .a(n_6287), .o(g62969_sb) );
na02m01 TIMEBOOST_cell_68530 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q), .b(n_3764), .o(TIMEBOOST_net_21473) );
na02m10 TIMEBOOST_cell_45323 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q), .o(TIMEBOOST_net_13556) );
no02f10 TIMEBOOST_cell_3418 ( .a(FE_OCPN1843_n_16033), .b(n_15999), .o(TIMEBOOST_net_269) );
in01f01 g62970_u0 ( .a(FE_OFN1257_n_4143), .o(g62970_sb) );
na03s01 TIMEBOOST_cell_41657 ( .a(g57953_sb), .b(FE_OFN217_n_9889), .c(g57953_db), .o(n_9855) );
na02m02 TIMEBOOST_cell_3072 ( .a(parchk_pci_par_en_in), .b(n_1089), .o(TIMEBOOST_net_96) );
in01f02 g62971_u0 ( .a(FE_OFN1234_n_6391), .o(g62971_sb) );
no02f20 TIMEBOOST_cell_44074 ( .a(TIMEBOOST_net_12931), .b(FE_RN_67_0), .o(n_15403) );
na02f08 TIMEBOOST_cell_3563 ( .a(TIMEBOOST_net_341), .b(n_3202), .o(n_3193) );
in01m01 g62972_u0 ( .a(FE_OFN1218_n_6886), .o(g62972_sb) );
na03s02 TIMEBOOST_cell_41654 ( .a(g57922_sb), .b(FE_OFN219_n_9853), .c(g57922_db), .o(n_9888) );
na02m02 TIMEBOOST_cell_3073 ( .a(TIMEBOOST_net_96), .b(n_12855), .o(n_13332) );
no02s02 TIMEBOOST_cell_3074 ( .a(n_1460), .b(n_169), .o(TIMEBOOST_net_97) );
in01f02 g62973_u0 ( .a(n_6232), .o(g62973_sb) );
no02f20 TIMEBOOST_cell_3419 ( .a(TIMEBOOST_net_269), .b(FE_RN_149_0), .o(n_16810) );
na02s01 g65797_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q), .b(FE_OFN1786_n_1699), .o(g65797_db) );
in01m01 g62974_u0 ( .a(FE_OFN1213_n_4151), .o(g62974_sb) );
na03f02 TIMEBOOST_cell_67997 ( .a(TIMEBOOST_net_20973), .b(FE_OFN1284_n_4097), .c(g62543_sb), .o(n_6480) );
no02f01 TIMEBOOST_cell_3075 ( .a(TIMEBOOST_net_97), .b(n_1696), .o(g59232_BP) );
na03s02 TIMEBOOST_cell_72644 ( .a(TIMEBOOST_net_21415), .b(n_8272), .c(g61929_sb), .o(n_7965) );
in01f02 g62975_u0 ( .a(FE_OFN1230_n_6391), .o(g62975_sb) );
na02s02 TIMEBOOST_cell_38440 ( .a(FE_OFN213_n_9124), .b(g57919_sb), .o(TIMEBOOST_net_10832) );
na02f04 TIMEBOOST_cell_3565 ( .a(TIMEBOOST_net_342), .b(n_2971), .o(n_3179) );
na02m02 TIMEBOOST_cell_43051 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q), .b(FE_OFN631_n_4454), .o(TIMEBOOST_net_12420) );
in01f01 g62976_u0 ( .a(FE_OFN1285_n_4097), .o(g62976_sb) );
na03f06 TIMEBOOST_cell_73249 ( .a(TIMEBOOST_net_22291), .b(g64140_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q), .o(TIMEBOOST_net_22436) );
na02m02 TIMEBOOST_cell_3077 ( .a(TIMEBOOST_net_98), .b(FE_OFN992_n_2373), .o(n_7397) );
na02s04 TIMEBOOST_cell_3078 ( .a(n_1690), .b(n_1187), .o(TIMEBOOST_net_99) );
in01f02 g62977_u0 ( .a(FE_OFN1236_n_6391), .o(g62977_sb) );
na03f02 TIMEBOOST_cell_66350 ( .a(TIMEBOOST_net_17075), .b(FE_OFN2064_n_6391), .c(g62381_sb), .o(n_6840) );
na02f02 TIMEBOOST_cell_44122 ( .a(TIMEBOOST_net_12955), .b(g63117_sb), .o(n_7117) );
na02f02 TIMEBOOST_cell_70987 ( .a(TIMEBOOST_net_22701), .b(g62334_sb), .o(n_6932) );
in01f02 g62978_u0 ( .a(n_6232), .o(g62978_sb) );
na02f04 TIMEBOOST_cell_3422 ( .a(n_1358), .b(conf_wb_err_addr_in_943), .o(TIMEBOOST_net_271) );
in01f02 g62979_u0 ( .a(n_6319), .o(g62979_sb) );
na02f06 TIMEBOOST_cell_3423 ( .a(TIMEBOOST_net_271), .b(n_2397), .o(n_2266) );
in01f02 g62980_u0 ( .a(FE_OFN1231_n_6391), .o(g62980_sb) );
na02m02 TIMEBOOST_cell_63063 ( .a(TIMEBOOST_net_20478), .b(g58097_sb), .o(TIMEBOOST_net_16672) );
na03f02 TIMEBOOST_cell_34814 ( .a(TIMEBOOST_net_9442), .b(FE_OFN1392_n_8567), .c(g57493_sb), .o(n_11243) );
na04f02 TIMEBOOST_cell_66034 ( .a(TIMEBOOST_net_315), .b(n_7039), .c(TIMEBOOST_net_399), .d(n_13679), .o(TIMEBOOST_net_11637) );
in01f02 g62981_u0 ( .a(FE_OFN1236_n_6391), .o(g62981_sb) );
na02m06 TIMEBOOST_cell_72218 ( .a(TIMEBOOST_net_10072), .b(configuration_wb_err_addr_541), .o(TIMEBOOST_net_23317) );
in01s01 TIMEBOOST_cell_73948 ( .a(wbm_dat_i_24_), .o(TIMEBOOST_net_23513) );
in01f02 g62982_u0 ( .a(FE_OFN1231_n_6391), .o(g62982_sb) );
na02s02 TIMEBOOST_cell_52427 ( .a(g58255_sb), .b(FE_OFN245_n_9114), .o(TIMEBOOST_net_16431) );
na02m10 TIMEBOOST_cell_28027 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q), .o(TIMEBOOST_net_8118) );
in01f02 g62983_u0 ( .a(FE_OFN1311_n_6624), .o(g62983_sb) );
in01s01 TIMEBOOST_cell_73984 ( .a(n_5790), .o(TIMEBOOST_net_23549) );
na02f02 TIMEBOOST_cell_69461 ( .a(TIMEBOOST_net_21938), .b(FE_OFN1797_n_2299), .o(n_2155) );
na02s01 TIMEBOOST_cell_53071 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q), .b(g57965_sb), .o(TIMEBOOST_net_16753) );
in01m01 g62984_u0 ( .a(FE_OFN1219_n_6886), .o(g62984_sb) );
na03s02 TIMEBOOST_cell_41661 ( .a(g58244_sb), .b(FE_OFN227_n_9841), .c(g58245_db), .o(n_9547) );
na02f02 TIMEBOOST_cell_3079 ( .a(TIMEBOOST_net_99), .b(n_1438), .o(n_2295) );
na02m10 TIMEBOOST_cell_3080 ( .a(n_1689), .b(n_1186), .o(TIMEBOOST_net_100) );
in01f02 g62985_u0 ( .a(FE_OFN1230_n_6391), .o(g62985_sb) );
na02s04 TIMEBOOST_cell_43754 ( .a(TIMEBOOST_net_12771), .b(g58100_sb), .o(n_9700) );
na04f04 TIMEBOOST_cell_73317 ( .a(n_4025), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q), .c(FE_OFN1112_g64577_p), .d(g62855_sb), .o(n_5258) );
in01f01 g62986_u0 ( .a(FE_OFN1207_n_6356), .o(g62986_sb) );
na03f02 TIMEBOOST_cell_73699 ( .a(TIMEBOOST_net_13515), .b(FE_OFN1762_n_10780), .c(FE_OFN1583_n_12306), .o(n_12747) );
na02m08 TIMEBOOST_cell_3081 ( .a(TIMEBOOST_net_100), .b(n_1476), .o(n_2275) );
no02f10 TIMEBOOST_cell_3082 ( .a(n_564), .b(n_2263), .o(TIMEBOOST_net_101) );
in01f02 g62987_u0 ( .a(FE_OFN1230_n_6391), .o(g62987_sb) );
na03s02 TIMEBOOST_cell_41660 ( .a(g58183_sb), .b(FE_OFN227_n_9841), .c(g58183_db), .o(n_9604) );
na02s01 TIMEBOOST_cell_63062 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q), .o(TIMEBOOST_net_20478) );
na03s02 TIMEBOOST_cell_69672 ( .a(TIMEBOOST_net_14079), .b(g65863_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q), .o(TIMEBOOST_net_22044) );
in01f02 g62988_u0 ( .a(FE_OFN1314_n_6624), .o(g62988_sb) );
in01m01 g62989_u0 ( .a(FE_OFN1295_n_4098), .o(g62989_sb) );
na02m02 TIMEBOOST_cell_49678 ( .a(TIMEBOOST_net_15056), .b(g61756_sb), .o(n_8302) );
no02f04 TIMEBOOST_cell_3084 ( .a(n_2263), .b(wishbone_slave_unit_pcim_sm_be_in_557), .o(TIMEBOOST_net_102) );
in01f02 g62990_u0 ( .a(n_6319), .o(g62990_sb) );
na02s02 TIMEBOOST_cell_68286 ( .a(TIMEBOOST_net_17200), .b(FE_OFN938_n_2292), .o(TIMEBOOST_net_21351) );
na03f02 TIMEBOOST_cell_73755 ( .a(n_13901), .b(TIMEBOOST_net_13697), .c(FE_OFN1593_n_13741), .o(g53276_p) );
na02s01 TIMEBOOST_cell_3426 ( .a(FE_OCPN1875_n_14526), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(TIMEBOOST_net_273) );
in01f01 g62991_u0 ( .a(FE_OFN1276_n_4096), .o(g62991_sb) );
na02s02 TIMEBOOST_cell_52428 ( .a(TIMEBOOST_net_16431), .b(g58255_db), .o(n_9041) );
na03f02 TIMEBOOST_cell_66909 ( .a(FE_OFN1735_n_16317), .b(TIMEBOOST_net_16002), .c(FE_OFN1741_n_11019), .o(n_12757) );
in01f02 g62992_u0 ( .a(n_6319), .o(g62992_sb) );
na02f02 TIMEBOOST_cell_3427 ( .a(n_15014), .b(TIMEBOOST_net_273), .o(n_7329) );
na02s01 TIMEBOOST_cell_45325 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q), .o(TIMEBOOST_net_13557) );
in01f01 g62993_u0 ( .a(FE_OFN1272_n_4096), .o(g62993_sb) );
na04f04 TIMEBOOST_cell_73318 ( .a(n_3955), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q), .c(FE_OFN1135_g64577_p), .d(g62813_sb), .o(n_5351) );
in01s01 TIMEBOOST_cell_45960 ( .a(TIMEBOOST_net_13921), .o(TIMEBOOST_net_13920) );
na02m04 TIMEBOOST_cell_68532 ( .a(n_3747), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q), .o(TIMEBOOST_net_21474) );
in01m01 g62994_u0 ( .a(FE_OFN1225_n_6391), .o(g62994_sb) );
na03s06 TIMEBOOST_cell_69252 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q), .c(FE_OFN956_n_1699), .o(TIMEBOOST_net_21834) );
na03f02 TIMEBOOST_cell_34769 ( .a(TIMEBOOST_net_9363), .b(FE_OFN1404_n_8567), .c(g57277_sb), .o(n_11477) );
na03f02 TIMEBOOST_cell_34773 ( .a(TIMEBOOST_net_9353), .b(FE_OFN1413_n_8567), .c(g57056_sb), .o(n_10508) );
in01m01 g62995_u0 ( .a(FE_OFN1193_n_6935), .o(g62995_sb) );
na03s02 TIMEBOOST_cell_33425 ( .a(FE_OFN270_n_9836), .b(g57996_sb), .c(g57996_db), .o(n_9798) );
na04s01 TIMEBOOST_cell_68002 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN529_n_9899), .c(FE_OFN207_n_9865), .d(g58008_sb), .o(n_9786) );
in01f02 g62996_u0 ( .a(n_6319), .o(g62996_sb) );
na02m01 TIMEBOOST_cell_71888 ( .a(n_3761), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q), .o(TIMEBOOST_net_23152) );
na02m01 TIMEBOOST_cell_71852 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q), .b(n_3783), .o(TIMEBOOST_net_23134) );
in01s01 TIMEBOOST_cell_63543 ( .a(TIMEBOOST_net_20723), .o(TIMEBOOST_net_20722) );
in01m01 g62997_u0 ( .a(FE_OFN1225_n_6391), .o(g62997_sb) );
na02m10 TIMEBOOST_cell_45403 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q), .o(TIMEBOOST_net_13596) );
na02m01 TIMEBOOST_cell_3095 ( .a(TIMEBOOST_net_107), .b(g65907_sb), .o(n_2151) );
in01f02 g62998_u0 ( .a(FE_OFN1320_n_6436), .o(g62998_sb) );
na02f01 TIMEBOOST_cell_44308 ( .a(TIMEBOOST_net_13048), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_11360) );
na02m03 TIMEBOOST_cell_69318 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q), .b(n_4482), .o(TIMEBOOST_net_21867) );
in01f02 g62999_u0 ( .a(FE_OFN1200_n_4090), .o(g62999_sb) );
na04f04 TIMEBOOST_cell_73319 ( .a(n_4045), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q), .c(FE_OFN1139_g64577_p), .d(g62748_sb), .o(n_5483) );
na02s01 TIMEBOOST_cell_44021 ( .a(FE_OFN555_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q), .o(TIMEBOOST_net_12905) );
in01s08 TIMEBOOST_cell_45930 ( .a(TIMEBOOST_net_13890), .o(TIMEBOOST_net_13891) );
in01f02 g63000_u0 ( .a(FE_OFN1230_n_6391), .o(g63000_sb) );
in01s01 TIMEBOOST_cell_63579 ( .a(TIMEBOOST_net_20758), .o(TIMEBOOST_net_20759) );
na03s02 TIMEBOOST_cell_65098 ( .a(g58264_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q), .c(TIMEBOOST_net_10772), .o(TIMEBOOST_net_9335) );
in01f01 g63001_u0 ( .a(FE_OFN1214_n_4151), .o(g63001_sb) );
na02m01 TIMEBOOST_cell_3099 ( .a(TIMEBOOST_net_109), .b(g65810_sb), .o(n_2186) );
in01f02 g63002_u0 ( .a(FE_OFN1272_n_4096), .o(g63002_sb) );
na02m02 TIMEBOOST_cell_54500 ( .a(TIMEBOOST_net_17467), .b(FE_OFN1242_n_4092), .o(TIMEBOOST_net_15818) );
na02m01 TIMEBOOST_cell_68450 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q), .b(FE_OFN671_n_4505), .o(TIMEBOOST_net_21433) );
in01f02 g63003_u0 ( .a(n_6645), .o(g63003_sb) );
na03f02 TIMEBOOST_cell_73576 ( .a(TIMEBOOST_net_17375), .b(FE_OFN1213_n_4151), .c(g62586_sb), .o(n_6379) );
na02m02 TIMEBOOST_cell_3431 ( .a(TIMEBOOST_net_275), .b(n_3437), .o(n_4591) );
na02m02 TIMEBOOST_cell_30935 ( .a(n_9710), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q), .o(TIMEBOOST_net_9572) );
in01f02 g63004_u0 ( .a(FE_OFN1317_n_6624), .o(g63004_sb) );
na02m02 TIMEBOOST_cell_54233 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q), .b(TIMEBOOST_net_13201), .o(TIMEBOOST_net_17334) );
na02s01 TIMEBOOST_cell_38042 ( .a(FE_OFN225_n_9122), .b(g57958_sb), .o(TIMEBOOST_net_10633) );
in01f02 g63005_u0 ( .a(FE_OFN1234_n_6391), .o(g63005_sb) );
na02m01 TIMEBOOST_cell_44077 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(FE_OFN1055_n_4727), .o(TIMEBOOST_net_12933) );
na03f02 TIMEBOOST_cell_66894 ( .a(FE_OFN1747_n_12004), .b(n_12010), .c(TIMEBOOST_net_13552), .o(n_12615) );
na03f02 TIMEBOOST_cell_73629 ( .a(TIMEBOOST_net_16813), .b(n_16748), .c(g52643_sb), .o(n_14747) );
in01f02 g63006_u0 ( .a(FE_OFN1196_n_4090), .o(g63006_sb) );
na04m06 TIMEBOOST_cell_72917 ( .a(TIMEBOOST_net_21171), .b(FE_OFN1041_n_2037), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q), .d(g65887_sb), .o(n_1862) );
na03m02 TIMEBOOST_cell_64497 ( .a(FE_OFN576_n_9902), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q), .c(TIMEBOOST_net_10855), .o(TIMEBOOST_net_9493) );
in01f02 g63007_u0 ( .a(FE_OFN1258_n_4143), .o(g63007_sb) );
na03s02 TIMEBOOST_cell_67910 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q), .b(g65844_sb), .c(TIMEBOOST_net_14840), .o(n_1876) );
na02m10 TIMEBOOST_cell_53015 ( .a(configuration_pci_err_data_518), .b(wbm_dat_o_17_), .o(TIMEBOOST_net_16725) );
in01f02 g63008_u0 ( .a(FE_OFN1311_n_6624), .o(g63008_sb) );
na02s01 TIMEBOOST_cell_42797 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q), .o(TIMEBOOST_net_12293) );
na03f01 TIMEBOOST_cell_66862 ( .a(FE_OFN1584_n_12306), .b(FE_OFN1761_n_10780), .c(TIMEBOOST_net_13692), .o(n_12614) );
in01f02 g63009_u0 ( .a(FE_OFN1235_n_6391), .o(g63009_sb) );
na02m01 TIMEBOOST_cell_43565 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q), .o(TIMEBOOST_net_12677) );
na02f02 TIMEBOOST_cell_68719 ( .a(TIMEBOOST_net_21567), .b(g64327_sb), .o(TIMEBOOST_net_13044) );
in01m01 g63010_u0 ( .a(FE_OFN1134_g64577_p), .o(g63010_sb) );
na03f02 TIMEBOOST_cell_73516 ( .a(TIMEBOOST_net_13370), .b(n_6431), .c(g62647_sb), .o(n_6254) );
na02m01 TIMEBOOST_cell_68832 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q), .b(FE_OFN623_n_4409), .o(TIMEBOOST_net_21624) );
in01f01 g63011_u0 ( .a(FE_OFN1207_n_6356), .o(g63011_sb) );
na02m01 TIMEBOOST_cell_68552 ( .a(wishbone_slave_unit_pci_initiator_if_current_byte_address_36), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_384), .o(TIMEBOOST_net_21484) );
na02m02 TIMEBOOST_cell_64057 ( .a(TIMEBOOST_net_21014), .b(g58398_sb), .o(n_9436) );
in01m01 g63012_u0 ( .a(FE_OFN1121_g64577_p), .o(g63012_sb) );
na03m02 TIMEBOOST_cell_72925 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q), .b(g65368_sb), .c(TIMEBOOST_net_23241), .o(TIMEBOOST_net_17451) );
na02f01 TIMEBOOST_cell_71977 ( .a(TIMEBOOST_net_23196), .b(FE_OFN660_n_4392), .o(TIMEBOOST_net_14434) );
na03m06 TIMEBOOST_cell_68370 ( .a(FE_OFN906_n_4736), .b(TIMEBOOST_net_12324), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q), .o(TIMEBOOST_net_21393) );
in01m01 g63013_u0 ( .a(FE_OFN1104_g64577_p), .o(g63013_sb) );
na02m02 TIMEBOOST_cell_30681 ( .a(n_8998), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q), .o(TIMEBOOST_net_9445) );
na02m10 TIMEBOOST_cell_28995 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q), .o(TIMEBOOST_net_8602) );
in01f01 g63014_u0 ( .a(FE_OFN2105_g64577_p), .o(g63014_sb) );
na02s01 TIMEBOOST_cell_29255 ( .a(FE_OFN1654_n_9502), .b(FE_OFN227_n_9841), .o(TIMEBOOST_net_8732) );
na04f04 TIMEBOOST_cell_73320 ( .a(n_4075), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q), .c(FE_OFN2105_g64577_p), .d(g62722_sb), .o(n_5539) );
in01f02 g63015_u0 ( .a(FE_OFN1122_g64577_p), .o(g63015_sb) );
na03m02 TIMEBOOST_cell_72567 ( .a(TIMEBOOST_net_23146), .b(FE_OFN665_n_4495), .c(TIMEBOOST_net_21527), .o(TIMEBOOST_net_13367) );
na02s03 TIMEBOOST_cell_42998 ( .a(TIMEBOOST_net_12393), .b(g58787_sb), .o(n_9836) );
na03f01 TIMEBOOST_cell_73399 ( .a(TIMEBOOST_net_16734), .b(FE_OFN1185_n_3476), .c(g60607_sb), .o(n_4847) );
in01f01 g63016_u0 ( .a(FE_OFN1100_g64577_p), .o(g63016_sb) );
na04m02 TIMEBOOST_cell_67237 ( .a(FE_OFN651_n_4508), .b(g65408_sb), .c(TIMEBOOST_net_20241), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q), .o(TIMEBOOST_net_17134) );
na02f02 TIMEBOOST_cell_71691 ( .a(TIMEBOOST_net_23053), .b(FE_OFN1601_n_13995), .o(n_14451) );
in01f01 g63017_u0 ( .a(FE_OFN1134_g64577_p), .o(g63017_sb) );
na02m04 TIMEBOOST_cell_68422 ( .a(g64769_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q), .o(TIMEBOOST_net_21419) );
na02f01 TIMEBOOST_cell_54234 ( .a(TIMEBOOST_net_17334), .b(g58280_db), .o(TIMEBOOST_net_9510) );
na04f04 TIMEBOOST_cell_73195 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q), .b(FE_OFN1104_g64577_p), .c(n_3900), .d(g63058_sb), .o(n_5134) );
in01f01 g63018_u0 ( .a(FE_OFN2104_g64577_p), .o(g63018_sb) );
na03f02 TIMEBOOST_cell_73176 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q), .b(g64323_sb), .c(g64323_db), .o(n_3853) );
in01f02 g63019_u0 ( .a(FE_OFN2105_g64577_p), .o(g63019_sb) );
na02s02 TIMEBOOST_cell_63841 ( .a(TIMEBOOST_net_20906), .b(g58219_sb), .o(TIMEBOOST_net_20454) );
na02s02 TIMEBOOST_cell_39727 ( .a(TIMEBOOST_net_11475), .b(g57907_db), .o(n_9220) );
in01m01 g63020_u0 ( .a(FE_OFN1100_g64577_p), .o(g63020_sb) );
na04m06 TIMEBOOST_cell_67418 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q), .b(g58028_sb), .c(FE_OFN235_n_9834), .d(g58028_db), .o(TIMEBOOST_net_16839) );
na03s02 TIMEBOOST_cell_46606 ( .a(TIMEBOOST_net_12835), .b(g63614_sb), .c(g63614_db), .o(n_7147) );
in01m01 g63021_u0 ( .a(FE_OFN1116_g64577_p), .o(g63021_sb) );
na03f02 TIMEBOOST_cell_73630 ( .a(TIMEBOOST_net_13445), .b(n_16748), .c(g52651_sb), .o(n_14671) );
na02s01 TIMEBOOST_cell_63122 ( .a(FE_OFN551_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q), .o(TIMEBOOST_net_20508) );
in01m01 g63022_u0 ( .a(FE_OFN882_g64577_p), .o(g63022_sb) );
na02m01 TIMEBOOST_cell_62824 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q), .o(TIMEBOOST_net_20359) );
na02s03 TIMEBOOST_cell_48095 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q), .b(pci_target_unit_fifos_pcir_data_in_170), .o(TIMEBOOST_net_14265) );
na03f02 TIMEBOOST_cell_35064 ( .a(TIMEBOOST_net_9610), .b(FE_OFN1438_n_9372), .c(g58481_sb), .o(n_8977) );
in01m01 g63023_u0 ( .a(FE_OFN882_g64577_p), .o(g63023_sb) );
na04f04 TIMEBOOST_cell_73321 ( .a(n_3954), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q), .c(FE_OFN1115_g64577_p), .d(g62864_sb), .o(n_5237) );
na02f01 TIMEBOOST_cell_69653 ( .a(TIMEBOOST_net_22034), .b(FE_OFN707_n_8119), .o(TIMEBOOST_net_14794) );
na02m08 TIMEBOOST_cell_62468 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q), .b(pci_target_unit_fifos_pciw_cbe_in_154), .o(TIMEBOOST_net_20181) );
in01f02 g63024_u0 ( .a(FE_OFN1122_g64577_p), .o(g63024_sb) );
na02s01 TIMEBOOST_cell_64192 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q), .o(TIMEBOOST_net_21082) );
na03s02 TIMEBOOST_cell_65599 ( .a(n_1921), .b(TIMEBOOST_net_20600), .c(g61768_sb), .o(n_8274) );
na03f02 TIMEBOOST_cell_72954 ( .a(pci_target_unit_del_sync_addr_in_220), .b(g65246_sb), .c(TIMEBOOST_net_7158), .o(n_2636) );
na02s01 TIMEBOOST_cell_68910 ( .a(g57964_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q), .o(TIMEBOOST_net_21663) );
na02f02 TIMEBOOST_cell_70699 ( .a(TIMEBOOST_net_22557), .b(g63172_sb), .o(n_4951) );
in01f02 g63026_u0 ( .a(FE_OFN1122_g64577_p), .o(g63026_sb) );
in01m01 g63027_u0 ( .a(FE_OFN877_g64577_p), .o(g63027_sb) );
na02s02 TIMEBOOST_cell_68268 ( .a(TIMEBOOST_net_21147), .b(g65701_sb), .o(TIMEBOOST_net_21342) );
na02s01 TIMEBOOST_cell_54049 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q), .o(TIMEBOOST_net_17242) );
in01f01 g63028_u0 ( .a(FE_OFN1123_g64577_p), .o(g63028_sb) );
na02f02 TIMEBOOST_cell_71104 ( .a(TIMEBOOST_net_17480), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_22760) );
na02s02 TIMEBOOST_cell_48340 ( .a(TIMEBOOST_net_14387), .b(TIMEBOOST_net_10775), .o(TIMEBOOST_net_9527) );
na03f02 TIMEBOOST_cell_73700 ( .a(TIMEBOOST_net_13516), .b(FE_OFN1762_n_10780), .c(FE_OFN1583_n_12306), .o(n_12598) );
in01f02 g63029_u0 ( .a(n_6645), .o(g63029_sb) );
na02f02 TIMEBOOST_cell_3433 ( .a(TIMEBOOST_net_276), .b(n_3335), .o(n_3498) );
na02m01 TIMEBOOST_cell_62546 ( .a(pci_target_unit_fifos_pciw_addr_data_in_123), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_20220) );
in01f01 g63030_u0 ( .a(FE_OFN1118_g64577_p), .o(g63030_sb) );
na02f02 TIMEBOOST_cell_27191 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_7700) );
in01f01 g63031_u0 ( .a(FE_OFN1123_g64577_p), .o(g63031_sb) );
na02s02 TIMEBOOST_cell_37430 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(g65790_sb), .o(TIMEBOOST_net_10327) );
in01m01 g63032_u0 ( .a(FE_OFN1131_g64577_p), .o(g63032_sb) );
na02s01 TIMEBOOST_cell_29241 ( .a(configuration_wb_err_data_571), .b(parchk_pci_ad_out_in_1168), .o(TIMEBOOST_net_8725) );
na02s01 TIMEBOOST_cell_51865 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q), .b(FE_OFN205_n_9140), .o(TIMEBOOST_net_16150) );
na02m02 g65346_u1 ( .a(g65346_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q), .o(g65346_da) );
in01f04 g63033_u0 ( .a(FE_OFN1121_g64577_p), .o(g63033_sb) );
na02m01 TIMEBOOST_cell_29247 ( .a(n_3744), .b(FE_OFN1642_n_4671), .o(TIMEBOOST_net_8728) );
na02s01 TIMEBOOST_cell_48127 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q), .b(FE_OFN585_n_9692), .o(TIMEBOOST_net_14281) );
na02f02 TIMEBOOST_cell_50715 ( .a(FE_OFN1000_n_15978), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_394), .o(TIMEBOOST_net_15575) );
in01f02 g63034_u0 ( .a(FE_OFN1116_g64577_p), .o(g63034_sb) );
na03m02 TIMEBOOST_cell_72472 ( .a(FE_OFN1786_n_1699), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q), .c(TIMEBOOST_net_21409), .o(TIMEBOOST_net_17296) );
in01s01 TIMEBOOST_cell_64260 ( .a(TIMEBOOST_net_21116), .o(wishbone_slave_unit_del_sync_sync_req_comp_pending) );
na03f06 TIMEBOOST_cell_73250 ( .a(TIMEBOOST_net_16394), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .c(g52631_sb), .o(TIMEBOOST_net_7472) );
in01f01 g63035_u0 ( .a(FE_OFN1127_g64577_p), .o(g63035_sb) );
na02m10 TIMEBOOST_cell_28013 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q), .o(TIMEBOOST_net_8111) );
in01f02 g63036_u0 ( .a(FE_OFN1120_g64577_p), .o(g63036_sb) );
na02f01 TIMEBOOST_cell_26063 ( .a(pci_target_unit_pcit_if_strd_addr_in_705), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7136) );
in01s01 TIMEBOOST_cell_73894 ( .a(n_8178), .o(TIMEBOOST_net_23459) );
in01f04 g63037_u0 ( .a(FE_OFN1121_g64577_p), .o(g63037_sb) );
na02f01 TIMEBOOST_cell_68901 ( .a(TIMEBOOST_net_21658), .b(n_4442), .o(TIMEBOOST_net_20843) );
in01m01 g63038_u0 ( .a(FE_OFN1122_g64577_p), .o(g63038_sb) );
in01f01 g63039_u0 ( .a(FE_OFN1097_g64577_p), .o(g63039_sb) );
na02f02 TIMEBOOST_cell_69121 ( .a(TIMEBOOST_net_21768), .b(g63543_db), .o(TIMEBOOST_net_17284) );
na03m02 TIMEBOOST_cell_68886 ( .a(g64838_sb), .b(n_4442), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q), .o(TIMEBOOST_net_21651) );
in01m01 g63040_u0 ( .a(FE_OFN1133_g64577_p), .o(g63040_sb) );
na02s01 TIMEBOOST_cell_38516 ( .a(FE_OFN211_n_9858), .b(g58202_sb), .o(TIMEBOOST_net_10870) );
na03f02 TIMEBOOST_cell_47402 ( .a(FE_OFN1588_n_13736), .b(TIMEBOOST_net_13712), .c(FE_OCP_RBN1995_n_13971), .o(n_14295) );
in01m01 g63041_u0 ( .a(FE_OFN1133_g64577_p), .o(g63041_sb) );
in01f02 g63042_u0 ( .a(FE_OFN2064_n_6391), .o(g63042_sb) );
na02s03 TIMEBOOST_cell_68626 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_21521) );
na04m04 TIMEBOOST_cell_67832 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(FE_OFN918_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q), .d(g64340_sb), .o(n_3838) );
in01m06 g63043_u0 ( .a(FE_OFN1119_g64577_p), .o(g63043_sb) );
na02s01 TIMEBOOST_cell_28009 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q), .o(TIMEBOOST_net_8109) );
na03f10 TIMEBOOST_cell_46082 ( .a(FE_OFN2059_n_13447), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_385), .o(TIMEBOOST_net_13130) );
in01f01 g63044_u0 ( .a(FE_OFN1128_g64577_p), .o(g63044_sb) );
na02m02 TIMEBOOST_cell_69519 ( .a(TIMEBOOST_net_21967), .b(TIMEBOOST_net_10596), .o(TIMEBOOST_net_20526) );
na03m06 TIMEBOOST_cell_69062 ( .a(FE_OFN1010_n_4734), .b(pci_target_unit_fifos_pciw_addr_data_in_127), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q), .o(TIMEBOOST_net_21739) );
in01m04 g63045_u0 ( .a(FE_OFN1097_g64577_p), .o(g63045_sb) );
in01f01 g63046_u0 ( .a(FE_OFN1123_g64577_p), .o(g63046_sb) );
na03f02 TIMEBOOST_cell_73724 ( .a(FE_OFN1559_n_12042), .b(TIMEBOOST_net_13627), .c(FE_OFN1577_n_12028), .o(n_12689) );
in01s01 g63047_u0 ( .a(FE_OFN881_g64577_p), .o(g63047_sb) );
na02s01 TIMEBOOST_cell_54737 ( .a(g57947_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q), .o(TIMEBOOST_net_17586) );
na02m01 g63047_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q), .b(FE_OFN881_g64577_p), .o(g63047_db) );
na02s01 TIMEBOOST_cell_54738 ( .a(TIMEBOOST_net_17586), .b(TIMEBOOST_net_12966), .o(TIMEBOOST_net_9472) );
in01f01 g63048_u0 ( .a(FE_OFN1094_g64577_p), .o(g63048_sb) );
na03m08 TIMEBOOST_cell_68948 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q), .b(g65302_sb), .c(FE_OFN639_n_4669), .o(TIMEBOOST_net_21682) );
na03m02 TIMEBOOST_cell_72512 ( .a(TIMEBOOST_net_21372), .b(g65377_sb), .c(TIMEBOOST_net_21646), .o(TIMEBOOST_net_17402) );
in01f01 g63049_u0 ( .a(FE_OFN1129_g64577_p), .o(g63049_sb) );
na02f02 TIMEBOOST_cell_49158 ( .a(TIMEBOOST_net_14796), .b(g61882_sb), .o(n_8066) );
in01m01 g63050_u0 ( .a(FE_OFN1112_g64577_p), .o(g63050_sb) );
na04f04 TIMEBOOST_cell_67919 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q), .b(FE_OFN2081_n_8176), .c(g61950_sb), .d(n_1564), .o(n_7925) );
na03s01 TIMEBOOST_cell_42110 ( .a(g57992_sb), .b(FE_OFN268_n_9880), .c(g57992_db), .o(n_9804) );
na02s01 TIMEBOOST_cell_38522 ( .a(g58198_sb), .b(FE_OFN207_n_9865), .o(TIMEBOOST_net_10873) );
in01f08 g63051_u0 ( .a(FE_OFN1134_g64577_p), .o(g63051_sb) );
na02s02 TIMEBOOST_cell_38524 ( .a(g58000_sb), .b(FE_OFN241_n_9830), .o(TIMEBOOST_net_10874) );
na02s02 TIMEBOOST_cell_38526 ( .a(FE_OFN215_n_9856), .b(g58204_sb), .o(TIMEBOOST_net_10875) );
in01m01 g63052_u0 ( .a(FE_OFN881_g64577_p), .o(g63052_sb) );
na02s02 TIMEBOOST_cell_68283 ( .a(TIMEBOOST_net_21349), .b(TIMEBOOST_net_14158), .o(n_2205) );
na03s02 TIMEBOOST_cell_64900 ( .a(TIMEBOOST_net_14135), .b(g65717_db), .c(TIMEBOOST_net_14520), .o(n_8193) );
na03f02 TIMEBOOST_cell_65163 ( .a(TIMEBOOST_net_14428), .b(g64161_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q), .o(TIMEBOOST_net_15059) );
in01f02 g63053_u0 ( .a(FE_OFN1135_g64577_p), .o(g63053_sb) );
na03f04 TIMEBOOST_cell_46017 ( .a(parchk_pci_cbe_out_in_1202), .b(parchk_pci_cbe_en_in), .c(g67045_da), .o(n_1847) );
na02m02 TIMEBOOST_cell_69808 ( .a(g65035_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q), .o(TIMEBOOST_net_22112) );
in01f01 g63054_u0 ( .a(FE_OFN1128_g64577_p), .o(g63054_sb) );
na04f04 TIMEBOOST_cell_73322 ( .a(n_4047), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q), .c(FE_OFN1124_g64577_p), .d(g62751_sb), .o(n_5478) );
na02s01 TIMEBOOST_cell_38528 ( .a(g58162_sb), .b(FE_OFN241_n_9830), .o(TIMEBOOST_net_10876) );
in01f01 g63055_u0 ( .a(FE_OFN1115_g64577_p), .o(g63055_sb) );
na03f02 TIMEBOOST_cell_72488 ( .a(n_3783), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q), .c(TIMEBOOST_net_21554), .o(TIMEBOOST_net_13235) );
na03m02 TIMEBOOST_cell_72514 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q), .b(TIMEBOOST_net_13881), .c(FE_OFN2109_n_2047), .o(TIMEBOOST_net_21951) );
na04m02 TIMEBOOST_cell_67412 ( .a(TIMEBOOST_net_17241), .b(g65360_sb), .c(FE_OFN1678_n_4655), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q), .o(TIMEBOOST_net_17127) );
in01s01 g63056_u0 ( .a(FE_OFN1104_g64577_p), .o(g63056_sb) );
in01f02 g63058_u0 ( .a(FE_OFN1104_g64577_p), .o(g63058_sb) );
na02s04 TIMEBOOST_cell_72220 ( .a(conf_wb_err_addr_in_961), .b(configuration_wb_err_addr_552), .o(TIMEBOOST_net_23318) );
in01m01 g63059_u0 ( .a(FE_OFN882_g64577_p), .o(g63059_sb) );
na02m01 TIMEBOOST_cell_62431 ( .a(TIMEBOOST_net_20162), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q), .o(TIMEBOOST_net_12307) );
in01m01 g63060_u0 ( .a(FE_OFN877_g64577_p), .o(g63060_sb) );
na02f02 TIMEBOOST_cell_49924 ( .a(TIMEBOOST_net_15179), .b(g63041_sb), .o(n_5168) );
na04f02 TIMEBOOST_cell_72620 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q), .b(FE_OFN1010_n_4734), .c(TIMEBOOST_net_14420), .d(g64146_sb), .o(TIMEBOOST_net_9971) );
na02s01 g58434_u2 ( .a(FE_OFN270_n_9836), .b(FE_OFN1650_n_9428), .o(g58434_db) );
in01f02 g63061_u0 ( .a(FE_OFN1140_g64577_p), .o(g63061_sb) );
in01f02 g63062_u0 ( .a(FE_OFN1122_g64577_p), .o(g63062_sb) );
in01f01 g63063_u0 ( .a(FE_OFN1122_g64577_p), .o(g63063_sb) );
na03f02 TIMEBOOST_cell_72970 ( .a(TIMEBOOST_net_21525), .b(TIMEBOOST_net_10432), .c(FE_OFN1232_n_6391), .o(TIMEBOOST_net_22807) );
na02f01 g63063_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q), .b(FE_OFN1106_g64577_p), .o(g63063_db) );
na02s01 g58421_u2 ( .a(FE_OFN260_n_9860), .b(FE_OFN523_n_9428), .o(g58421_db) );
in01f02 g63064_u0 ( .a(FE_OFN1135_g64577_p), .o(g63064_sb) );
na02s01 TIMEBOOST_cell_43188 ( .a(TIMEBOOST_net_12488), .b(g58176_db), .o(n_9613) );
na03f06 TIMEBOOST_cell_73251 ( .a(TIMEBOOST_net_16960), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .c(g52635_sb), .o(TIMEBOOST_net_5686) );
in01f02 g63065_u0 ( .a(FE_OFN1140_g64577_p), .o(g63065_sb) );
na02m02 TIMEBOOST_cell_38031 ( .a(TIMEBOOST_net_10627), .b(g58182_sb), .o(n_9060) );
na02f02 TIMEBOOST_cell_39435 ( .a(TIMEBOOST_net_11329), .b(g63073_sb), .o(n_5104) );
na02m01 TIMEBOOST_cell_69526 ( .a(n_4447), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q), .o(TIMEBOOST_net_21971) );
in01f02 g63066_u0 ( .a(FE_OFN2105_g64577_p), .o(g63066_sb) );
na03f02 TIMEBOOST_cell_67999 ( .a(TIMEBOOST_net_20617), .b(FE_OFN1248_n_4093), .c(g62929_sb), .o(n_6023) );
in01m01 g63067_u0 ( .a(FE_OFN877_g64577_p), .o(g63067_sb) );
na02f01 TIMEBOOST_cell_49682 ( .a(TIMEBOOST_net_15058), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_13145) );
na02s01 TIMEBOOST_cell_47632 ( .a(TIMEBOOST_net_14033), .b(TIMEBOOST_net_9650), .o(TIMEBOOST_net_12838) );
na02f02 TIMEBOOST_cell_39953 ( .a(TIMEBOOST_net_11588), .b(g62411_sb), .o(n_6776) );
in01f01 g63068_u0 ( .a(FE_OFN1123_g64577_p), .o(g63068_sb) );
no03f06 TIMEBOOST_cell_73342 ( .a(n_4145), .b(n_12595), .c(n_4807), .o(g60339_p) );
na02s01 TIMEBOOST_cell_47881 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q), .b(FE_OFN938_n_2292), .o(TIMEBOOST_net_14158) );
in01f01 g63069_u0 ( .a(FE_OFN1137_g64577_p), .o(g63069_sb) );
na02s01 TIMEBOOST_cell_38423 ( .a(TIMEBOOST_net_10823), .b(g57981_db), .o(n_9818) );
in01m01 g63070_u0 ( .a(FE_OFN882_g64577_p), .o(g63070_sb) );
na03f02 TIMEBOOST_cell_73725 ( .a(FE_OFN1559_n_12042), .b(TIMEBOOST_net_13631), .c(FE_OFN1577_n_12028), .o(n_12659) );
na04f04 TIMEBOOST_cell_67680 ( .a(TIMEBOOST_net_21071), .b(g52400_db), .c(TIMEBOOST_net_13206), .d(g52400_sb), .o(n_14819) );
in01f01 g63071_u0 ( .a(FE_OFN1131_g64577_p), .o(g63071_sb) );
na02m08 TIMEBOOST_cell_45539 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q), .o(TIMEBOOST_net_13664) );
na03f02 TIMEBOOST_cell_73517 ( .a(TIMEBOOST_net_13373), .b(n_6431), .c(g63186_sb), .o(n_5780) );
na02f02 TIMEBOOST_cell_49382 ( .a(TIMEBOOST_net_14908), .b(FE_RN_437_0), .o(TIMEBOOST_net_451) );
in01f01 g63072_u0 ( .a(FE_OFN1121_g64577_p), .o(g63072_sb) );
na03m02 TIMEBOOST_cell_68896 ( .a(n_4498), .b(g64933_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q), .o(TIMEBOOST_net_21656) );
na02m02 TIMEBOOST_cell_63011 ( .a(TIMEBOOST_net_20452), .b(g58090_db), .o(TIMEBOOST_net_9505) );
in01f02 g63073_u0 ( .a(FE_OFN1116_g64577_p), .o(g63073_sb) );
in01f01 g63074_u0 ( .a(FE_OFN1136_g64577_p), .o(g63074_sb) );
na02s06 TIMEBOOST_cell_17922 ( .a(TIMEBOOST_net_5324), .b(n_1690), .o(TIMEBOOST_net_187) );
na03f02 TIMEBOOST_cell_34816 ( .a(TIMEBOOST_net_9443), .b(FE_OFN1421_n_8567), .c(g57491_sb), .o(n_11245) );
in01m01 g63075_u0 ( .a(FE_OFN1129_g64577_p), .o(g63075_sb) );
na02m02 TIMEBOOST_cell_38066 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q), .b(g58401_sb), .o(TIMEBOOST_net_10645) );
na02s01 TIMEBOOST_cell_48183 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q), .b(pci_target_unit_fifos_pcir_control_in_192), .o(TIMEBOOST_net_14309) );
na02m01 TIMEBOOST_cell_48187 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q), .b(pci_target_unit_fifos_pcir_data_in_184), .o(TIMEBOOST_net_14311) );
in01f01 g63076_u0 ( .a(FE_OFN1130_g64577_p), .o(g63076_sb) );
na02m01 TIMEBOOST_cell_52433 ( .a(configuration_pci_err_data_515), .b(wbm_dat_o_14_), .o(TIMEBOOST_net_16434) );
in01m01 g63077_u0 ( .a(FE_OFN1097_g64577_p), .o(g63077_sb) );
na03f06 TIMEBOOST_cell_66262 ( .a(TIMEBOOST_net_15270), .b(n_3290), .c(n_3039), .o(TIMEBOOST_net_8003) );
na02s01 TIMEBOOST_cell_45451 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q), .o(TIMEBOOST_net_13620) );
na02s01 TIMEBOOST_cell_52603 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q), .o(TIMEBOOST_net_16519) );
in01f01 g63078_u0 ( .a(FE_OFN1133_g64577_p), .o(g63078_sb) );
na02s01 TIMEBOOST_cell_63217 ( .a(TIMEBOOST_net_20555), .b(FE_OFN563_n_9895), .o(TIMEBOOST_net_14586) );
na02f02 TIMEBOOST_cell_71016 ( .a(TIMEBOOST_net_17491), .b(FE_OFN1269_n_4095), .o(TIMEBOOST_net_22716) );
in01m02 g63079_u0 ( .a(FE_OFN1132_g64577_p), .o(g63079_sb) );
na03f02 TIMEBOOST_cell_66812 ( .a(TIMEBOOST_net_16845), .b(FE_OFN1345_n_8567), .c(g57140_sb), .o(n_11609) );
in01f02 g63080_u0 ( .a(FE_OFN1119_g64577_p), .o(g63080_sb) );
na02s01 TIMEBOOST_cell_45107 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_), .o(TIMEBOOST_net_13448) );
na03f02 TIMEBOOST_cell_66732 ( .a(TIMEBOOST_net_16828), .b(FE_OFN1305_n_13124), .c(g54366_sb), .o(n_13076) );
na03f01 TIMEBOOST_cell_72426 ( .a(TIMEBOOST_net_14008), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q), .c(wbu_addr_in_261), .o(n_9126) );
in01f01 g63081_u0 ( .a(FE_OFN2106_g64577_p), .o(g63081_sb) );
na03f06 TIMEBOOST_cell_73252 ( .a(TIMEBOOST_net_20409), .b(FE_OFN2076_FE_OCPUNCON1952_FE_OFN697_n_16760), .c(g52632_sb), .o(TIMEBOOST_net_5685) );
in01m01 g63082_u0 ( .a(FE_OFN1133_g64577_p), .o(g63082_sb) );
na03f10 TIMEBOOST_cell_33773 ( .a(n_16521), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q), .c(FE_OCPN1823_n_16560), .o(n_16442) );
na02m02 TIMEBOOST_cell_68285 ( .a(TIMEBOOST_net_21350), .b(g65685_sb), .o(n_2210) );
na03f02 TIMEBOOST_cell_67921 ( .a(TIMEBOOST_net_9970), .b(FE_OFN1100_g64577_p), .c(g62807_sb), .o(n_5366) );
in01f01 g63083_u0 ( .a(FE_OFN1120_g64577_p), .o(g63083_sb) );
no04f04 TIMEBOOST_cell_72578 ( .a(TIMEBOOST_net_14103), .b(wishbone_slave_unit_pcim_if_del_we_in), .c(n_1827), .d(TIMEBOOST_net_594), .o(g61618_p) );
in01f01 g63084_u0 ( .a(FE_OFN1123_g64577_p), .o(g63084_sb) );
na02s01 TIMEBOOST_cell_48821 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q), .o(TIMEBOOST_net_14628) );
in01s01 g63085_u0 ( .a(FE_OFN881_g64577_p), .o(g63085_sb) );
in01m01 TIMEBOOST_cell_67781 ( .a(pci_target_unit_fifos_pcir_data_in_163), .o(TIMEBOOST_net_21208) );
na03m02 TIMEBOOST_cell_70000 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q), .b(FE_OFN2081_n_8176), .c(n_1589), .o(TIMEBOOST_net_22208) );
na02s01 TIMEBOOST_cell_52605 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q), .o(TIMEBOOST_net_16520) );
in01f01 g63086_u0 ( .a(FE_OFN1094_g64577_p), .o(g63086_sb) );
na02f01 TIMEBOOST_cell_69374 ( .a(wbu_latency_tim_val_in_244), .b(n_6986), .o(TIMEBOOST_net_21895) );
na02f01 g63086_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q), .b(FE_OFN1094_g64577_p), .o(g63086_db) );
in01f01 g63087_u0 ( .a(FE_OFN1123_g64577_p), .o(g63087_sb) );
na03f02 TIMEBOOST_cell_73400 ( .a(TIMEBOOST_net_16745), .b(FE_OFN1185_n_3476), .c(g60642_sb), .o(n_5687) );
na03m01 TIMEBOOST_cell_72438 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q), .b(FE_OFN936_n_2292), .c(TIMEBOOST_net_21167), .o(TIMEBOOST_net_21344) );
na02m02 TIMEBOOST_cell_49768 ( .a(TIMEBOOST_net_15101), .b(g61725_sb), .o(n_8371) );
in01m01 g63088_u0 ( .a(FE_OFN1137_g64577_p), .o(g63088_sb) );
na02f01 TIMEBOOST_cell_49684 ( .a(TIMEBOOST_net_15059), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_13161) );
na02f04 TIMEBOOST_cell_26218 ( .a(TIMEBOOST_net_7213), .b(n_7040), .o(FE_RN_267_0) );
na03m02 TIMEBOOST_cell_72690 ( .a(TIMEBOOST_net_21526), .b(g64793_sb), .c(TIMEBOOST_net_21783), .o(TIMEBOOST_net_17129) );
in01m01 g63089_u0 ( .a(FE_OFN1104_g64577_p), .o(g63089_sb) );
na04f04 TIMEBOOST_cell_67706 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q), .b(n_12369), .c(FE_OFN1559_n_12042), .d(n_12238), .o(TIMEBOOST_net_16064) );
na02m10 TIMEBOOST_cell_52435 ( .a(configuration_pci_err_data_516), .b(wbm_dat_o_15_), .o(TIMEBOOST_net_16435) );
in01f04 g63090_u0 ( .a(FE_OFN1131_g64577_p), .o(g63090_sb) );
na03f02 TIMEBOOST_cell_41755 ( .a(TIMEBOOST_net_10571), .b(g64182_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q), .o(TIMEBOOST_net_8325) );
na03f02 TIMEBOOST_cell_72428 ( .a(n_2308), .b(n_3108), .c(n_4743), .o(TIMEBOOST_net_365) );
in01m01 g63091_u0 ( .a(FE_OFN1104_g64577_p), .o(g63091_sb) );
na03f02 TIMEBOOST_cell_73401 ( .a(TIMEBOOST_net_8837), .b(FE_OFN1183_n_3476), .c(g60673_sb), .o(n_5646) );
na02m10 TIMEBOOST_cell_45785 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q), .o(TIMEBOOST_net_13787) );
na02f01 g60664_u2 ( .a(configuration_pci_err_data_504), .b(FE_OFN1183_n_3476), .o(g60664_db) );
in01f01 g63092_u0 ( .a(FE_OFN2106_g64577_p), .o(g63092_sb) );
na02f02 TIMEBOOST_cell_52432 ( .a(TIMEBOOST_net_16433), .b(n_13814), .o(n_14073) );
na03f02 TIMEBOOST_cell_65965 ( .a(n_3963), .b(g62852_sb), .c(g62852_db), .o(n_5265) );
na02s01 TIMEBOOST_cell_45327 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q), .o(TIMEBOOST_net_13558) );
in01f02 g63093_u0 ( .a(FE_OFN1119_g64577_p), .o(g63093_sb) );
na02f02 TIMEBOOST_cell_69373 ( .a(TIMEBOOST_net_21894), .b(g60674_sb), .o(TIMEBOOST_net_5477) );
na03f01 TIMEBOOST_cell_72429 ( .a(TIMEBOOST_net_10179), .b(FE_OFN945_n_2248), .c(g65857_sb), .o(n_1648) );
na03f02 TIMEBOOST_cell_73785 ( .a(TIMEBOOST_net_13752), .b(FE_OFN1601_n_13995), .c(FE_OFN1605_n_13997), .o(n_14512) );
in01f02 g63094_u0 ( .a(FE_OFN1200_n_4090), .o(g63094_sb) );
na03f02 TIMEBOOST_cell_66204 ( .a(TIMEBOOST_net_17553), .b(FE_OFN1284_n_4097), .c(g62357_sb), .o(n_6885) );
in01m01 g63095_u0 ( .a(FE_OFN1106_g64577_p), .o(g63095_sb) );
in01s02 TIMEBOOST_cell_45931 ( .a(TIMEBOOST_net_13949), .o(TIMEBOOST_net_13892) );
na02f01 g63095_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q), .b(FE_OFN1106_g64577_p), .o(g63095_db) );
in01m01 g63096_u0 ( .a(FE_OFN881_g64577_p), .o(g63096_sb) );
na02m04 TIMEBOOST_cell_42822 ( .a(TIMEBOOST_net_12305), .b(g58786_sb), .o(n_9876) );
na03f02 TIMEBOOST_cell_73701 ( .a(TIMEBOOST_net_13517), .b(FE_OFN1762_n_10780), .c(FE_OFN1583_n_12306), .o(n_12763) );
in01m01 g63097_u0 ( .a(FE_OFN1134_g64577_p), .o(g63097_sb) );
na02f08 TIMEBOOST_cell_45108 ( .a(TIMEBOOST_net_13448), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_11821) );
na02m02 TIMEBOOST_cell_68620 ( .a(pci_target_unit_fifos_pciw_addr_data_in_144), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q), .o(TIMEBOOST_net_21518) );
in01m02 g63098_u0 ( .a(FE_OFN1135_g64577_p), .o(g63098_sb) );
na02m02 TIMEBOOST_cell_43851 ( .a(g65363_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_12820) );
na02m02 TIMEBOOST_cell_49670 ( .a(TIMEBOOST_net_15052), .b(g61827_sb), .o(n_8132) );
na02m01 TIMEBOOST_cell_47991 ( .a(n_3747), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q), .o(TIMEBOOST_net_14213) );
in01f01 g63099_u0 ( .a(FE_OFN2106_g64577_p), .o(g63099_sb) );
na02f02 TIMEBOOST_cell_30453 ( .a(n_9009), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q), .o(TIMEBOOST_net_9331) );
in01f02 g63100_u0 ( .a(FE_OFN877_g64577_p), .o(g63100_sb) );
na02s02 TIMEBOOST_cell_48829 ( .a(g57942_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q), .o(TIMEBOOST_net_14632) );
na04m04 TIMEBOOST_cell_73060 ( .a(n_1581), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q), .c(FE_OFN710_n_8232), .d(g61946_sb), .o(n_7933) );
na02m02 TIMEBOOST_cell_71136 ( .a(n_1594), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q), .o(TIMEBOOST_net_22776) );
in01f02 g63101_u0 ( .a(FE_OFN1139_g64577_p), .o(g63101_sb) );
na02f01 g63101_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q), .b(FE_OFN1107_g64577_p), .o(g63101_db) );
na03m02 TIMEBOOST_cell_66089 ( .a(TIMEBOOST_net_20935), .b(FE_OFN1655_n_9502), .c(g58310_sb), .o(n_9026) );
in01m01 g63102_u0 ( .a(FE_OFN1123_g64577_p), .o(g63102_sb) );
na03s01 TIMEBOOST_cell_72363 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_96), .b(wishbone_slave_unit_pci_initiator_if_data_source), .c(g54160_sb), .o(TIMEBOOST_net_13984) );
na03f02 TIMEBOOST_cell_65364 ( .a(TIMEBOOST_net_8277), .b(n_5633), .c(g62094_sb), .o(n_5611) );
in01f02 g63103_u0 ( .a(FE_OFN2104_g64577_p), .o(g63103_sb) );
in01f02 g63104_u0 ( .a(FE_OFN1140_g64577_p), .o(g63104_sb) );
na02f02 TIMEBOOST_cell_50528 ( .a(TIMEBOOST_net_15481), .b(g62488_sb), .o(n_6610) );
na02m02 TIMEBOOST_cell_71398 ( .a(n_1859), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q), .o(TIMEBOOST_net_22907) );
in01s02 g63105_u0 ( .a(FE_OFN2105_g64577_p), .o(g63105_sb) );
na04f02 TIMEBOOST_cell_67923 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_), .b(FE_OFN1092_g64577_p), .c(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .d(g63572_sb), .o(n_4109) );
na02m01 TIMEBOOST_cell_48075 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q), .o(TIMEBOOST_net_14255) );
in01f02 g63106_u0 ( .a(FE_OFN877_g64577_p), .o(g63106_sb) );
na02f01 TIMEBOOST_cell_70708 ( .a(TIMEBOOST_net_13067), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_22562) );
in01s01 TIMEBOOST_cell_17870 ( .a(TIMEBOOST_net_5281), .o(TIMEBOOST_net_5280) );
in01s01 TIMEBOOST_cell_73985 ( .a(TIMEBOOST_net_23549), .o(TIMEBOOST_net_23550) );
in01f01 g63107_u0 ( .a(FE_OFN1115_g64577_p), .o(g63107_sb) );
na02s01 TIMEBOOST_cell_52743 ( .a(pci_target_unit_pcit_if_strd_addr_in_698), .b(pci_target_unit_del_sync_addr_in_216), .o(TIMEBOOST_net_16589) );
in01f01 g63108_u0 ( .a(FE_OFN1242_n_4092), .o(g63108_sb) );
na02f20 TIMEBOOST_cell_3109 ( .a(TIMEBOOST_net_114), .b(n_15922), .o(n_15927) );
in01m01 g63109_u0 ( .a(FE_OFN1118_g64577_p), .o(g63109_sb) );
na04f04 TIMEBOOST_cell_24182 ( .a(n_9089), .b(g57204_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q), .d(FE_OFN1384_n_8567), .o(n_10443) );
na02m04 TIMEBOOST_cell_17906 ( .a(TIMEBOOST_net_5316), .b(pci_target_unit_wishbone_master_reset_rty_cnt), .o(TIMEBOOST_net_158) );
in01m01 g63110_u0 ( .a(FE_OFN1134_g64577_p), .o(g63110_sb) );
na04f02 TIMEBOOST_cell_72476 ( .a(FE_OFN905_n_4736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q), .c(pci_target_unit_fifos_pciw_addr_data_in_138), .d(g64189_sb), .o(n_3978) );
na02s01 TIMEBOOST_cell_17905 ( .a(n_1280), .b(wbm_rty_i), .o(TIMEBOOST_net_5316) );
in01s01 TIMEBOOST_cell_17886 ( .a(TIMEBOOST_net_5297), .o(TIMEBOOST_net_5296) );
in01f06 g63111_u0 ( .a(FE_OFN1131_g64577_p), .o(g63111_sb) );
na03f02 TIMEBOOST_cell_63488 ( .a(n_12002), .b(FE_OFN1559_n_12042), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q), .o(TIMEBOOST_net_20691) );
na04f04 TIMEBOOST_cell_25007 ( .a(n_9321), .b(n_10985), .c(n_9322), .d(n_10198), .o(n_12162) );
in01s01 TIMEBOOST_cell_17904 ( .a(TIMEBOOST_net_5315), .o(TIMEBOOST_net_5314) );
in01f01 g63112_u0 ( .a(FE_OFN1121_g64577_p), .o(g63112_sb) );
na02f01 TIMEBOOST_cell_70698 ( .a(TIMEBOOST_net_13106), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_22557) );
in01s01 TIMEBOOST_cell_17903 ( .a(TIMEBOOST_net_5314), .o(wbs_sel_i_3_) );
in01s01 TIMEBOOST_cell_17902 ( .a(TIMEBOOST_net_5313), .o(TIMEBOOST_net_5312) );
in01f01 g63113_u0 ( .a(FE_OFN1137_g64577_p), .o(g63113_sb) );
na04f04 TIMEBOOST_cell_36829 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q), .b(FE_OFN1414_n_8567), .c(n_9700), .d(g57123_sb), .o(n_11623) );
in01s01 TIMEBOOST_cell_17901 ( .a(TIMEBOOST_net_5312), .o(wbs_sel_i_2_) );
in01f01 g63114_u0 ( .a(FE_OFN1130_g64577_p), .o(g63114_sb) );
na03m02 TIMEBOOST_cell_72066 ( .a(n_3749), .b(FE_OFN644_n_4677), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q), .o(TIMEBOOST_net_23241) );
in01f01 g63115_u0 ( .a(FE_OFN1137_g64577_p), .o(g63115_sb) );
na02s01 TIMEBOOST_cell_54095 ( .a(TIMEBOOST_net_12624), .b(FE_OFN1043_n_2037), .o(TIMEBOOST_net_17265) );
na04f04 TIMEBOOST_cell_73323 ( .a(n_4046), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q), .c(FE_OFN2106_g64577_p), .d(g62725_sb), .o(n_5531) );
na02f01 TIMEBOOST_cell_52933 ( .a(TIMEBOOST_net_13078), .b(FE_OFN1134_g64577_p), .o(TIMEBOOST_net_16684) );
in01m02 g63116_u0 ( .a(FE_OFN1130_g64577_p), .o(g63116_sb) );
na04f04 TIMEBOOST_cell_68001 ( .a(n_3290), .b(pciu_bar0_in_375), .c(n_3050), .d(n_2842), .o(n_4647) );
in01m01 g63117_u0 ( .a(FE_OFN1095_g64577_p), .o(g63117_sb) );
na03f02 TIMEBOOST_cell_66462 ( .a(TIMEBOOST_net_16775), .b(FE_OFN1317_n_6624), .c(g62451_sb), .o(n_6695) );
na02m01 TIMEBOOST_cell_39180 ( .a(g58078_sb), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_11202) );
in01f01 g63118_u0 ( .a(FE_OFN1136_g64577_p), .o(g63118_sb) );
na02m01 TIMEBOOST_cell_68202 ( .a(FE_OFN276_n_9941), .b(n_135), .o(TIMEBOOST_net_21309) );
na02f01 TIMEBOOST_cell_70910 ( .a(TIMEBOOST_net_16729), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_22663) );
in01f02 g63119_u0 ( .a(FE_OFN1132_g64577_p), .o(g63119_sb) );
na02m08 TIMEBOOST_cell_53017 ( .a(configuration_pci_err_data_513), .b(wbm_dat_o_12_), .o(TIMEBOOST_net_16726) );
na02s01 TIMEBOOST_cell_45329 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q), .o(TIMEBOOST_net_13559) );
in01m02 g63120_u0 ( .a(FE_OFN1119_g64577_p), .o(g63120_sb) );
na02s02 TIMEBOOST_cell_63839 ( .a(TIMEBOOST_net_20905), .b(g58090_sb), .o(TIMEBOOST_net_20452) );
na03f02 TIMEBOOST_cell_35066 ( .a(TIMEBOOST_net_9612), .b(FE_OFN1439_n_9372), .c(g58469_sb), .o(n_8983) );
na03m02 TIMEBOOST_cell_33800 ( .a(n_2197), .b(g61717_sb), .c(g61717_db), .o(n_8391) );
in01f01 g63121_u0 ( .a(FE_OFN1125_g64577_p), .o(g63121_sb) );
na04f02 TIMEBOOST_cell_67588 ( .a(n_14738), .b(n_14839), .c(TIMEBOOST_net_20554), .d(g52451_sb), .o(n_14840) );
in01f01 g63122_u0 ( .a(FE_OFN1112_g64577_p), .o(g63122_sb) );
na04f20 TIMEBOOST_cell_20761 ( .a(g75024_sb), .b(conf_w_addr_in_931), .c(n_16027), .d(conf_w_addr_in), .o(n_16393) );
na03f02 TIMEBOOST_cell_35068 ( .a(TIMEBOOST_net_9594), .b(FE_OFN1440_n_9372), .c(g58480_sb), .o(n_9355) );
na03s02 TIMEBOOST_cell_65303 ( .a(g58055_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q), .c(TIMEBOOST_net_12807), .o(TIMEBOOST_net_9399) );
in01m01 g63123_u0 ( .a(FE_OFN1131_g64577_p), .o(g63123_sb) );
na03m02 TIMEBOOST_cell_73108 ( .a(TIMEBOOST_net_10707), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q), .c(TIMEBOOST_net_8754), .o(TIMEBOOST_net_17467) );
na03f02 TIMEBOOST_cell_35070 ( .a(TIMEBOOST_net_9595), .b(FE_OFN1440_n_9372), .c(g58477_sb), .o(n_8979) );
na03f02 TIMEBOOST_cell_35072 ( .a(TIMEBOOST_net_9611), .b(FE_OFN1440_n_9372), .c(g58472_sb), .o(n_8981) );
in01f01 g63124_u0 ( .a(FE_OFN1106_g64577_p), .o(g63124_sb) );
na02f01 g63124_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q), .b(FE_OFN1106_g64577_p), .o(g63124_db) );
na02m10 TIMEBOOST_cell_52607 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q), .o(TIMEBOOST_net_16521) );
in01m01 g63125_u0 ( .a(FE_OFN1134_g64577_p), .o(g63125_sb) );
na02s02 TIMEBOOST_cell_26051 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q), .b(g65874_sb), .o(TIMEBOOST_net_7130) );
in01m01 g63126_u0 ( .a(FE_OFN1106_g64577_p), .o(g63126_sb) );
na02f01 g63126_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q), .b(FE_OFN1106_g64577_p), .o(g63126_db) );
na02f01 g63127_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q), .b(FE_OFN1107_g64577_p), .o(g63127_db) );
na03f02 TIMEBOOST_cell_66589 ( .a(TIMEBOOST_net_17112), .b(FE_OFN1314_n_6624), .c(g62518_sb), .o(n_6541) );
in01f01 g63128_u0 ( .a(FE_OFN1115_g64577_p), .o(g63128_sb) );
na04f04 TIMEBOOST_cell_67709 ( .a(n_12372), .b(n_12116), .c(n_12243), .d(n_12244), .o(n_12901) );
na03f02 TIMEBOOST_cell_35074 ( .a(TIMEBOOST_net_9587), .b(FE_OFN1436_n_9372), .c(g58475_sb), .o(n_9366) );
na02f02 TIMEBOOST_cell_17992 ( .a(TIMEBOOST_net_5359), .b(g67040_sb), .o(n_1649) );
na02m02 TIMEBOOST_cell_38068 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q), .b(g65318_sb), .o(TIMEBOOST_net_10646) );
na02f02 TIMEBOOST_cell_71484 ( .a(wbm_adr_o_10_), .b(g59123_sb), .o(TIMEBOOST_net_22950) );
in01f02 g63130_u0 ( .a(FE_OFN877_g64577_p), .o(g63130_sb) );
na02s01 TIMEBOOST_cell_48866 ( .a(TIMEBOOST_net_14650), .b(g58159_db), .o(TIMEBOOST_net_9531) );
na02f01 TIMEBOOST_cell_70608 ( .a(TIMEBOOST_net_17320), .b(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_22512) );
na03f02 TIMEBOOST_cell_73253 ( .a(TIMEBOOST_net_23272), .b(g64183_sb), .c(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_22465) );
in01f01 g63131_u0 ( .a(FE_OFN1115_g64577_p), .o(g63131_sb) );
in01s01 TIMEBOOST_cell_73895 ( .a(TIMEBOOST_net_23459), .o(TIMEBOOST_net_23460) );
na03m04 TIMEBOOST_cell_73007 ( .a(FE_OFN1049_n_16657), .b(TIMEBOOST_net_16620), .c(g64137_sb), .o(n_4025) );
in01m01 g63132_u0 ( .a(FE_OFN1118_g64577_p), .o(g63132_sb) );
na03f02 TIMEBOOST_cell_73631 ( .a(TIMEBOOST_net_16816), .b(n_16748), .c(g52648_sb), .o(n_14740) );
in01m01 g63133_u0 ( .a(FE_OFN1131_g64577_p), .o(g63133_sb) );
na02f02 TIMEBOOST_cell_50871 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_4__Q), .b(n_13221), .o(TIMEBOOST_net_15653) );
na04s02 TIMEBOOST_cell_64484 ( .a(TIMEBOOST_net_10231), .b(g65802_sb), .c(g61709_sb), .d(g61709_db), .o(n_8409) );
in01f02 g63134_u0 ( .a(FE_OFN1137_g64577_p), .o(g63134_sb) );
na02s01 TIMEBOOST_cell_70430 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q), .o(TIMEBOOST_net_22423) );
in01s01 TIMEBOOST_cell_45996 ( .a(TIMEBOOST_net_13957), .o(TIMEBOOST_net_13956) );
in01s01 TIMEBOOST_cell_17866 ( .a(TIMEBOOST_net_5277), .o(TIMEBOOST_net_5276) );
in01f02 g63135_u0 ( .a(FE_OFN1137_g64577_p), .o(g63135_sb) );
na02f04 TIMEBOOST_cell_17950 ( .a(TIMEBOOST_net_5338), .b(n_3083), .o(TIMEBOOST_net_154) );
in01f02 g63136_u0 ( .a(FE_OFN2105_g64577_p), .o(g63136_sb) );
na02s01 TIMEBOOST_cell_62544 ( .a(g61705_sb), .b(g61953_db), .o(TIMEBOOST_net_20219) );
na03f02 TIMEBOOST_cell_73807 ( .a(TIMEBOOST_net_16553), .b(FE_OFN1775_n_13800), .c(FE_OFN1769_n_14054), .o(g53239_p) );
in01m01 g63137_u0 ( .a(FE_OFN1120_g64577_p), .o(g63137_sb) );
in01m06 g63138_u0 ( .a(FE_OFN881_g64577_p), .o(g63138_sb) );
in01s01 TIMEBOOST_cell_45985 ( .a(TIMEBOOST_net_13946), .o(TIMEBOOST_net_13851) );
na03s02 TIMEBOOST_cell_68416 ( .a(TIMEBOOST_net_8190), .b(g65860_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_21416) );
in01f01 g63139_u0 ( .a(FE_OFN1125_g64577_p), .o(g63139_sb) );
na02f02 TIMEBOOST_cell_70589 ( .a(TIMEBOOST_net_22502), .b(g63082_sb), .o(n_7119) );
na03f02 TIMEBOOST_cell_73402 ( .a(TIMEBOOST_net_17425), .b(FE_OFN1288_n_4098), .c(g63157_sb), .o(n_5824) );
in01f01 g63140_u0 ( .a(FE_OFN1129_g64577_p), .o(g63140_sb) );
na02s01 TIMEBOOST_cell_43917 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q), .o(TIMEBOOST_net_12853) );
na03s01 TIMEBOOST_cell_64392 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q), .b(FE_OFN602_n_9687), .c(TIMEBOOST_net_17475), .o(TIMEBOOST_net_14666) );
in01m01 g63141_u0 ( .a(FE_OFN881_g64577_p), .o(g63141_sb) );
na02f02 TIMEBOOST_cell_17988 ( .a(TIMEBOOST_net_5357), .b(g67040_sb), .o(n_1277) );
na02f01 g63141_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q), .b(FE_OFN881_g64577_p), .o(g63141_db) );
in01f01 g63142_u0 ( .a(FE_OFN1121_g64577_p), .o(g63142_sb) );
na02m02 TIMEBOOST_cell_52437 ( .a(configuration_pci_err_addr_498), .b(wbm_adr_o_28_), .o(TIMEBOOST_net_16436) );
na03f02 TIMEBOOST_cell_73726 ( .a(FE_OFN1559_n_12042), .b(TIMEBOOST_net_13626), .c(FE_OFN1577_n_12028), .o(n_12603) );
in01f01 g63143_u0 ( .a(FE_OFN1129_g64577_p), .o(g63143_sb) );
no04f08 TIMEBOOST_cell_20883 ( .a(FE_RN_677_0), .b(FE_RN_678_0), .c(n_376), .d(n_2844), .o(TIMEBOOST_net_116) );
na03m02 TIMEBOOST_cell_69420 ( .a(n_4493), .b(g65002_db), .c(n_139), .o(TIMEBOOST_net_21918) );
in01f02 g63144_u0 ( .a(FE_OFN1236_n_6391), .o(g63144_sb) );
na03f02 TIMEBOOST_cell_34818 ( .a(TIMEBOOST_net_9461), .b(FE_OFN1387_n_8567), .c(g57253_sb), .o(n_11502) );
in01s01 TIMEBOOST_cell_67718 ( .a(TIMEBOOST_net_21144), .o(TIMEBOOST_net_21145) );
na02s01 TIMEBOOST_cell_54173 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q), .o(TIMEBOOST_net_17304) );
in01f01 g63145_u0 ( .a(FE_OFN1202_n_4090), .o(g63145_sb) );
na02m04 TIMEBOOST_cell_68958 ( .a(g64764_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_21687) );
na03f02 TIMEBOOST_cell_66208 ( .a(TIMEBOOST_net_20966), .b(FE_OFN369_n_4092), .c(g62506_sb), .o(n_6567) );
in01f02 g63146_u0 ( .a(FE_OFN1197_n_4090), .o(g63146_sb) );
na02s02 TIMEBOOST_cell_63061 ( .a(TIMEBOOST_net_20477), .b(g58214_sb), .o(TIMEBOOST_net_16670) );
no02f02 TIMEBOOST_cell_3113 ( .a(TIMEBOOST_net_116), .b(FE_RN_682_0), .o(FE_RN_683_0) );
in01f01 g63147_u0 ( .a(FE_OFN1214_n_4151), .o(g63147_sb) );
na03f02 TIMEBOOST_cell_73727 ( .a(TIMEBOOST_net_13623), .b(FE_OFN1559_n_12042), .c(FE_OFN1575_n_12028), .o(n_12678) );
no02f06 TIMEBOOST_cell_3115 ( .a(TIMEBOOST_net_117), .b(FE_RN_689_0), .o(FE_RN_691_0) );
na03f02 TIMEBOOST_cell_70776 ( .a(n_740), .b(FE_OFN1698_n_5751), .c(wbm_adr_o_3_), .o(TIMEBOOST_net_22596) );
in01m01 g63148_u0 ( .a(FE_OFN1270_n_4095), .o(g63148_sb) );
na03f02 TIMEBOOST_cell_73728 ( .a(TIMEBOOST_net_13632), .b(FE_OCP_RBN2272_n_10268), .c(FE_OFN1751_n_12086), .o(n_12674) );
no02f02 TIMEBOOST_cell_3119 ( .a(TIMEBOOST_net_119), .b(FE_RN_670_0), .o(FE_RN_675_0) );
in01m01 g63149_u0 ( .a(FE_OFN1203_n_4090), .o(g63149_sb) );
na03m02 TIMEBOOST_cell_73109 ( .a(TIMEBOOST_net_22048), .b(g65361_sb), .c(TIMEBOOST_net_22170), .o(TIMEBOOST_net_20949) );
in01s01 TIMEBOOST_cell_63582 ( .a(pciu_cache_lsize_not_zero_in), .o(TIMEBOOST_net_20762) );
na02s01 TIMEBOOST_cell_43827 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q), .b(FE_OFN211_n_9858), .o(TIMEBOOST_net_12808) );
in01m01 g63150_u0 ( .a(FE_OFN1216_n_4151), .o(g63150_sb) );
na02f04 TIMEBOOST_cell_70141 ( .a(TIMEBOOST_net_22278), .b(g64125_sb), .o(n_4037) );
na02m01 TIMEBOOST_cell_68812 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q), .b(FE_OFN659_n_4392), .o(TIMEBOOST_net_21614) );
na02s01 TIMEBOOST_cell_30481 ( .a(n_9642), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q), .o(TIMEBOOST_net_9345) );
in01f01 g63151_u0 ( .a(FE_OFN1276_n_4096), .o(g63151_sb) );
na02f02 TIMEBOOST_cell_50604 ( .a(TIMEBOOST_net_15519), .b(g63171_sb), .o(n_5800) );
na02f08 TIMEBOOST_cell_3123 ( .a(TIMEBOOST_net_121), .b(n_2238), .o(n_2954) );
na02f04 TIMEBOOST_cell_3124 ( .a(n_1362), .b(wbu_addr_in_251), .o(TIMEBOOST_net_122) );
in01f01 g63152_u0 ( .a(FE_OFN2104_g64577_p), .o(g63152_sb) );
in01s01 TIMEBOOST_cell_67711 ( .a(pci_target_unit_fifos_pcir_data_in_187), .o(TIMEBOOST_net_21138) );
in01m01 g63153_u0 ( .a(FE_OFN1215_n_4151), .o(g63153_sb) );
na03f02 TIMEBOOST_cell_72212 ( .a(TIMEBOOST_net_11095), .b(FE_OFN1151_n_13249), .c(TIMEBOOST_net_20893), .o(TIMEBOOST_net_23314) );
na02f06 TIMEBOOST_cell_3125 ( .a(TIMEBOOST_net_122), .b(n_2244), .o(n_2716) );
na02f06 TIMEBOOST_cell_3126 ( .a(n_2243), .b(n_2225), .o(TIMEBOOST_net_123) );
in01f01 g63154_u0 ( .a(FE_OFN1192_n_6935), .o(g63154_sb) );
na02s01 TIMEBOOST_cell_70388 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q), .o(TIMEBOOST_net_22402) );
na02f02 g63154_u2 ( .a(n_3568), .b(FE_OFN1192_n_6935), .o(g63154_db) );
in01f02 g63155_u0 ( .a(FE_OFN1233_n_6391), .o(g63155_sb) );
na03f02 TIMEBOOST_cell_34820 ( .a(TIMEBOOST_net_9358), .b(FE_OFN1421_n_8567), .c(g57480_sb), .o(n_11256) );
na03f02 TIMEBOOST_cell_72238 ( .a(n_3838), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q), .c(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_23327) );
in01f01 g63156_u0 ( .a(FE_OFN1272_n_4096), .o(g63156_sb) );
na02s01 TIMEBOOST_cell_45575 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q), .o(TIMEBOOST_net_13682) );
na02f06 TIMEBOOST_cell_3127 ( .a(TIMEBOOST_net_123), .b(n_2244), .o(n_2712) );
in01f02 g63157_u0 ( .a(FE_OFN1288_n_4098), .o(g63157_sb) );
na02m10 TIMEBOOST_cell_52439 ( .a(configuration_pci_err_addr_490), .b(wbm_adr_o_20_), .o(TIMEBOOST_net_16437) );
na02f01 TIMEBOOST_cell_3129 ( .a(n_2238), .b(TIMEBOOST_net_124), .o(n_2714) );
na02s01 TIMEBOOST_cell_63220 ( .a(FE_OFN601_n_9687), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_20557) );
in01f01 g63158_u0 ( .a(FE_OFN1243_n_4092), .o(g63158_sb) );
na02m01 TIMEBOOST_cell_3131 ( .a(TIMEBOOST_net_125), .b(n_2708), .o(n_2709) );
na03m02 TIMEBOOST_cell_73254 ( .a(TIMEBOOST_net_8781), .b(FE_OFN719_n_8060), .c(g62023_sb), .o(n_7851) );
in01f02 g63159_u0 ( .a(FE_OFN1316_n_6624), .o(g63159_sb) );
na02m02 TIMEBOOST_cell_70153 ( .a(TIMEBOOST_net_22284), .b(g65251_sb), .o(n_3591) );
in01f04 g63160_u0 ( .a(FE_OFN1313_n_6624), .o(g63160_sb) );
na02f01 TIMEBOOST_cell_49686 ( .a(TIMEBOOST_net_15060), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_13162) );
na02f02 TIMEBOOST_cell_70092 ( .a(g65338_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q), .o(TIMEBOOST_net_22254) );
na02s01 TIMEBOOST_cell_38043 ( .a(TIMEBOOST_net_10633), .b(g57960_db), .o(n_9123) );
in01f02 g63161_u0 ( .a(FE_OFN1317_n_6624), .o(g63161_sb) );
na02s01 TIMEBOOST_cell_45331 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q), .o(TIMEBOOST_net_13560) );
in01s01 TIMEBOOST_cell_67713 ( .a(pci_target_unit_fifos_pcir_data_in_167), .o(TIMEBOOST_net_21140) );
na02f02 TIMEBOOST_cell_70097 ( .a(TIMEBOOST_net_22256), .b(FE_OFN1092_g64577_p), .o(TIMEBOOST_net_15151) );
in01m01 g63162_u0 ( .a(FE_OFN1242_n_4092), .o(g63162_sb) );
na02f04 TIMEBOOST_cell_3133 ( .a(TIMEBOOST_net_126), .b(n_1630), .o(n_1994) );
in01f02 g63163_u0 ( .a(FE_OFN1279_n_4097), .o(g63163_sb) );
na02m10 TIMEBOOST_cell_52441 ( .a(configuration_pci_err_data_510), .b(wbm_dat_o_9_), .o(TIMEBOOST_net_16438) );
no02f02 TIMEBOOST_cell_31850 ( .a(TIMEBOOST_net_10029), .b(n_13348), .o(g53084_p) );
in01m01 g63164_u0 ( .a(FE_OFN1225_n_6391), .o(g63164_sb) );
in01m01 g63165_u0 ( .a(FE_OFN881_g64577_p), .o(g63165_sb) );
na02f20 TIMEBOOST_cell_17975 ( .a(n_15923), .b(n_2016), .o(TIMEBOOST_net_5351) );
in01s02 TIMEBOOST_cell_45967 ( .a(pci_target_unit_fifos_pcir_data_in_162), .o(TIMEBOOST_net_13928) );
in01m01 g63166_u0 ( .a(FE_OFN1295_n_4098), .o(g63166_sb) );
na02m08 TIMEBOOST_cell_52745 ( .a(pci_target_unit_pcit_if_strd_addr_in_687), .b(n_2515), .o(TIMEBOOST_net_16590) );
na03f02 TIMEBOOST_cell_66185 ( .a(TIMEBOOST_net_16435), .b(FE_OFN1179_n_3476), .c(g60646_sb), .o(n_5681) );
na04f04 TIMEBOOST_cell_42515 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_776), .c(FE_OFN2134_n_13124), .d(g54340_sb), .o(n_12976) );
in01f01 g63167_u0 ( .a(FE_OFN1276_n_4096), .o(g63167_sb) );
na02s01 TIMEBOOST_cell_45573 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q), .o(TIMEBOOST_net_13681) );
na02m02 TIMEBOOST_cell_64004 ( .a(wbm_adr_o_22_), .b(g58800_sb), .o(TIMEBOOST_net_20988) );
na02m02 TIMEBOOST_cell_64038 ( .a(n_1960), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q), .o(TIMEBOOST_net_21005) );
in01m01 g63168_u0 ( .a(FE_OFN1242_n_4092), .o(g63168_sb) );
na02f02 g59797_u2 ( .a(n_3472), .b(FE_OFN1698_n_5751), .o(g59797_db) );
na02f02 TIMEBOOST_cell_50374 ( .a(TIMEBOOST_net_15404), .b(g62609_sb), .o(n_6335) );
na02m06 TIMEBOOST_cell_68825 ( .a(TIMEBOOST_net_21620), .b(n_4465), .o(TIMEBOOST_net_10641) );
in01f01 g63169_u0 ( .a(FE_OFN1132_g64577_p), .o(g63169_sb) );
na02m02 TIMEBOOST_cell_30539 ( .a(n_9026), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q), .o(TIMEBOOST_net_9374) );
in01m02 g63170_u0 ( .a(FE_OFN1118_g64577_p), .o(g63170_sb) );
na02m02 TIMEBOOST_cell_68726 ( .a(FE_OFN660_n_4392), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q), .o(TIMEBOOST_net_21571) );
na02f02 TIMEBOOST_cell_69679 ( .a(TIMEBOOST_net_22047), .b(TIMEBOOST_net_14604), .o(TIMEBOOST_net_17116) );
na02m02 TIMEBOOST_cell_39535 ( .a(TIMEBOOST_net_11379), .b(g63137_sb), .o(n_4975) );
in01m01 g63171_u0 ( .a(FE_OFN1225_n_6391), .o(g63171_sb) );
na02f02 TIMEBOOST_cell_63789 ( .a(TIMEBOOST_net_20880), .b(FE_OFN1151_n_13249), .o(TIMEBOOST_net_20430) );
in01f01 g63172_u0 ( .a(FE_OFN1112_g64577_p), .o(g63172_sb) );
na02s01 TIMEBOOST_cell_49385 ( .a(pci_target_unit_del_sync_addr_in_219), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_14910) );
na03s02 TIMEBOOST_cell_67664 ( .a(TIMEBOOST_net_14930), .b(g58068_sb), .c(TIMEBOOST_net_15082), .o(TIMEBOOST_net_9330) );
na03m02 TIMEBOOST_cell_72734 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q), .b(FE_OFN646_n_4497), .c(TIMEBOOST_net_21996), .o(TIMEBOOST_net_17575) );
in01f01 g63173_u0 ( .a(FE_OFN1194_n_6935), .o(g63173_sb) );
na02f02 TIMEBOOST_cell_70541 ( .a(TIMEBOOST_net_22478), .b(g63076_sb), .o(n_5098) );
na02m02 TIMEBOOST_cell_53468 ( .a(TIMEBOOST_net_16951), .b(g62009_sb), .o(n_7877) );
na03f02 TIMEBOOST_cell_42469 ( .a(TIMEBOOST_net_9190), .b(FE_OFN1326_n_13547), .c(g53930_sb), .o(n_13515) );
in01f01 g63174_u0 ( .a(FE_OFN1206_n_6356), .o(g63174_sb) );
na02f02 TIMEBOOST_cell_27185 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_7697) );
na03f02 TIMEBOOST_cell_73403 ( .a(TIMEBOOST_net_17413), .b(FE_OFN1200_n_4090), .c(g62572_sb), .o(n_6410) );
in01f01 g63175_u0 ( .a(FE_OFN1136_g64577_p), .o(g63175_sb) );
na03m04 TIMEBOOST_cell_72825 ( .a(g65428_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q), .c(TIMEBOOST_net_14413), .o(TIMEBOOST_net_13373) );
na02s02 TIMEBOOST_cell_43105 ( .a(FE_OFN223_n_9844), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q), .o(TIMEBOOST_net_12447) );
in01m01 g63176_u0 ( .a(FE_OFN1116_g64577_p), .o(g63176_sb) );
na02f02 TIMEBOOST_cell_50190 ( .a(TIMEBOOST_net_15312), .b(g60640_sb), .o(n_5689) );
na02m02 TIMEBOOST_cell_48915 ( .a(FE_OFN231_n_9839), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q), .o(TIMEBOOST_net_14675) );
na03f02 TIMEBOOST_cell_73632 ( .a(TIMEBOOST_net_23378), .b(FE_OCPN1847_n_14981), .c(g59110_sb), .o(n_8708) );
in01f02 g63177_u0 ( .a(FE_OFN1230_n_6391), .o(g63177_sb) );
na03f02 TIMEBOOST_cell_34822 ( .a(TIMEBOOST_net_9482), .b(FE_OFN1421_n_8567), .c(g57114_sb), .o(n_11632) );
na04f04 TIMEBOOST_cell_68003 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q), .b(g62963_sb), .c(n_4225), .d(FE_OFN1223_n_6391), .o(n_5956) );
na04f04 TIMEBOOST_cell_73663 ( .a(n_4051), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q), .c(FE_OFN1118_g64577_p), .d(g62745_sb), .o(n_5491) );
in01f02 g63178_u0 ( .a(FE_OFN1310_n_6624), .o(g63178_sb) );
na02m01 TIMEBOOST_cell_69262 ( .a(n_4645), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q), .o(TIMEBOOST_net_21839) );
na03f02 TIMEBOOST_cell_66591 ( .a(TIMEBOOST_net_17128), .b(FE_OFN1323_n_6436), .c(g62967_sb), .o(n_5948) );
na02f02 TIMEBOOST_cell_69845 ( .a(TIMEBOOST_net_22130), .b(FE_OFN713_n_8140), .o(TIMEBOOST_net_16370) );
in01m01 g63179_u0 ( .a(FE_OFN1095_g64577_p), .o(g63179_sb) );
na02m01 TIMEBOOST_cell_17986 ( .a(TIMEBOOST_net_5356), .b(g67051_sb), .o(n_1495) );
na02f01 g63179_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q), .b(FE_OFN1095_g64577_p), .o(g63179_db) );
in01m01 g63180_u0 ( .a(FE_OFN1215_n_4151), .o(g63180_sb) );
na03s02 TIMEBOOST_cell_72443 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(FE_OFN946_n_2248), .c(TIMEBOOST_net_21346), .o(n_1573) );
na02f01 TIMEBOOST_cell_62543 ( .a(TIMEBOOST_net_20218), .b(FE_OFN918_n_4725), .o(TIMEBOOST_net_14335) );
na03f02 TIMEBOOST_cell_73404 ( .a(TIMEBOOST_net_21005), .b(FE_OFN1264_n_4095), .c(g62754_sb), .o(n_6129) );
in01f01 g63181_u0 ( .a(FE_OFN1272_n_4096), .o(g63181_sb) );
in01s01 TIMEBOOST_cell_45891 ( .a(TIMEBOOST_net_13852), .o(wbs_adr_i_8_) );
na03f06 TIMEBOOST_cell_64314 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q), .b(n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_389), .o(TIMEBOOST_net_17291) );
na03m02 TIMEBOOST_cell_72843 ( .a(g65297_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q), .c(TIMEBOOST_net_16268), .o(TIMEBOOST_net_20954) );
in01f01 g63182_u0 ( .a(FE_OFN1130_g64577_p), .o(g63182_sb) );
in01s01 TIMEBOOST_cell_73920 ( .a(wbm_dat_i_11_), .o(TIMEBOOST_net_23485) );
na04f04 TIMEBOOST_cell_24815 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q), .b(g58822_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q), .d(FE_OFN2153_n_16439), .o(n_8619) );
in01f01 g63183_u0 ( .a(FE_OFN1194_n_6935), .o(g63183_sb) );
in01m01 TIMEBOOST_cell_45932 ( .a(TIMEBOOST_net_13892), .o(TIMEBOOST_net_13893) );
na02s01 TIMEBOOST_cell_53497 ( .a(FE_OFN258_n_9862), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q), .o(TIMEBOOST_net_16966) );
in01f01 g63184_u0 ( .a(FE_OFN1212_n_4151), .o(g63184_sb) );
na02s01 TIMEBOOST_cell_45345 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q), .o(TIMEBOOST_net_13567) );
na04f02 TIMEBOOST_cell_36825 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q), .b(FE_OFN1394_n_8567), .c(n_8554), .d(g58594_sb), .o(n_8902) );
na03f02 TIMEBOOST_cell_65944 ( .a(TIMEBOOST_net_16404), .b(FE_OFN1163_n_5615), .c(g62099_sb), .o(n_5604) );
in01m01 g63185_u0 ( .a(FE_OFN1203_n_4090), .o(g63185_sb) );
na02s01 TIMEBOOST_cell_3161 ( .a(TIMEBOOST_net_140), .b(g65849_sb), .o(n_1574) );
in01f02 g63186_u0 ( .a(n_6431), .o(g63186_sb) );
na02f08 TIMEBOOST_cell_52937 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_767), .b(FE_RN_578_0), .o(TIMEBOOST_net_16686) );
na02s01 TIMEBOOST_cell_54183 ( .a(configuration_wb_err_addr_559), .b(conf_wb_err_addr_in_968), .o(TIMEBOOST_net_17309) );
in01f01 g63187_u0 ( .a(FE_OFN1285_n_4097), .o(g63187_sb) );
na02m02 TIMEBOOST_cell_69224 ( .a(FE_OFN643_n_4677), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q), .o(TIMEBOOST_net_21820) );
na02f01 TIMEBOOST_cell_63096 ( .a(n_16867), .b(n_4085), .o(TIMEBOOST_net_20495) );
na02s01 TIMEBOOST_cell_45405 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_13597) );
in01f01 g63188_u0 ( .a(FE_OFN1130_g64577_p), .o(g63188_sb) );
na04f04 TIMEBOOST_cell_73405 ( .a(n_4354), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q), .c(FE_OFN1250_n_4093), .d(g62503_sb), .o(n_6575) );
na02f10 TIMEBOOST_cell_17948 ( .a(TIMEBOOST_net_5337), .b(n_15923), .o(TIMEBOOST_net_114) );
na02m08 TIMEBOOST_cell_17949 ( .a(wbs_we_i), .b(n_1347), .o(TIMEBOOST_net_5338) );
in01f02 g63189_u0 ( .a(FE_OFN1269_n_4095), .o(g63189_sb) );
na02m10 TIMEBOOST_cell_53019 ( .a(configuration_pci_err_data_519), .b(wbm_dat_o_18_), .o(TIMEBOOST_net_16727) );
in01f01 g63190_u0 ( .a(FE_OFN1212_n_4151), .o(g63190_sb) );
na02m10 TIMEBOOST_cell_53053 ( .a(configuration_pci_err_data_522), .b(wbm_dat_o_21_), .o(TIMEBOOST_net_16744) );
na02f04 TIMEBOOST_cell_3165 ( .a(TIMEBOOST_net_142), .b(n_2236), .o(n_2948) );
na02f01 TIMEBOOST_cell_18093 ( .a(pci_target_unit_pcit_if_strd_addr_in_709), .b(FE_OFN784_n_2678), .o(TIMEBOOST_net_5410) );
in01f01 g63191_u0 ( .a(FE_OFN1121_g64577_p), .o(g63191_sb) );
na04m10 TIMEBOOST_cell_64339 ( .a(g56933_sb), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q), .c(pci_target_unit_fifos_pcir_flush_in), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q), .o(TIMEBOOST_net_15867) );
na02f06 TIMEBOOST_cell_17947 ( .a(n_15924), .b(n_2078), .o(TIMEBOOST_net_5337) );
na02f02 TIMEBOOST_cell_18212 ( .a(TIMEBOOST_net_5469), .b(n_4660), .o(n_5713) );
in01f01 g63192_u0 ( .a(FE_OFN1202_n_4090), .o(g63192_sb) );
in01s01 TIMEBOOST_cell_63550 ( .a(TIMEBOOST_net_20730), .o(TIMEBOOST_net_10058) );
na03f02 TIMEBOOST_cell_73786 ( .a(TIMEBOOST_net_16536), .b(FE_OFN1599_n_13995), .c(FE_OFN1606_n_13997), .o(g53231_p) );
in01f02 g63193_u0 ( .a(FE_OFN1142_n_15261), .o(g63193_sb) );
na02m10 TIMEBOOST_cell_29003 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q), .o(TIMEBOOST_net_8606) );
na02f04 TIMEBOOST_cell_51026 ( .a(TIMEBOOST_net_15730), .b(n_3413), .o(n_4894) );
in01m01 g63194_u0 ( .a(n_5546), .o(g63194_sb) );
na04f04 TIMEBOOST_cell_24621 ( .a(n_9233), .b(g57059_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q), .d(FE_OFN2182_n_8567), .o(n_10848) );
na04f04 TIMEBOOST_cell_24645 ( .a(n_9686), .b(g57245_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q), .d(FE_OFN2179_n_8567), .o(n_11512) );
in01f02 g63195_u0 ( .a(FE_OFN1142_n_15261), .o(g63195_sb) );
na02m06 TIMEBOOST_cell_45817 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q), .o(TIMEBOOST_net_13803) );
na02f02 TIMEBOOST_cell_69111 ( .a(TIMEBOOST_net_21763), .b(g64160_db), .o(n_4005) );
in01f02 g63196_u0 ( .a(FE_OFN1143_n_15261), .o(g63196_sb) );
in01f01 g63197_u0 ( .a(FE_OFN1192_n_6935), .o(g63197_sb) );
na02f06 TIMEBOOST_cell_3337 ( .a(TIMEBOOST_net_228), .b(n_2424), .o(n_2490) );
in01f01 g63198_u0 ( .a(FE_OFN1192_n_6935), .o(g63198_sb) );
na02m10 TIMEBOOST_cell_45245 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q), .o(TIMEBOOST_net_13517) );
na02f02 g63198_u2 ( .a(n_1199), .b(FE_OFN1192_n_6935), .o(g63198_db) );
na02m02 TIMEBOOST_cell_68704 ( .a(n_3761), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q), .o(TIMEBOOST_net_21560) );
in01f01 g63199_u0 ( .a(FE_OFN1192_n_6935), .o(g63199_sb) );
na02f02 TIMEBOOST_cell_39497 ( .a(TIMEBOOST_net_11360), .b(g62793_sb), .o(n_5402) );
na02f01 g63199_u2 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .b(FE_OFN1192_n_6935), .o(g63199_db) );
na02m02 TIMEBOOST_cell_69264 ( .a(n_4672), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q), .o(TIMEBOOST_net_21840) );
no02f04 g63200_u0 ( .a(wbm_adr_o_16_), .b(n_2442), .o(g63200_p) );
ao12f02 g63200_u1 ( .a(g63200_p), .b(wbm_adr_o_16_), .c(n_2442), .o(n_3152) );
no02f02 g63201_u0 ( .a(wbu_addr_in_265), .b(n_2438), .o(g63201_p) );
ao12f02 g63201_u1 ( .a(g63201_p), .b(wbu_addr_in_265), .c(n_2438), .o(n_3151) );
in01f01 g63202_u0 ( .a(FE_OFN1697_n_5751), .o(g63202_sb) );
na02s01 TIMEBOOST_cell_45453 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q), .o(TIMEBOOST_net_13621) );
na02f02 TIMEBOOST_cell_69191 ( .a(TIMEBOOST_net_21803), .b(g64271_sb), .o(TIMEBOOST_net_14984) );
na04f04 TIMEBOOST_cell_73255 ( .a(n_2154), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q), .c(FE_OFN2212_n_8407), .d(g62014_sb), .o(n_7867) );
in01f01 g63203_u0 ( .a(FE_OFN1697_n_5751), .o(g63203_sb) );
na03f02 TIMEBOOST_cell_46741 ( .a(TIMEBOOST_net_10947), .b(g64237_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q), .o(TIMEBOOST_net_13018) );
in01f02 g63204_u0 ( .a(FE_OFN1700_n_5751), .o(g63204_sb) );
na02s06 TIMEBOOST_cell_47565 ( .a(wbs_dat_i_4_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q), .o(TIMEBOOST_net_14000) );
na02m10 TIMEBOOST_cell_68332 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_5__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_388), .o(TIMEBOOST_net_21374) );
na02f01 TIMEBOOST_cell_64076 ( .a(n_1094), .b(wishbone_slave_unit_fifos_outGreyCount_1_), .o(TIMEBOOST_net_21024) );
no02m02 g63206_u0 ( .a(n_416), .b(n_1659), .o(g63206_p) );
ao12m02 g63206_u1 ( .a(g63206_p), .b(n_416), .c(n_1659), .o(n_2014) );
no02f02 g63207_u0 ( .a(pci_target_unit_fifos_pciw_inTransactionCount_0_), .b(n_5546), .o(g63207_p) );
ao12f01 g63207_u1 ( .a(g63207_p), .b(pci_target_unit_fifos_pciw_inTransactionCount_0_), .c(n_5546), .o(n_4797) );
no02f02 g63208_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_10_), .b(n_2473), .o(g63208_p) );
ao12f01 g63208_u1 ( .a(g63208_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_10_), .c(n_2473), .o(n_2965) );
no02m04 g63209_u0 ( .a(n_207), .b(n_2477), .o(g63209_p) );
ao12m02 g63209_u1 ( .a(g63209_p), .b(n_207), .c(n_2477), .o(n_2964) );
in01f01 g63213_u0 ( .a(FE_OFN191_n_1193), .o(n_2284) );
ao22f40 g63214_u0 ( .a(pci_irdy_i), .b(n_961), .c(parchk_pci_irdy_en_in), .d(out_bckp_irdy_out), .o(n_1193) );
no02f04 g63215_u0 ( .a(n_2254), .b(n_2249), .o(g63215_p) );
ao12f04 g63215_u1 ( .a(g63215_p), .b(n_2254), .c(n_2249), .o(n_2963) );
no02f08 g63216_u0 ( .a(n_2253), .b(n_2251), .o(g63216_p) );
ao12f08 g63216_u1 ( .a(g63216_p), .b(n_2253), .c(n_2251), .o(n_2962) );
no02f04 g63217_u0 ( .a(n_2252), .b(n_2255), .o(g63217_p) );
ao12f08 g63217_u1 ( .a(g63217_p), .b(n_2252), .c(n_2255), .o(n_2961) );
na02s01 g63226_u0 ( .a(n_4795), .b(n_1684), .o(n_4796) );
no02m02 g63227_u0 ( .a(n_2959), .b(n_2412), .o(n_2960) );
in01f01 g63228_u0 ( .a(n_3157), .o(n_2958) );
no02f06 g63229_u0 ( .a(n_15390), .b(n_705), .o(TIMEBOOST_net_10066) );
in01f20 g63230_u0 ( .a(n_4149), .o(n_5592) );
in01f10 g63245_u0 ( .a(n_4149), .o(n_5633) );
no02f20 g63250_u0 ( .a(n_3120), .b(FE_OCPN1838_n_1238), .o(n_4149) );
na02f04 g63251_u0 ( .a(n_3271), .b(n_4743), .o(n_8450) );
na02f10 g63252_u0 ( .a(n_2013), .b(wbu_addr_in_254), .o(g63252_p) );
in01f08 g63252_u1 ( .a(g63252_p), .o(n_2487) );
na02f20 g63253_u0 ( .a(n_2012), .b(wbm_adr_o_5_), .o(g63253_p) );
in01f10 g63253_u1 ( .a(g63253_p), .o(n_2485) );
na02f40 g63254_u0 ( .a(n_1669), .b(conf_wb_err_addr_in_946), .o(n_2035) );
na02f02 g63255_u0 ( .a(FE_OFN2245_n_4792), .b(n_2950), .o(n_4793) );
na02f20 g63256_u0 ( .a(n_2897), .b(n_4743), .o(g63256_p) );
in01f20 g63256_u1 ( .a(g63256_p), .o(n_16916) );
na04f04 TIMEBOOST_cell_73406 ( .a(n_4345), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q), .c(FE_OFN1214_n_4151), .d(g62616_sb), .o(n_6325) );
na03f02 TIMEBOOST_cell_66913 ( .a(FE_OFN1733_n_16317), .b(TIMEBOOST_net_13577), .c(FE_OFN1738_n_11019), .o(n_12722) );
na02f08 g63259_u0 ( .a(n_1438), .b(pci_target_unit_del_sync_comp_cycle_count_3_), .o(g63259_p) );
in01f06 g63259_u1 ( .a(g63259_p), .o(n_1692) );
no02s02 g63261_u0 ( .a(n_1226), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(n_1714) );
na02f20 g63263_u0 ( .a(n_1476), .b(wishbone_slave_unit_del_sync_comp_cycle_count_3_), .o(g63263_p) );
in01f10 g63263_u1 ( .a(g63263_p), .o(n_1694) );
na02f02 g63264_u0 ( .a(n_4939), .b(FE_OFN1192_n_6935), .o(n_7136) );
in01f06 g63265_u0 ( .a(n_2956), .o(n_2957) );
no02f10 g63266_u0 ( .a(n_15390), .b(n_2215), .o(n_2956) );
no02f02 g63267_u0 ( .a(n_15390), .b(n_3267), .o(n_4177) );
na02f02 g63268_u0 ( .a(n_3406), .b(n_5230), .o(g63268_p) );
in01f02 g63268_u1 ( .a(g63268_p), .o(n_4654) );
na02f02 g63269_u0 ( .a(n_3117), .b(n_3245), .o(n_4146) );
na02f01 g63270_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(n_3455) );
no02f10 g63271_u0 ( .a(n_15390), .b(n_2966), .o(g63271_p) );
in01f08 g63271_u1 ( .a(g63271_p), .o(n_3342) );
no02f04 g63272_u0 ( .a(n_8440), .b(n_3388), .o(n_7809) );
na02s01 TIMEBOOST_cell_54515 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q), .o(TIMEBOOST_net_17475) );
no02f10 g63275_u0 ( .a(n_3090), .b(n_8440), .o(n_7803) );
na02s01 g63276_u0 ( .a(n_8440), .b(configuration_interrupt_line_39), .o(n_7565) );
na02s01 g63277_u0 ( .a(n_8440), .b(configuration_interrupt_line_40), .o(n_7564) );
na02s01 g63278_u0 ( .a(n_8440), .b(configuration_interrupt_line_41), .o(n_7562) );
na02s01 TIMEBOOST_cell_52609 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q), .o(TIMEBOOST_net_16522) );
in01f40 g63280_u0 ( .a(n_4685), .o(n_7398) );
in01f40 g63284_u0 ( .a(n_15919), .o(n_4685) );
na02f02 g63287_u0 ( .a(n_3109), .b(n_3247), .o(n_4144) );
na02s01 g63288_u0 ( .a(n_8440), .b(configuration_interrupt_line_43), .o(n_7561) );
na02f08 g63289_u0 ( .a(n_3409), .b(n_16160), .o(n_7321) );
na02s01 TIMEBOOST_cell_48871 ( .a(FE_OFN596_n_9694), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_14653) );
na02f02 g63291_u0 ( .a(n_2920), .b(n_3116), .o(g63291_p) );
in01f02 g63291_u1 ( .a(g63291_p), .o(n_3454) );
na02f10 g63292_u0 ( .a(n_2013), .b(n_964), .o(g63292_p) );
in01f10 g63292_u1 ( .a(g63292_p), .o(n_2680) );
no02m02 g63293_u0 ( .a(n_8440), .b(n_4720), .o(g63293_p) );
in01f02 g63293_u1 ( .a(g63293_p), .o(n_8446) );
na02s01 g63294_u0 ( .a(n_8440), .b(wbu_cache_line_size_in_208), .o(n_7560) );
na03f02 TIMEBOOST_cell_73061 ( .a(TIMEBOOST_net_22039), .b(FE_OFN717_n_8176), .c(g61750_sb), .o(n_8316) );
na02f06 g63297_u0 ( .a(n_2954), .b(wbu_addr_in_273), .o(n_2955) );
na02f04 g63298_u0 ( .a(n_3147), .b(wbu_addr_in_276), .o(n_3148) );
na02f02 TIMEBOOST_cell_18230 ( .a(TIMEBOOST_net_5478), .b(n_4663), .o(n_6987) );
no02f20 g63301_u0 ( .a(n_8440), .b(n_3278), .o(n_7466) );
na03f02 TIMEBOOST_cell_73518 ( .a(TIMEBOOST_net_17484), .b(n_6554), .c(g62919_sb), .o(n_6041) );
na02m02 TIMEBOOST_cell_38072 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q), .b(g65334_sb), .o(TIMEBOOST_net_10648) );
in01f02 g63307_u1 ( .a(g63307_p), .o(n_3450) );
na04f02 TIMEBOOST_cell_72698 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q), .b(FE_OFN660_n_4392), .c(g64930_sb), .d(n_3741), .o(n_3678) );
na02s01 g63309_u0 ( .a(n_8440), .b(wbu_cache_line_size_in_207), .o(n_7559) );
na02f02 g63310_u0 ( .a(n_853), .b(n_5546), .o(n_5545) );
in01s01 g63313_u0 ( .a(n_3448), .o(n_3449) );
no02f08 g63314_u0 ( .a(n_16280), .b(n_3319), .o(n_3448) );
na02f10 g63315_u0 ( .a(FE_OFN1143_n_15261), .b(n_4535), .o(g63315_p) );
in01f10 g63315_u1 ( .a(g63315_p), .o(n_13825) );
na02f04 g63316_u0 ( .a(conf_wb_err_addr_in_943), .b(FE_OFN1142_n_15261), .o(n_3327) );
in01f06 g63318_u0 ( .a(n_2011), .o(n_2458) );
na02s01 TIMEBOOST_cell_47587 ( .a(g58775_sb), .b(n_8831), .o(TIMEBOOST_net_14011) );
no02f01 g63320_u0 ( .a(n_1424), .b(FE_OFN778_n_4152), .o(n_2953) );
no02f01 g63321_u0 ( .a(FE_OCPN1841_n_16089), .b(n_8498), .o(n_2725) );
no02f01 g63322_u0 ( .a(n_2423), .b(FE_OFN778_n_4152), .o(n_2952) );
no02f04 g63323_u0 ( .a(n_1673), .b(FE_OFN1143_n_15261), .o(n_3326) );
ao12f01 g63324_u0 ( .a(n_4536), .b(n_2370), .c(n_4718), .o(n_4936) );
no02f10 g63338_u0 ( .a(n_15054), .b(n_2354), .o(g63338_p) );
in01f08 g63338_u1 ( .a(g63338_p), .o(n_5763) );
na02s01 g63339_u0 ( .a(n_8440), .b(wbu_cache_line_size_in_209), .o(n_7558) );
na02f04 g63340_u0 ( .a(n_2280), .b(FE_OFN199_n_3298), .o(g63340_p) );
in01f02 g63340_u1 ( .a(g63340_p), .o(n_4142) );
na02f04 g63341_u0 ( .a(n_3324), .b(wbm_adr_o_27_), .o(n_3325) );
na02f04 g63342_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_), .b(n_4662), .o(n_3447) );
na02f06 g63343_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_), .o(n_3446) );
na02f06 g63344_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_), .o(n_3445) );
na02s02 TIMEBOOST_cell_48872 ( .a(TIMEBOOST_net_14653), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_12817) );
na02f10 g63348_u0 ( .a(n_2012), .b(n_1116), .o(g63348_p) );
in01f10 g63348_u1 ( .a(g63348_p), .o(n_2738) );
na02f10 g63349_u0 ( .a(n_2950), .b(n_1435), .o(n_2951) );
na02f04 g63350_u0 ( .a(n_2018), .b(pci_target_unit_wishbone_master_rty_counter_7_), .o(n_2019) );
no02f04 g63351_u0 ( .a(n_2395), .b(FE_OFN1142_n_15261), .o(n_3323) );
na02s01 g63352_u0 ( .a(n_8440), .b(wbu_cache_line_size_in_211), .o(n_7557) );
na02f04 g63353_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(n_3444) );
na02m01 g63354_u0 ( .a(n_3020), .b(parity_checker_check_for_serr_on_second), .o(n_7396) );
na02f04 g63355_u0 ( .a(n_2948), .b(wbm_adr_o_24_), .o(n_2949) );
na02m02 g63356_u0 ( .a(n_4662), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_), .o(n_3443) );
in01f02 g63358_u0 ( .a(n_7795), .o(n_7785) );
no02f10 g63359_u0 ( .a(n_8440), .b(n_3261), .o(n_7795) );
na02m02 TIMEBOOST_cell_70213 ( .a(TIMEBOOST_net_22314), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_15049) );
na02s01 g63361_u0 ( .a(wishbone_slave_unit_del_sync_comp_rty_exp_clr), .b(wishbone_slave_unit_del_sync_comp_rty_exp_reg), .o(g63361_p) );
in01s01 g63361_u1 ( .a(g63361_p), .o(n_4140) );
na02f02 g63362_u0 ( .a(n_15733), .b(n_5230), .o(g63362_p) );
in01f02 g63362_u1 ( .a(g63362_p), .o(n_4641) );
na04f06 TIMEBOOST_cell_65975 ( .a(FE_OFN237_n_9118), .b(g58251_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q), .d(g58251_db), .o(TIMEBOOST_net_16841) );
no02m02 g63364_u0 ( .a(n_8440), .b(FE_OFN2100_n_3281), .o(g63364_p) );
in01f02 g63364_u1 ( .a(g63364_p), .o(n_8444) );
na02m02 TIMEBOOST_cell_69708 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q), .b(n_4482), .o(TIMEBOOST_net_22062) );
na02f04 g63373_u0 ( .a(n_2921), .b(n_2625), .o(n_3321) );
ao12f02 g63374_u0 ( .a(n_3111), .b(configuration_wb_err_addr_560), .c(n_15444), .o(n_3440) );
ao12f02 g63375_u0 ( .a(n_3114), .b(configuration_wb_err_addr_562), .c(n_15444), .o(n_3438) );
na02s01 TIMEBOOST_cell_49415 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q), .o(TIMEBOOST_net_14925) );
na02f02 g63377_u0 ( .a(n_3417), .b(n_4637), .o(n_4638) );
in01f02 g63378_u0 ( .a(FE_OFN1117_g64577_p), .o(g63378_sb) );
in01s01 TIMEBOOST_cell_63598 ( .a(TIMEBOOST_net_20778), .o(TIMEBOOST_net_20747) );
na02s02 TIMEBOOST_cell_25482 ( .a(TIMEBOOST_net_5361), .b(TIMEBOOST_net_6845), .o(n_9856) );
in01f02 g63379_u0 ( .a(n_4137), .o(n_4636) );
ao12f04 g63380_u0 ( .a(n_4131), .b(FE_OFN1117_g64577_p), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_), .o(n_4137) );
na02f04 g63381_u0 ( .a(n_3297), .b(n_2624), .o(n_4136) );
na02f06 TIMEBOOST_cell_18358 ( .a(TIMEBOOST_net_5542), .b(n_14967), .o(n_16161) );
na02f04 g63383_u0 ( .a(n_3294), .b(n_2620), .o(n_4135) );
no02f08 g63385_u0 ( .a(n_2432), .b(n_1372), .o(n_2947) );
in01m01 g63386_u0 ( .a(n_3436), .o(n_3437) );
na02m01 TIMEBOOST_cell_69308 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q), .o(TIMEBOOST_net_21862) );
na02m02 TIMEBOOST_cell_68854 ( .a(n_4452), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q), .o(TIMEBOOST_net_21635) );
ao12f02 g63390_u0 ( .a(n_2443), .b(n_3260), .c(conf_wb_err_bc_in), .o(n_4635) );
in01f02 g63392_u0 ( .a(FE_OFN1117_g64577_p), .o(g63392_sb) );
na03f01 TIMEBOOST_cell_65024 ( .a(n_4488), .b(TIMEBOOST_net_237), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q), .o(TIMEBOOST_net_17101) );
na02s02 TIMEBOOST_cell_68287 ( .a(TIMEBOOST_net_21351), .b(g65692_sb), .o(n_2206) );
na02f02 TIMEBOOST_cell_39637 ( .a(TIMEBOOST_net_11430), .b(g62787_sb), .o(n_5416) );
na02m02 TIMEBOOST_cell_69725 ( .a(TIMEBOOST_net_22070), .b(g65358_sb), .o(TIMEBOOST_net_10803) );
in01f02 g63394_u0 ( .a(n_4132), .o(n_4634) );
ao12f04 g63395_u0 ( .a(n_4131), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .c(FE_OFN1117_g64577_p), .o(n_4132) );
in01m01 g63397_u0 ( .a(FE_OFN1117_g64577_p), .o(g63397_sb) );
na02m01 TIMEBOOST_cell_43918 ( .a(TIMEBOOST_net_12853), .b(FE_OFN1074_n_4740), .o(TIMEBOOST_net_11133) );
na03f02 TIMEBOOST_cell_73407 ( .a(TIMEBOOST_net_17451), .b(FE_OFN1197_n_4090), .c(g63146_sb), .o(n_5848) );
oa12s01 g63398_u0 ( .a(n_16330), .b(n_653), .c(FE_OFN2093_n_2301), .o(n_2946) );
na02m10 TIMEBOOST_cell_25615 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52), .b(pci_target_unit_pcit_if_strd_addr_in_688), .o(TIMEBOOST_net_6912) );
in01f02 g63400_u0 ( .a(n_3160), .o(n_2943) );
na02s01 TIMEBOOST_cell_43194 ( .a(TIMEBOOST_net_12491), .b(FE_OFN250_n_9789), .o(n_9591) );
no02f08 g63402_u0 ( .a(n_2434), .b(n_1382), .o(n_2942) );
ao12f02 g63403_u0 ( .a(n_3112), .b(configuration_wb_err_addr_559), .c(n_15444), .o(n_17049) );
oa12f02 g63404_u0 ( .a(n_2701), .b(n_3304), .c(n_1998), .o(n_3432) );
ao12f02 g63406_u0 ( .a(n_3110), .b(configuration_wb_err_addr_561), .c(n_15444), .o(n_17040) );
no02f06 g63407_u0 ( .a(n_2930), .b(n_880), .o(n_3318) );
no02s02 g63409_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_13_), .b(n_1990), .o(g63409_p) );
ao12s02 g63409_u1 ( .a(g63409_p), .b(pci_target_unit_del_sync_comp_cycle_count_13_), .c(n_1990), .o(n_2721) );
ao12m02 g63410_u0 ( .a(n_3384), .b(n_4783), .c(configuration_interrupt_line_40), .o(n_4785) );
ao12f04 g63411_u0 ( .a(n_3381), .b(n_4783), .c(configuration_interrupt_line_39), .o(n_4784) );
ao12f04 g63412_u0 ( .a(n_3389), .b(n_4783), .c(configuration_interrupt_line_41), .o(n_4782) );
ao12m02 g63413_u0 ( .a(n_3387), .b(n_4783), .c(configuration_interrupt_line_43), .o(n_4781) );
oa12f02 g63414_u0 ( .a(n_2935), .b(n_2934), .c(wbm_adr_o_19_), .o(n_3317) );
oa12f02 g63415_u0 ( .a(n_2717), .b(n_2716), .c(wbu_addr_in_268), .o(n_3140) );
oa12f01 g63416_u0 ( .a(n_2715), .b(n_2714), .c(wbu_addr_in_269), .o(n_3139) );
ao12f04 g63417_u0 ( .a(n_3276), .b(n_4630), .c(wbu_cache_line_size_in_209), .o(n_4633) );
oa12f02 g63418_u0 ( .a(n_2713), .b(n_2712), .c(wbu_addr_in_272), .o(n_3138) );
oa12f02 g63419_u0 ( .a(n_3419), .b(n_1752), .c(FE_OFN1117_g64577_p), .o(n_4632) );
oa12f02 g63420_u0 ( .a(n_2707), .b(n_2706), .c(wbm_adr_o_20_), .o(n_3137) );
ao12f02 g63421_u0 ( .a(n_3274), .b(n_4630), .c(wbu_cache_line_size_in_208), .o(n_4631) );
no02f04 g63422_u0 ( .a(conf_wb_err_addr_in_964), .b(n_2398), .o(g63422_p) );
ao12f02 g63422_u1 ( .a(g63422_p), .b(conf_wb_err_addr_in_964), .c(n_2398), .o(n_3136) );
no02f04 g63423_u0 ( .a(conf_wb_err_addr_in_961), .b(n_2230), .o(g63423_p) );
ao12f02 g63423_u1 ( .a(g63423_p), .b(conf_wb_err_addr_in_961), .c(n_2230), .o(n_2941) );
no02f04 g63424_u0 ( .a(conf_wb_err_addr_in_960), .b(n_2266), .o(g63424_p) );
ao12f02 g63424_u1 ( .a(g63424_p), .b(conf_wb_err_addr_in_960), .c(n_2266), .o(n_2940) );
ao12f04 g63425_u0 ( .a(n_3279), .b(n_4630), .c(wbu_cache_line_size_in_207), .o(n_4629) );
no02m02 g63426_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_6_), .b(n_2009), .o(g63426_p) );
ao12m02 g63426_u1 ( .a(g63426_p), .b(pci_target_unit_del_sync_comp_cycle_count_6_), .c(n_2009), .o(n_2010) );
ao12f02 g63427_u0 ( .a(n_3266), .b(n_4630), .c(wbu_cache_line_size_in_211), .o(n_4628) );
no02f04 g63428_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q), .b(n_1994), .o(g63428_p) );
ao12f02 g63428_u1 ( .a(g63428_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q), .c(n_1994), .o(n_2731) );
no02m01 g63429_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_6_), .b(n_2007), .o(g63429_p) );
ao12m01 g63429_u1 ( .a(g63429_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_6_), .c(n_2007), .o(n_2008) );
no02f08 g63430_u0 ( .a(n_2227), .b(n_1399), .o(g63430_p) );
in01m01 g63431_u0 ( .a(FE_OFN1126_g64577_p), .o(g63431_sb) );
na02m10 TIMEBOOST_cell_69104 ( .a(FE_OFN1640_n_4671), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q), .o(TIMEBOOST_net_21760) );
na03f02 TIMEBOOST_cell_34897 ( .a(TIMEBOOST_net_9356), .b(FE_OFN1421_n_8567), .c(g57045_sb), .o(n_11689) );
na04f04 TIMEBOOST_cell_73324 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q), .b(FE_OFN1121_g64577_p), .c(n_3840), .d(g63037_sb), .o(n_5174) );
in01m01 g63432_u0 ( .a(FE_OFN1133_g64577_p), .o(g63432_sb) );
na02f08 TIMEBOOST_cell_53972 ( .a(TIMEBOOST_net_17203), .b(n_2769), .o(n_3008) );
na02f02 TIMEBOOST_cell_49591 ( .a(TIMEBOOST_net_86), .b(n_2132), .o(TIMEBOOST_net_15013) );
in01m01 g63433_u0 ( .a(FE_OFN1126_g64577_p), .o(g63433_sb) );
na03m02 TIMEBOOST_cell_68954 ( .a(FE_OFN654_n_4508), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q), .c(n_4473), .o(TIMEBOOST_net_21685) );
na02s01 TIMEBOOST_cell_71364 ( .a(FE_OFN203_n_9228), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q), .o(TIMEBOOST_net_22890) );
na02f02 TIMEBOOST_cell_52198 ( .a(TIMEBOOST_net_16316), .b(FE_OFN1032_n_4732), .o(TIMEBOOST_net_14919) );
in01f01 g63434_u0 ( .a(FE_OFN1126_g64577_p), .o(g63434_sb) );
na03f02 TIMEBOOST_cell_66814 ( .a(TIMEBOOST_net_16841), .b(FE_OFN1344_n_8567), .c(g57394_sb), .o(n_10374) );
na03f02 TIMEBOOST_cell_42142 ( .a(TIMEBOOST_net_8785), .b(FE_OFN1169_n_5592), .c(g62081_sb), .o(n_5628) );
in01f01 g63435_u0 ( .a(FE_OFN1125_g64577_p), .o(g63435_sb) );
na02m02 TIMEBOOST_cell_69223 ( .a(TIMEBOOST_net_21819), .b(g65278_sb), .o(TIMEBOOST_net_15242) );
na04f04 TIMEBOOST_cell_73325 ( .a(n_4053), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q), .c(FE_OFN877_g64577_p), .d(g62726_sb), .o(n_5528) );
na02s01 TIMEBOOST_cell_48509 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN525_n_9899), .o(TIMEBOOST_net_14472) );
in01m01 g63436_u0 ( .a(FE_OFN1124_g64577_p), .o(g63436_sb) );
na02s01 TIMEBOOST_cell_48511 ( .a(FE_OFN517_n_9697), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q), .o(TIMEBOOST_net_14473) );
in01m01 g63437_u0 ( .a(FE_OFN1128_g64577_p), .o(g63437_sb) );
na03m02 TIMEBOOST_cell_65058 ( .a(TIMEBOOST_net_14318), .b(g65085_sb), .c(TIMEBOOST_net_20342), .o(TIMEBOOST_net_9942) );
in01f01 g63438_u0 ( .a(FE_OFN1125_g64577_p), .o(g63438_sb) );
no04f80 TIMEBOOST_cell_20784 ( .a(FE_RN_60_0), .b(FE_RN_61_0), .c(wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_), .d(wishbone_slave_unit_fifos_outGreyCount_1_), .o(n_1829) );
na03f01 TIMEBOOST_cell_72440 ( .a(FE_OFN197_n_2683), .b(FE_OFN992_n_2373), .c(g65995_da), .o(n_2374) );
na04f04 TIMEBOOST_cell_73408 ( .a(n_4456), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q), .c(FE_OFN1246_n_4093), .d(g62713_sb), .o(n_6144) );
in01f03 g63458_u0 ( .a(n_7350), .o(n_8272) );
in01m06 g63463_u0 ( .a(n_7350), .o(n_7845) );
in01f40 g63466_u0 ( .a(n_7350), .o(n_8069) );
in01f03 g63479_u0 ( .a(n_7350), .o(n_8119) );
in01f03 g63488_u0 ( .a(n_7350), .o(n_8232) );
in01f03 g63511_u0 ( .a(n_7350), .o(n_8140) );
in01f03 g63516_u0 ( .a(n_7350), .o(n_8176) );
in01m06 g63517_u0 ( .a(n_7350), .o(n_8060) );
in01f03 g63519_u0 ( .a(n_7350), .o(n_8407) );
in01f40 g63523_u0 ( .a(n_7102), .o(n_7350) );
ao22f40 g63524_u0 ( .a(n_1036), .b(pci_target_unit_fifos_pcir_wenable_in), .c(n_659), .d(pci_target_unit_fifos_pcir_wenable_in), .o(n_7102) );
no02f04 g63525_u0 ( .a(wbm_adr_o_23_), .b(n_2414), .o(g63525_p) );
ao12f02 g63525_u1 ( .a(g63525_p), .b(wbm_adr_o_23_), .c(n_2414), .o(n_3135) );
ao12f02 g63528_u0 ( .a(n_3301), .b(n_16543), .c(configuration_wb_err_cs_bit9), .o(n_4125) );
ao12f02 g63529_u0 ( .a(n_3407), .b(FE_OFN1066_n_15808), .c(configuration_pci_err_data_503), .o(n_4619) );
in01f02 g63530_u0 ( .a(n_15262), .o(g63530_sb) );
na02s02 TIMEBOOST_cell_49287 ( .a(g58125_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q), .o(TIMEBOOST_net_14861) );
na02f02 TIMEBOOST_cell_50364 ( .a(TIMEBOOST_net_15399), .b(g62397_sb), .o(n_6806) );
na03s02 TIMEBOOST_cell_64482 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q), .b(g65923_sb), .c(g65923_db), .o(n_1565) );
ao12f02 g63531_u0 ( .a(n_3302), .b(FE_OCPN1845_n_16427), .c(n_3592), .o(n_4123) );
ao12f02 g63532_u0 ( .a(n_4088), .b(FE_OFN1695_n_3368), .c(wbu_cache_line_size_in_210), .o(n_4780) );
in01f06 g63533_u0 ( .a(FE_OFN1148_n_13249), .o(g63533_sb) );
na02s02 TIMEBOOST_cell_71133 ( .a(TIMEBOOST_net_22774), .b(TIMEBOOST_net_12471), .o(TIMEBOOST_net_15218) );
na02f08 g63533_u2 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q), .b(FE_OFN1148_n_13249), .o(g63533_db) );
na02s01 TIMEBOOST_cell_43467 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q), .o(TIMEBOOST_net_12628) );
ao12f02 g63534_u0 ( .a(n_3306), .b(n_16791), .c(pciu_bar0_in_361), .o(n_4119) );
in01m01 g63537_u0 ( .a(FE_OFN904_n_4736), .o(g63537_sb) );
na02f02 TIMEBOOST_cell_50673 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q), .b(g58292_sb), .o(TIMEBOOST_net_15554) );
na04f04 TIMEBOOST_cell_73409 ( .a(n_4369), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q), .c(FE_OFN1202_n_4090), .d(g62675_sb), .o(n_6189) );
na02s01 TIMEBOOST_cell_49476 ( .a(TIMEBOOST_net_14955), .b(g57929_db), .o(n_9881) );
in01m01 g63538_u0 ( .a(FE_OFN1074_n_4740), .o(g63538_sb) );
na03f02 TIMEBOOST_cell_64894 ( .a(TIMEBOOST_net_16587), .b(FE_OFN785_n_2678), .c(g65227_sb), .o(n_2660) );
na02f01 g63538_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q), .b(FE_OFN1074_n_4740), .o(g63538_db) );
na03f02 TIMEBOOST_cell_73410 ( .a(TIMEBOOST_net_20974), .b(FE_OFN1278_n_4097), .c(g62350_sb), .o(n_6900) );
no02f01 g63539_u0 ( .a(wbm_adr_o_12_), .b(n_2441), .o(g63539_p) );
ao12f01 g63539_u1 ( .a(g63539_p), .b(wbm_adr_o_12_), .c(n_2441), .o(n_2720) );
oa12f01 g63540_u0 ( .a(n_3420), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_), .c(FE_OFN1117_g64577_p), .o(n_4616) );
oa12f02 g63541_u0 ( .a(n_3416), .b(n_3415), .c(FE_OFN1117_g64577_p), .o(n_4614) );
no02f02 g63542_u0 ( .a(wbu_addr_in_261), .b(n_2437), .o(g63542_p) );
ao12f02 g63542_u1 ( .a(g63542_p), .b(wbu_addr_in_261), .c(n_2437), .o(n_2719) );
in01f01 g63543_u0 ( .a(FE_OFN1013_n_4734), .o(g63543_sb) );
na03f02 TIMEBOOST_cell_66750 ( .a(TIMEBOOST_net_16830), .b(FE_OFN1306_n_13124), .c(g54363_sb), .o(n_13079) );
na02f01 g63543_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q), .b(FE_OFN1013_n_4734), .o(g63543_db) );
na02m04 TIMEBOOST_cell_43919 ( .a(pci_target_unit_fifos_pciw_addr_data_in_126), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q), .o(TIMEBOOST_net_12854) );
in01f01 g63544_u0 ( .a(FE_OFN1074_n_4740), .o(g63544_sb) );
na04f04 TIMEBOOST_cell_73326 ( .a(n_3929), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q), .c(FE_OFN2105_g64577_p), .d(g63026_sb), .o(n_5194) );
na02f01 g63544_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q), .b(FE_OFN1074_n_4740), .o(g63544_db) );
in01s01 TIMEBOOST_cell_45892 ( .a(TIMEBOOST_net_13853), .o(TIMEBOOST_net_13852) );
in01m02 g63545_u0 ( .a(FE_OFN1013_n_4734), .o(g63545_sb) );
na02m01 TIMEBOOST_cell_62430 ( .a(FE_OFN2054_n_8831), .b(g58791_sb), .o(TIMEBOOST_net_20162) );
in01s01 TIMEBOOST_cell_67760 ( .a(TIMEBOOST_net_21186), .o(TIMEBOOST_net_21187) );
no02f02 g63546_u0 ( .a(n_2931), .b(wbm_adr_o_15_), .o(g63546_p) );
ao12f02 g63546_u1 ( .a(g63546_p), .b(wbm_adr_o_15_), .c(n_2931), .o(n_3134) );
in01m01 g63547_u0 ( .a(FE_OFN1046_n_16657), .o(g63547_sb) );
na02s01 g63547_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN1046_n_16657), .o(g63547_db) );
na02f01 TIMEBOOST_cell_37305 ( .a(TIMEBOOST_net_10264), .b(TIMEBOOST_net_9662), .o(n_3118) );
in01m02 g63548_u0 ( .a(FE_OFN904_n_4736), .o(g63548_sb) );
na02f04 g63548_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q), .b(FE_OFN904_n_4736), .o(g63548_db) );
na02s01 TIMEBOOST_cell_54050 ( .a(TIMEBOOST_net_17242), .b(FE_OFN1668_n_9477), .o(TIMEBOOST_net_11288) );
in01m01 g63549_u0 ( .a(FE_OFN1046_n_16657), .o(g63549_sb) );
na02f01 g63549_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q), .b(FE_OFN1046_n_16657), .o(g63549_db) );
na02f01 TIMEBOOST_cell_37309 ( .a(TIMEBOOST_net_10266), .b(TIMEBOOST_net_9663), .o(n_2718) );
in01s01 g63550_u0 ( .a(FE_OFN1125_g64577_p), .o(g63550_sb) );
no04f80 TIMEBOOST_cell_20785 ( .a(FE_RN_63_0), .b(FE_RN_64_0), .c(wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_), .d(wishbone_slave_unit_fifos_outGreyCount_0_), .o(n_1828) );
na03f02 TIMEBOOST_cell_47307 ( .a(FE_OFN1551_n_12104), .b(TIMEBOOST_net_13592), .c(FE_OCPN1827_n_14995), .o(n_12654) );
in01f01 g63551_u0 ( .a(FE_OFN1128_g64577_p), .o(g63551_sb) );
na02m01 TIMEBOOST_cell_45455 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q), .o(TIMEBOOST_net_13622) );
na02s01 TIMEBOOST_cell_25303 ( .a(pci_ad_i_30_), .b(n_2509), .o(TIMEBOOST_net_6756) );
in01m01 g63552_u0 ( .a(FE_OFN1133_g64577_p), .o(g63552_sb) );
na02s01 TIMEBOOST_cell_48818 ( .a(TIMEBOOST_net_14626), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_9495) );
na03m02 TIMEBOOST_cell_42007 ( .a(g58400_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q), .c(g58400_db), .o(n_9208) );
na02f06 TIMEBOOST_cell_63812 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_401), .b(FE_OFN2057_n_2117), .o(TIMEBOOST_net_20892) );
in01f01 g63553_u0 ( .a(FE_OFN1128_g64577_p), .o(g63553_sb) );
na03f02 TIMEBOOST_cell_73256 ( .a(TIMEBOOST_net_23310), .b(TIMEBOOST_net_16365), .c(FE_OFN1135_g64577_p), .o(TIMEBOOST_net_22491) );
na02m04 TIMEBOOST_cell_69232 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q), .b(FE_OFN642_n_4677), .o(TIMEBOOST_net_21824) );
na02f02 TIMEBOOST_cell_72243 ( .a(TIMEBOOST_net_23329), .b(g59371_sb), .o(n_7692) );
in01m01 g63554_u0 ( .a(FE_OFN1133_g64577_p), .o(g63554_sb) );
na02f04 TIMEBOOST_cell_45456 ( .a(FE_OFN1558_n_12042), .b(TIMEBOOST_net_13622), .o(TIMEBOOST_net_12027) );
na03f02 TIMEBOOST_cell_42036 ( .a(TIMEBOOST_net_5273), .b(g62106_sb), .c(g62106_db), .o(n_5594) );
na03s02 TIMEBOOST_cell_72877 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q), .b(g63568_sb), .c(g63568_db), .o(n_4594) );
in01m01 g63555_u0 ( .a(FE_OFN1126_g64577_p), .o(g63555_sb) );
na03m02 TIMEBOOST_cell_64958 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q), .b(g64241_sb), .c(g64241_db), .o(n_3931) );
in01f01 g63556_u0 ( .a(FE_OFN1125_g64577_p), .o(g63556_sb) );
na02m01 g65888_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q), .b(FE_OFN682_n_4460), .o(g65888_db) );
na03f02 TIMEBOOST_cell_42042 ( .a(TIMEBOOST_net_5271), .b(g62134_sb), .c(g62134_db), .o(n_5559) );
na02f02 TIMEBOOST_cell_49592 ( .a(TIMEBOOST_net_15013), .b(TIMEBOOST_net_118), .o(n_4680) );
in01m01 g63557_u0 ( .a(FE_OFN1126_g64577_p), .o(g63557_sb) );
na03m02 TIMEBOOST_cell_70160 ( .a(FE_OFN1077_n_4740), .b(pci_target_unit_fifos_pciw_addr_data_in_147), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q), .o(TIMEBOOST_net_22288) );
na03m02 TIMEBOOST_cell_72803 ( .a(TIMEBOOST_net_21559), .b(g64891_sb), .c(TIMEBOOST_net_21829), .o(TIMEBOOST_net_17413) );
ao12f02 g63558_u0 ( .a(n_3125), .b(n_15808), .c(configuration_pci_err_data), .o(n_3428) );
in01f04 g63559_u0 ( .a(FE_OFN1117_g64577_p), .o(g63559_sb) );
na03s02 TIMEBOOST_cell_41908 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q), .b(g58276_sb), .c(g58276_db), .o(n_9034) );
na02s01 g58377_u2 ( .a(FE_OFN260_n_9860), .b(FE_OFN579_n_9531), .o(g58377_db) );
in01f02 g63560_u0 ( .a(FE_OFN1092_g64577_p), .o(g63560_sb) );
na02s01 TIMEBOOST_cell_68499 ( .a(TIMEBOOST_net_21457), .b(g66403_db), .o(n_2537) );
in01s01 TIMEBOOST_cell_67776 ( .a(TIMEBOOST_net_21202), .o(TIMEBOOST_net_21203) );
in01f02 g63561_u0 ( .a(FE_OFN1092_g64577_p), .o(g63561_sb) );
na02m08 TIMEBOOST_cell_17982 ( .a(TIMEBOOST_net_5354), .b(n_785), .o(TIMEBOOST_net_171) );
na02m08 TIMEBOOST_cell_17981 ( .a(n_245), .b(n_193), .o(TIMEBOOST_net_5354) );
in01f01 g63562_u0 ( .a(FE_OFN1092_g64577_p), .o(g63562_sb) );
na04f03 TIMEBOOST_cell_67880 ( .a(FE_OFN642_n_4677), .b(n_4493), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q), .d(g65292_sb), .o(n_4283) );
na02f01 TIMEBOOST_cell_17979 ( .a(n_2742), .b(n_3503), .o(TIMEBOOST_net_5353) );
in01m02 g63563_u0 ( .a(FE_OFN1058_n_4727), .o(g63563_sb) );
na04m08 TIMEBOOST_cell_72566 ( .a(FE_OFN659_n_4392), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q), .c(n_3780), .d(g64938_sb), .o(n_3676) );
in01s01 g63564_u0 ( .a(FE_OFN1057_n_4727), .o(g63564_sb) );
na02f02 TIMEBOOST_cell_37603 ( .a(TIMEBOOST_net_10413), .b(g58094_db), .o(n_9082) );
in01m01 g63565_u0 ( .a(FE_OFN918_n_4725), .o(g63565_sb) );
na02s01 TIMEBOOST_cell_43625 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q), .b(FE_OFN539_n_9690), .o(TIMEBOOST_net_12707) );
na02m02 g63565_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(FE_OFN918_n_4725), .o(g63565_db) );
na03m02 TIMEBOOST_cell_73411 ( .a(TIMEBOOST_net_21002), .b(FE_OFN1279_n_4097), .c(g62390_sb), .o(n_6819) );
in01m01 g63566_u0 ( .a(FE_OFN1031_n_4732), .o(g63566_sb) );
na03s02 TIMEBOOST_cell_73676 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q), .b(g57975_sb), .c(FE_OFN252_n_9868), .o(TIMEBOOST_net_16754) );
na04f02 TIMEBOOST_cell_73257 ( .a(n_2153), .b(FE_OFN2212_n_8407), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q), .d(g62019_sb), .o(n_7857) );
in01m01 g63567_u0 ( .a(FE_OFN929_n_4730), .o(g63567_sb) );
na03f02 TIMEBOOST_cell_66286 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q), .b(g62580_sb), .c(g62580_db), .o(n_6393) );
na02m01 g63567_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(FE_OFN929_n_4730), .o(g63567_db) );
na02f02 TIMEBOOST_cell_43933 ( .a(conf_wb_err_addr_in_958), .b(n_3347), .o(TIMEBOOST_net_12861) );
in01s01 g63568_u0 ( .a(FE_OFN929_n_4730), .o(g63568_sb) );
na02m01 TIMEBOOST_cell_69290 ( .a(n_4442), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q), .o(TIMEBOOST_net_21853) );
na02s01 g63568_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_121), .b(FE_OFN929_n_4730), .o(g63568_db) );
na02m04 TIMEBOOST_cell_68724 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q), .b(FE_OFN687_n_4417), .o(TIMEBOOST_net_21570) );
in01m01 g63569_u0 ( .a(FE_OFN1031_n_4732), .o(g63569_sb) );
na02f02 TIMEBOOST_cell_70331 ( .a(TIMEBOOST_net_22373), .b(FE_OFN1812_n_7845), .o(TIMEBOOST_net_15100) );
na02s06 TIMEBOOST_cell_47553 ( .a(wbs_dat_i_6_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q), .o(TIMEBOOST_net_13994) );
in01m01 g63570_u0 ( .a(FE_OFN918_n_4725), .o(g63570_sb) );
na03s02 TIMEBOOST_cell_65259 ( .a(TIMEBOOST_net_14544), .b(g65766_sb), .c(TIMEBOOST_net_14588), .o(n_8173) );
na02m01 g63570_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(FE_OFN918_n_4725), .o(g63570_db) );
na03s01 TIMEBOOST_cell_72501 ( .a(FE_OFN527_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q), .c(FE_OFN211_n_9858), .o(TIMEBOOST_net_12762) );
in01f04 g63571_u0 ( .a(FE_OFN1117_g64577_p), .o(g63571_sb) );
na03m02 TIMEBOOST_cell_72502 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q), .b(g65425_sb), .c(g65425_db), .o(n_3510) );
na02f02 TIMEBOOST_cell_70215 ( .a(TIMEBOOST_net_22315), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_15052) );
in01f01 g63572_u0 ( .a(FE_OFN1092_g64577_p), .o(g63572_sb) );
na02s02 TIMEBOOST_cell_68397 ( .a(TIMEBOOST_net_21406), .b(TIMEBOOST_net_16145), .o(TIMEBOOST_net_14167) );
na03s02 TIMEBOOST_cell_72657 ( .a(TIMEBOOST_net_21123), .b(FE_OFN1015_n_2053), .c(TIMEBOOST_net_14488), .o(TIMEBOOST_net_22358) );
na04f04 TIMEBOOST_cell_73258 ( .a(n_1862), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q), .c(FE_OFN2212_n_8407), .d(g61907_sb), .o(n_8007) );
in01f02 g63573_u0 ( .a(FE_OFN1092_g64577_p), .o(g63573_sb) );
na02f20 TIMEBOOST_cell_17976 ( .a(TIMEBOOST_net_5351), .b(n_2028), .o(TIMEBOOST_net_166) );
na02s02 TIMEBOOST_cell_38436 ( .a(FE_OFN252_n_9868), .b(g57944_sb), .o(TIMEBOOST_net_10830) );
in01f02 g63574_u0 ( .a(FE_OFN1092_g64577_p), .o(g63574_sb) );
na02m02 TIMEBOOST_cell_48801 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q), .b(g58279_sb), .o(TIMEBOOST_net_14618) );
ao22s01 g63575_u0 ( .a(n_1180), .b(n_1999), .c(n_3250), .d(pci_target_unit_wishbone_master_read_count_reg_2__Q), .o(n_3316) );
in01f02 g63576_u0 ( .a(FE_OFN1698_n_5751), .o(g63576_sb) );
na02f02 TIMEBOOST_cell_69375 ( .a(TIMEBOOST_net_21895), .b(g60671_sb), .o(TIMEBOOST_net_5478) );
na04m02 TIMEBOOST_cell_67206 ( .a(TIMEBOOST_net_10314), .b(g65286_sb), .c(n_4479), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q), .o(TIMEBOOST_net_17422) );
in01f02 g63577_u0 ( .a(FE_OFN1700_n_5751), .o(g63577_sb) );
in01m04 TIMEBOOST_cell_35481 ( .a(TIMEBOOST_net_10071), .o(TIMEBOOST_net_10072) );
na02m04 TIMEBOOST_cell_69088 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q), .b(n_3785), .o(TIMEBOOST_net_21752) );
no02f08 g63578_u0 ( .a(wbu_addr_in_264), .b(n_3132), .o(g63578_p) );
ao12f04 g63578_u1 ( .a(g63578_p), .b(wbu_addr_in_264), .c(n_3132), .o(n_3133) );
no02f04 g63579_u0 ( .a(conf_wb_err_addr_in_953), .b(n_2722), .o(g63579_p) );
ao12f02 g63579_u1 ( .a(g63579_p), .b(conf_wb_err_addr_in_953), .c(n_2722), .o(n_2744) );
no02f04 g63580_u0 ( .a(conf_wb_err_addr_in_956), .b(n_3130), .o(g63580_p) );
ao12f02 g63580_u1 ( .a(g63580_p), .b(conf_wb_err_addr_in_956), .c(n_3130), .o(n_3131) );
no02f04 g63581_u0 ( .a(FE_OFN1698_n_5751), .b(wbm_adr_o_2_), .o(g63581_p) );
ao12f02 g63581_u1 ( .a(g63581_p), .b(wbm_adr_o_2_), .c(FE_OFN1698_n_5751), .o(n_3425) );
in01s01 g63582_u0 ( .a(FE_OFN1021_n_11877), .o(g63582_sb) );
na02f01 g63582_u2 ( .a(wbu_addr_in), .b(FE_OFN1021_n_11877), .o(g63582_db) );
na03f02 TIMEBOOST_cell_66534 ( .a(g53921_sb), .b(FE_OFN1331_n_13547), .c(TIMEBOOST_net_16796), .o(n_13523) );
na02s02 TIMEBOOST_cell_37997 ( .a(TIMEBOOST_net_10610), .b(g58120_sb), .o(n_9076) );
in01s01 g63584_u0 ( .a(FE_OFN1025_n_11877), .o(g63584_sb) );
na03s02 TIMEBOOST_cell_72584 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q), .b(TIMEBOOST_net_20577), .c(FE_OFN233_n_9876), .o(TIMEBOOST_net_16763) );
na02s01 g63584_u2 ( .a(wbu_sel_in), .b(FE_OFN1025_n_11877), .o(g63584_db) );
na02s01 TIMEBOOST_cell_38417 ( .a(TIMEBOOST_net_10820), .b(g57951_db), .o(n_9125) );
na03f02 TIMEBOOST_cell_47285 ( .a(FE_OFN1736_n_16317), .b(TIMEBOOST_net_13582), .c(FE_OFN1741_n_11019), .o(n_12617) );
na02s01 g63585_u2 ( .a(wbu_sel_in_312), .b(FE_OFN1025_n_11877), .o(g63585_db) );
na02f04 TIMEBOOST_cell_54253 ( .a(TIMEBOOST_net_13130), .b(n_2120), .o(TIMEBOOST_net_17344) );
in01s01 g63586_u0 ( .a(FE_OFN1025_n_11877), .o(g63586_sb) );
na03s02 TIMEBOOST_cell_72399 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_92), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .c(g54209_sb), .o(TIMEBOOST_net_20795) );
na02s01 g63586_u2 ( .a(wbu_sel_in_313), .b(FE_OFN1025_n_11877), .o(g63586_db) );
na02m01 TIMEBOOST_cell_38003 ( .a(TIMEBOOST_net_10613), .b(g58082_db), .o(n_9085) );
na04f04 TIMEBOOST_cell_73062 ( .a(n_1593), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q), .c(FE_OFN714_n_8140), .d(g61805_sb), .o(n_8184) );
na02s01 g63587_u2 ( .a(wbu_sel_in_314), .b(FE_OFN1025_n_11877), .o(g63587_db) );
no03f02 TIMEBOOST_cell_73729 ( .a(TIMEBOOST_net_13633), .b(FE_RN_723_0), .c(FE_OCP_RBN2291_FE_OFN1575_n_12028), .o(n_12725) );
in01m01 g63588_u0 ( .a(FE_OFN9_n_11877), .o(g63588_sb) );
na02m02 TIMEBOOST_cell_38076 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q), .b(g65343_sb), .o(TIMEBOOST_net_10650) );
na02f01 g63588_u2 ( .a(n_16945), .b(FE_OFN9_n_11877), .o(g63588_db) );
in01m01 g63589_u0 ( .a(FE_OFN2_n_4778), .o(g63589_sb) );
na03m06 TIMEBOOST_cell_69596 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q), .b(g65412_sb), .c(FE_OFN639_n_4669), .o(TIMEBOOST_net_22006) );
na02s02 TIMEBOOST_cell_38438 ( .a(FE_OFN215_n_9856), .b(g57920_sb), .o(TIMEBOOST_net_10831) );
in01f04 g63590_u0 ( .a(FE_OFN989_n_574), .o(g63590_sb) );
na03m02 TIMEBOOST_cell_73008 ( .a(TIMEBOOST_net_21863), .b(FE_OFN1810_n_4454), .c(TIMEBOOST_net_22120), .o(TIMEBOOST_net_17393) );
na02s01 g63590_u2 ( .a(pci_inti_conf_int_in), .b(FE_OFN989_n_574), .o(g63590_db) );
in01m01 g63591_u0 ( .a(FE_OFN2021_n_4778), .o(g63591_sb) );
na02s02 TIMEBOOST_cell_48784 ( .a(TIMEBOOST_net_14609), .b(TIMEBOOST_net_11084), .o(TIMEBOOST_net_9468) );
na03s02 TIMEBOOST_cell_33801 ( .a(n_2191), .b(g61703_sb), .c(g61703_db), .o(n_8421) );
na03f02 TIMEBOOST_cell_47281 ( .a(FE_OFN1735_n_16317), .b(TIMEBOOST_net_13579), .c(FE_OFN1739_n_11019), .o(n_12743) );
in01m01 g63592_u0 ( .a(FE_OFN2_n_4778), .o(g63592_sb) );
na02f02 TIMEBOOST_cell_39549 ( .a(TIMEBOOST_net_11386), .b(g62764_sb), .o(n_5467) );
na02s01 TIMEBOOST_cell_63216 ( .a(TIMEBOOST_net_12567), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q), .o(TIMEBOOST_net_20555) );
na02s02 TIMEBOOST_cell_38442 ( .a(FE_OFN215_n_9856), .b(g57983_sb), .o(TIMEBOOST_net_10833) );
in01m01 g63593_u0 ( .a(FE_OFN2_n_4778), .o(g63593_sb) );
na03f02 TIMEBOOST_cell_65924 ( .a(TIMEBOOST_net_20895), .b(n_13825), .c(g61843_sb), .o(n_7212) );
in01s01 TIMEBOOST_cell_63534 ( .a(TIMEBOOST_net_20714), .o(wbs_adr_i_12_) );
in01m01 g63594_u0 ( .a(FE_OFN2021_n_4778), .o(g63594_sb) );
na02s01 TIMEBOOST_cell_42729 ( .a(g58793_sb), .b(n_8831), .o(TIMEBOOST_net_12259) );
na02f02 TIMEBOOST_cell_71080 ( .a(TIMEBOOST_net_20636), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_22748) );
na04f04 TIMEBOOST_cell_67925 ( .a(TIMEBOOST_net_7283), .b(FE_OFN1149_n_13249), .c(TIMEBOOST_net_20892), .d(g54135_sb), .o(n_13670) );
in01m01 g63595_u0 ( .a(FE_OFN2_n_4778), .o(g63595_sb) );
na02s01 TIMEBOOST_cell_38444 ( .a(FE_OFN213_n_9124), .b(g57982_sb), .o(TIMEBOOST_net_10834) );
na03f02 TIMEBOOST_cell_73702 ( .a(TIMEBOOST_net_13685), .b(FE_OFN1760_n_10780), .c(FE_OFN1579_n_12306), .o(n_12734) );
in01m01 g63596_u0 ( .a(FE_OFN2_n_4778), .o(g63596_sb) );
na04m02 TIMEBOOST_cell_72926 ( .a(TIMEBOOST_net_12639), .b(FE_OFN1678_n_4655), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q), .d(g65897_sb), .o(TIMEBOOST_net_17030) );
na03f02 TIMEBOOST_cell_66834 ( .a(TIMEBOOST_net_16456), .b(g59382_db), .c(g52401_db), .o(n_14818) );
in01s01 g63597_u0 ( .a(FE_OFN1079_n_4778), .o(g63597_sb) );
na02s02 TIMEBOOST_cell_38600 ( .a(g58006_sb), .b(FE_OFN254_n_9825), .o(TIMEBOOST_net_10912) );
na02s01 TIMEBOOST_cell_52611 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q), .o(TIMEBOOST_net_16523) );
in01f01 g63598_u0 ( .a(FE_OFN2022_n_4778), .o(g63598_sb) );
na02m20 TIMEBOOST_cell_42717 ( .a(wishbone_slave_unit_pci_initiator_if_data_source), .b(g54160_sb), .o(TIMEBOOST_net_12253) );
na03s02 TIMEBOOST_cell_66379 ( .a(TIMEBOOST_net_14644), .b(g58180_sb), .c(TIMEBOOST_net_14849), .o(TIMEBOOST_net_9547) );
in01s01 g63599_u0 ( .a(FE_OFN1079_n_4778), .o(g63599_sb) );
na02f02 TIMEBOOST_cell_39381 ( .a(TIMEBOOST_net_11302), .b(g63559_sb), .o(n_4115) );
na02s01 g63599_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q), .b(FE_OFN1079_n_4778), .o(g63599_db) );
na02f02 TIMEBOOST_cell_49860 ( .a(TIMEBOOST_net_15147), .b(g63176_sb), .o(n_4947) );
in01m01 g63600_u0 ( .a(FE_OFN2021_n_4778), .o(g63600_sb) );
na03f02 TIMEBOOST_cell_35073 ( .a(TIMEBOOST_net_9591), .b(FE_OFN1440_n_9372), .c(g58486_sb), .o(n_9348) );
na02s01 TIMEBOOST_cell_38595 ( .a(TIMEBOOST_net_10909), .b(g58045_db), .o(n_9745) );
in01m01 g63601_u0 ( .a(FE_OFN2022_n_4778), .o(g63601_sb) );
na02s01 TIMEBOOST_cell_52613 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q), .o(TIMEBOOST_net_16524) );
na02s01 g63601_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q), .b(FE_OFN1079_n_4778), .o(g63601_db) );
na02s01 TIMEBOOST_cell_38450 ( .a(g58099_sb), .b(FE_OFN252_n_9868), .o(TIMEBOOST_net_10837) );
in01s01 g63602_u0 ( .a(FE_OFN1079_n_4778), .o(g63602_sb) );
na02s01 g63602_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q), .b(FE_OFN1079_n_4778), .o(g63602_db) );
in01s01 TIMEBOOST_cell_67715 ( .a(pci_target_unit_fifos_pcir_data_in_184), .o(TIMEBOOST_net_21142) );
in01s01 g63603_u0 ( .a(FE_OFN1079_n_4778), .o(g63603_sb) );
in01s01 TIMEBOOST_cell_67717 ( .a(pci_target_unit_fifos_pcir_data_in_187), .o(TIMEBOOST_net_21144) );
na02s01 g63603_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q), .b(FE_OFN1079_n_4778), .o(g63603_db) );
na04f04 TIMEBOOST_cell_36105 ( .a(parchk_pci_ad_out_in_1184), .b(g62087_sb), .c(configuration_wb_err_data_587), .d(FE_OFN1173_n_5592), .o(n_5620) );
in01m01 g63604_u0 ( .a(FE_OFN2021_n_4778), .o(g63604_sb) );
in01s01 TIMEBOOST_cell_63611 ( .a(TIMEBOOST_net_20791), .o(TIMEBOOST_net_20790) );
in01s01 g63605_u0 ( .a(FE_OFN1079_n_4778), .o(g63605_sb) );
na02s01 TIMEBOOST_cell_49510 ( .a(TIMEBOOST_net_14972), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9480) );
na02s01 g63605_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q), .b(FE_OFN1079_n_4778), .o(g63605_db) );
na02s02 TIMEBOOST_cell_54544 ( .a(TIMEBOOST_net_17489), .b(TIMEBOOST_net_12818), .o(TIMEBOOST_net_9422) );
in01m01 g63606_u0 ( .a(FE_OFN2_n_4778), .o(g63606_sb) );
na03m02 TIMEBOOST_cell_73009 ( .a(g65375_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q), .c(TIMEBOOST_net_7098), .o(TIMEBOOST_net_20532) );
in01s01 g63607_u0 ( .a(FE_OFN1079_n_4778), .o(g63607_sb) );
na02s01 g63607_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q), .b(FE_OFN1079_n_4778), .o(g63607_db) );
in01f01 g63608_u0 ( .a(FE_OFN2022_n_4778), .o(g63608_sb) );
na02s04 TIMEBOOST_cell_45599 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q), .o(TIMEBOOST_net_13694) );
na03m02 TIMEBOOST_cell_65141 ( .a(TIMEBOOST_net_16925), .b(g64876_sb), .c(TIMEBOOST_net_17260), .o(TIMEBOOST_net_13230) );
na02s01 TIMEBOOST_cell_62756 ( .a(g61708_sb), .b(g61708_db), .o(TIMEBOOST_net_20325) );
in01m01 g63609_u0 ( .a(FE_OFN2_n_4778), .o(g63609_sb) );
na02m01 TIMEBOOST_cell_62542 ( .a(pci_target_unit_fifos_pciw_addr_data_in_124), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_20218) );
in01m01 g63610_u0 ( .a(FE_OFN2021_n_4778), .o(g63610_sb) );
na03f02 TIMEBOOST_cell_35069 ( .a(TIMEBOOST_net_9614), .b(FE_OFN1439_n_9372), .c(g58482_sb), .o(n_8975) );
na02m01 TIMEBOOST_cell_43225 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_12507) );
na03f02 TIMEBOOST_cell_34765 ( .a(TIMEBOOST_net_9349), .b(FE_OFN1411_n_8567), .c(g57383_sb), .o(n_11362) );
in01s01 g63611_u0 ( .a(FE_OFN1079_n_4778), .o(g63611_sb) );
na02m02 TIMEBOOST_cell_68799 ( .a(TIMEBOOST_net_21607), .b(TIMEBOOST_net_10536), .o(TIMEBOOST_net_17521) );
na02s01 g63611_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q), .b(FE_OFN1079_n_4778), .o(g63611_db) );
na02s01 TIMEBOOST_cell_47965 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q), .o(TIMEBOOST_net_14200) );
in01s01 g63612_u0 ( .a(FE_OFN1079_n_4778), .o(g63612_sb) );
na02f02 TIMEBOOST_cell_70991 ( .a(TIMEBOOST_net_22703), .b(g62991_sb), .o(n_5900) );
na03f02 TIMEBOOST_cell_34870 ( .a(TIMEBOOST_net_9371), .b(FE_OFN1382_n_8567), .c(g57191_sb), .o(n_10447) );
in01s01 TIMEBOOST_cell_73896 ( .a(n_8166), .o(TIMEBOOST_net_23461) );
in01s01 g63613_u0 ( .a(FE_OFN1079_n_4778), .o(g63613_sb) );
na04f04 TIMEBOOST_cell_36852 ( .a(n_8560), .b(g58588_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q), .d(FE_OFN1403_n_8567), .o(n_8914) );
na02s01 g63613_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q), .b(FE_OFN1079_n_4778), .o(g63613_db) );
na02m01 TIMEBOOST_cell_69797 ( .a(TIMEBOOST_net_22106), .b(n_4450), .o(TIMEBOOST_net_17381) );
in01s01 g63614_u0 ( .a(FE_OFN1079_n_4778), .o(g63614_sb) );
na02s01 g63614_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q), .b(FE_OFN1079_n_4778), .o(g63614_db) );
na02f02 TIMEBOOST_cell_28008 ( .a(n_13901), .b(TIMEBOOST_net_8108), .o(TIMEBOOST_net_758) );
in01f01 g63615_u0 ( .a(FE_OFN2022_n_4778), .o(g63615_sb) );
na02s02 TIMEBOOST_cell_71908 ( .a(TIMEBOOST_net_20215), .b(FE_OFN953_n_2055), .o(TIMEBOOST_net_23162) );
na02m02 TIMEBOOST_cell_62540 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_130), .o(TIMEBOOST_net_20217) );
in01m01 g63616_u0 ( .a(FE_OFN2_n_4778), .o(g63616_sb) );
na03f02 TIMEBOOST_cell_73127 ( .a(TIMEBOOST_net_22135), .b(g64234_sb), .c(FE_OFN2104_g64577_p), .o(TIMEBOOST_net_22485) );
in01m01 g63617_u0 ( .a(FE_OFN2021_n_4778), .o(g63617_sb) );
na02f02 TIMEBOOST_cell_18030 ( .a(TIMEBOOST_net_5378), .b(n_4743), .o(TIMEBOOST_net_321) );
na02f01 TIMEBOOST_cell_18029 ( .a(n_3503), .b(n_2308), .o(TIMEBOOST_net_5378) );
in01m01 g63618_u0 ( .a(FE_OFN2022_n_4778), .o(g63618_sb) );
na03f02 TIMEBOOST_cell_73259 ( .a(TIMEBOOST_net_23311), .b(TIMEBOOST_net_16359), .c(FE_OFN1119_g64577_p), .o(TIMEBOOST_net_22492) );
na02s01 g63618_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q), .b(FE_OFN1079_n_4778), .o(g63618_db) );
na02f02 TIMEBOOST_cell_71742 ( .a(TIMEBOOST_net_13803), .b(n_13903), .o(TIMEBOOST_net_23079) );
in01s01 g63619_u0 ( .a(FE_OFN1079_n_4778), .o(g63619_sb) );
na02s01 TIMEBOOST_cell_42722 ( .a(TIMEBOOST_net_12255), .b(n_2373), .o(TIMEBOOST_net_10154) );
na02s01 g63619_u2 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q), .b(FE_OFN1079_n_4778), .o(g63619_db) );
na02s01 TIMEBOOST_cell_42724 ( .a(TIMEBOOST_net_12256), .b(n_2373), .o(TIMEBOOST_net_10157) );
in01f01 g63620_u0 ( .a(FE_OFN2022_n_4778), .o(g63620_sb) );
na03f02 TIMEBOOST_cell_35071 ( .a(TIMEBOOST_net_9586), .b(FE_OFN1436_n_9372), .c(g58461_sb), .o(n_9393) );
na03m02 TIMEBOOST_cell_72683 ( .a(g64788_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q), .c(TIMEBOOST_net_14278), .o(TIMEBOOST_net_13227) );
in01m01 g63621_u0 ( .a(FE_OFN2021_n_4778), .o(g63621_sb) );
na02f02 TIMEBOOST_cell_54388 ( .a(TIMEBOOST_net_17411), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_15455) );
in01f20 g63667_u0 ( .a(pciu_cache_lsize_not_zero_in), .o(n_3319) );
na02f02 g63682_u0 ( .a(n_1472), .b(n_3809), .o(n_4746) );
in01f06 g63695_u0 ( .a(FE_OFN1155_n_3464), .o(n_4098) );
in01f08 g63708_u0 ( .a(FE_OFN1154_n_3464), .o(n_4097) );
in01f04 g63721_u0 ( .a(FE_OFN1155_n_3464), .o(n_4096) );
in01f06 g63734_u0 ( .a(FE_OFN1154_n_3464), .o(n_4095) );
in01f06 g63747_u0 ( .a(FE_OFN1155_n_3464), .o(n_4143) );
in01f08 g63773_u0 ( .a(FE_OFN1154_n_3464), .o(n_4093) );
in01f06 g63786_u0 ( .a(FE_OFN1155_n_3464), .o(n_4092) );
in01f20 g63799_u0 ( .a(FE_OFN1155_n_3464), .o(n_6391) );
in01f04 g63803_u0 ( .a(FE_OFN1154_n_3464), .o(n_6886) );
in01f06 g63834_u0 ( .a(FE_OFN1154_n_3464), .o(n_4151) );
in01f04 g63838_u0 ( .a(FE_OFN1154_n_3464), .o(n_6356) );
in01f04 g63847_u0 ( .a(FE_OFN1155_n_3464), .o(n_4090) );
in01f10 g63853_u0 ( .a(n_4658), .o(n_6431) );
in01f20 g63860_u0 ( .a(n_4658), .o(n_6436) );
in01f10 g63861_u0 ( .a(n_4658), .o(n_6554) );
in01f10 g63862_u0 ( .a(n_4658), .o(n_6319) );
in01f10 g63864_u0 ( .a(n_4658), .o(n_6287) );
in01f10 g63868_u0 ( .a(n_4658), .o(n_6645) );
in01f20 g63870_u0 ( .a(n_4658), .o(n_6232) );
in01f80 g63881_u0 ( .a(n_4658), .o(n_6624) );
in01f80 g63888_u0 ( .a(FE_OFN1192_n_6935), .o(n_4658) );
in01f20 g63889_u0 ( .a(FE_OFN1155_n_3464), .o(n_6935) );
na02f10 g63890_u0 ( .a(n_3314), .b(n_3313), .o(n_3464) );
no02f08 g63891_u0 ( .a(n_868), .b(FE_OFN1117_g64577_p), .o(g63891_p) );
in01f04 g63891_u1 ( .a(g63891_p), .o(n_4637) );
na02f02 g63892_u0 ( .a(n_646), .b(n_1825), .o(g63892_p) );
in01s01 g63892_u1 ( .a(g63892_p), .o(n_2445) );
no02m01 g63894_u0 ( .a(n_963), .b(FE_OFN778_n_4152), .o(n_2938) );
na02f02 g63895_u0 ( .a(n_3053), .b(n_4806), .o(g63895_p) );
in01f02 g63895_u1 ( .a(g63895_p), .o(n_3424) );
in01m02 g63896_u0 ( .a(n_2950), .o(n_14389) );
no02f10 g63897_u0 ( .a(n_1964), .b(n_2443), .o(n_2950) );
na02f01 g63899_u0 ( .a(FE_OFN1024_n_11877), .b(n_16818), .o(n_3423) );
in01f06 g63900_u0 ( .a(n_3421), .o(n_3422) );
na02f08 g63902_u0 ( .a(n_2441), .b(n_2433), .o(g63902_p) );
in01f04 g63902_u1 ( .a(g63902_p), .o(n_2442) );
na02f01 g63905_u0 ( .a(n_2727), .b(FE_OFN1619_n_1787), .o(n_2728) );
na02f04 g63907_u0 ( .a(n_2813), .b(n_2814), .o(n_3306) );
no02f01 g63908_u0 ( .a(n_1701), .b(FE_OFN778_n_4152), .o(n_2937) );
na02f01 g63909_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_), .b(FE_OFN1117_g64577_p), .o(n_3420) );
na02f04 g63910_u0 ( .a(n_3235), .b(n_2847), .o(n_4088) );
na02f04 g63911_u0 ( .a(n_2716), .b(wbu_addr_in_268), .o(n_2717) );
na02f01 g63912_u0 ( .a(n_2714), .b(wbu_addr_in_269), .o(n_2715) );
no02s01 g63914_u0 ( .a(n_4533), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_0_), .o(n_4537) );
na02f04 g63915_u0 ( .a(n_2712), .b(wbu_addr_in_272), .o(n_2713) );
na02f08 g63916_u0 ( .a(n_2727), .b(wishbone_slave_unit_pci_initiator_if_current_byte_address), .o(g63916_p) );
in01f04 g63916_u1 ( .a(g63916_p), .o(n_2711) );
na02f06 g63919_u0 ( .a(FE_OFN1117_g64577_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_), .o(n_3419) );
na02f02 g63920_u0 ( .a(FE_OFN1092_g64577_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_), .o(n_3417) );
na02f04 g63921_u0 ( .a(n_3415), .b(FE_OFN1117_g64577_p), .o(n_3416) );
na02f01 g63922_u0 ( .a(n_2437), .b(n_2431), .o(g63922_p) );
in01f02 g63922_u1 ( .a(g63922_p), .o(n_2438) );
na02f01 TIMEBOOST_cell_37308 ( .a(n_1192), .b(FE_OFN989_n_574), .o(TIMEBOOST_net_10266) );
in01f01 g63924_u0 ( .a(n_4535), .o(n_4536) );
no02f10 g63925_u0 ( .a(wishbone_slave_unit_pcim_sm_rdy_in), .b(FE_OFN999_n_15978), .o(g63925_p) );
in01f08 g63925_u1 ( .a(g63925_p), .o(n_4535) );
no02f04 g63926_u0 ( .a(FE_OFN967_n_2233), .b(n_3080), .o(n_3413) );
no02f06 g63927_u0 ( .a(FE_OFN1117_g64577_p), .b(pci_target_unit_fifos_pciw_control_in), .o(n_5546) );
no02f04 g63929_u0 ( .a(n_2231), .b(n_2232), .o(n_2710) );
na02f08 g63930_u0 ( .a(n_2722), .b(n_2435), .o(n_2436) );
na02f04 g63933_u0 ( .a(n_2934), .b(wbm_adr_o_19_), .o(n_2935) );
no02f01 g63934_u0 ( .a(n_1204), .b(n_4533), .o(n_4534) );
no02f04 g63935_u0 ( .a(n_2402), .b(n_2401), .o(g63935_p) );
in01f02 g63935_u1 ( .a(g63935_p), .o(n_2933) );
no02f02 g63936_u0 ( .a(n_2400), .b(n_2876), .o(n_3305) );
no02f06 g63938_u0 ( .a(n_2214), .b(FE_OCP_RBN2239_g74749_p), .o(n_4642) );
na02f04 g63939_u0 ( .a(pci_target_unit_wishbone_master_burst_chopped), .b(FE_OCP_RBN2237_g74749_p), .o(g63939_p) );
in01f02 g63939_u1 ( .a(g63939_p), .o(n_3410) );
na02f06 g63940_u0 ( .a(n_3304), .b(n_16159), .o(n_4674) );
no02f08 g63941_u0 ( .a(n_1998), .b(FE_OCP_RBN2239_g74749_p), .o(n_3409) );
no02s01 g63942_u0 ( .a(FE_OFN778_n_4152), .b(pci_target_unit_del_sync_comp_cycle_count_0_), .o(n_2932) );
na02s01 TIMEBOOST_cell_49489 ( .a(FE_OFN262_n_9851), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q), .o(TIMEBOOST_net_14962) );
in01f02 g63943_u3 ( .a(g63943_p), .o(n_2264) );
no02f10 g63944_u0 ( .a(n_3047), .b(n_1192), .o(n_3408) );
na02f20 g63947_u0 ( .a(n_2218), .b(n_6986), .o(n_4662) );
no02f06 g63948_u0 ( .a(n_2009), .b(n_1484), .o(n_2477) );
na02s01 TIMEBOOST_cell_18417 ( .a(FE_RN_122_0), .b(FE_OFN9_n_11877), .o(TIMEBOOST_net_5572) );
no02f06 g63950_u0 ( .a(n_1485), .b(n_2007), .o(n_2473) );
na02f04 g63951_u0 ( .a(n_2706), .b(wbm_adr_o_20_), .o(n_2707) );
na02f04 g63952_u0 ( .a(n_1643), .b(n_1009), .o(n_5769) );
na02f04 g63954_u0 ( .a(n_5230), .b(n_3077), .o(n_3407) );
na02m02 TIMEBOOST_cell_29547 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_408), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_8878) );
ao12f02 g63957_u0 ( .a(n_3071), .b(FE_OCPN1845_n_16427), .c(n_3404), .o(n_3406) );
na02f04 g63958_u0 ( .a(n_2840), .b(n_2621), .o(n_3302) );
na02f04 g63959_u0 ( .a(FE_OFN1944_n_15813), .b(n_2984), .o(n_3301) );
na02f04 TIMEBOOST_cell_18357 ( .a(n_3410), .b(FE_RN_158_0), .o(TIMEBOOST_net_5542) );
ao12f02 g63963_u0 ( .a(n_3042), .b(FE_OCPN1845_n_16427), .c(n_3078), .o(n_3403) );
na02s02 TIMEBOOST_cell_49288 ( .a(TIMEBOOST_net_14861), .b(TIMEBOOST_net_10890), .o(TIMEBOOST_net_9452) );
ao12s01 g63965_u0 ( .a(pci_target_unit_del_sync_req_comp_pending_sample), .b(n_3795), .c(g66433_sb), .o(n_4532) );
na02s02 TIMEBOOST_cell_48873 ( .a(FE_OFN252_n_9868), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q), .o(TIMEBOOST_net_14654) );
in01s01 TIMEBOOST_cell_73986 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .o(TIMEBOOST_net_23551) );
oa12f01 g63969_u0 ( .a(n_4084), .b(n_3386), .c(FE_OFN2121_n_2687), .o(n_4085) );
na02s01 TIMEBOOST_cell_37105 ( .a(TIMEBOOST_net_10164), .b(g61943_sb), .o(TIMEBOOST_net_575) );
ao22f04 g63976_u0 ( .a(n_1013), .b(n_1626), .c(n_2430), .d(wishbone_slave_unit_pci_initiator_if_current_byte_address_36), .o(n_2959) );
na02s01 TIMEBOOST_cell_28001 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q), .o(TIMEBOOST_net_8105) );
ao12f02 g63980_u0 ( .a(n_3084), .b(n_3372), .c(wbu_pref_en_in_137), .o(n_3399) );
ao12f10 g63981_u0 ( .a(FE_OFN1125_g64577_p), .b(n_980), .c(n_813), .o(n_4131) );
ao12f10 g63982_u0 ( .a(n_3119), .b(n_4718), .c(n_2344), .o(n_3120) );
na03s02 TIMEBOOST_cell_72557 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q), .b(FE_OFN587_n_9692), .c(TIMEBOOST_net_20607), .o(TIMEBOOST_net_17526) );
oa12f01 g63985_u0 ( .a(n_1488), .b(n_4904), .c(FE_OFN672_n_4505), .o(n_4918) );
oa12m02 g63986_u0 ( .a(n_2138), .b(n_4904), .c(FE_OFN665_n_4495), .o(n_4917) );
oa12f02 g63987_u0 ( .a(n_4510), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583), .c(FE_OFN1640_n_4671), .o(n_4915) );
oa12m02 g63988_u0 ( .a(n_1642), .b(n_4904), .c(FE_OFN634_n_4454), .o(n_4914) );
no02f01 g63989_u0 ( .a(n_1417), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_), .o(g63989_p) );
ao12f02 g63989_u1 ( .a(g63989_p), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_), .c(n_1417), .o(n_2262) );
oa12m02 g63990_u0 ( .a(n_1559), .b(n_4904), .c(FE_OFN614_n_4501), .o(n_4913) );
oa12f01 g63991_u0 ( .a(n_1555), .b(n_4904), .c(FE_OFN622_n_4409), .o(n_4912) );
oa12m02 g63992_u0 ( .a(n_1546), .b(n_4904), .c(FE_OFN659_n_4392), .o(n_4911) );
oa12m02 g63993_u0 ( .a(n_4513), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466), .c(n_4677), .o(n_4909) );
ao22f02 g63_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q), .b(n_15568), .c(n_15566), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q), .o(n_15529) );
in01f20 g64011_u0 ( .a(n_4743), .o(n_8440) );
oa12m02 g64016_u0 ( .a(n_1553), .b(n_4904), .c(FE_OFN648_n_4497), .o(n_4908) );
oa12m02 g64017_u0 ( .a(n_4511), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310), .c(FE_OFN1678_n_4655), .o(n_4907) );
oa12f01 g64018_u0 ( .a(n_2131), .b(n_4904), .c(n_4417), .o(n_4906) );
oa12f04 g64019_u0 ( .a(n_1547), .b(n_4904), .c(FE_OFN1623_n_4438), .o(n_4905) );
oa12m02 g64020_u0 ( .a(n_4509), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622), .c(FE_OFN651_n_4508), .o(n_4903) );
oa12m02 g64021_u0 ( .a(n_4514), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544), .c(n_4669), .o(n_4902) );
no02f02 g64022_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_), .b(n_1015), .o(g64022_p) );
ao12f01 g64022_u1 ( .a(g64022_p), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_), .c(n_1015), .o(n_1688) );
oa12m02 g64023_u0 ( .a(n_1537), .b(n_4904), .c(FE_OFN682_n_4460), .o(n_4901) );
oa12f01 g64024_u0 ( .a(n_1377), .b(n_4904), .c(FE_OFN1660_n_4490), .o(n_4900) );
na02m02 TIMEBOOST_cell_63323 ( .a(TIMEBOOST_net_20608), .b(g58071_sb), .o(TIMEBOOST_net_14943) );
ao22f04 g64027_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_486), .c(configuration_wb_err_addr_548), .d(n_15445), .o(n_2927) );
ao22f04 g64028_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_492), .c(n_16791), .d(pciu_bar0_in_370), .o(n_2926) );
ao22f02 g64029_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_487), .c(n_16791), .d(pciu_bar0_in_365), .o(n_2925) );
ao22f02 g64030_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_488), .c(n_16791), .d(pciu_bar0_in_366), .o(n_2924) );
ao22f04 g64031_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_473), .c(configuration_interrupt_line_39), .d(n_3295), .o(n_3297) );
ao22f02 g64033_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_471), .c(configuration_interrupt_line_37), .d(n_3295), .o(n_3296) );
ao22f02 g64034_u0 ( .a(n_3115), .b(configuration_icr_bit_2961), .c(configuration_wb_err_addr_533), .d(n_15444), .o(n_3117) );
ao22f06 g64035_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_493), .c(configuration_wb_err_addr_555), .d(n_15445), .o(n_2922) );
ao22f06 g64036_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_495), .c(n_3252), .d(configuration_pci_err_cs_bit_464), .o(n_2921) );
in01f02 g64038_u0 ( .a(n_15645), .o(n_4795) );
ao22f02 g64041_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_501), .c(n_3252), .d(configuration_pci_err_cs_bit_470), .o(n_2920) );
ao22f02 g64042_u0 ( .a(n_3115), .b(pci_resi_conf_soft_res_in), .c(configuration_wb_err_addr_563), .d(n_15444), .o(n_3116) );
ao22f02 g64043_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_505), .c(FE_OFN1006_n_16288), .d(configuration_pci_err_addr_474), .o(n_2919) );
ao22f02 g64044_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_508), .c(FE_OFN1006_n_16288), .d(configuration_pci_err_addr_477), .o(n_2918) );
na02s01 TIMEBOOST_cell_38220 ( .a(n_8511), .b(g65240_sb), .o(TIMEBOOST_net_10722) );
na03f02 TIMEBOOST_cell_66480 ( .a(TIMEBOOST_net_16778), .b(FE_OFN1311_n_6624), .c(g62446_sb), .o(n_6703) );
na03f02 TIMEBOOST_cell_66743 ( .a(TIMEBOOST_net_17163), .b(FE_OFN1260_n_4143), .c(g62467_sb), .o(n_6659) );
ao22f04 g64048_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_475), .c(configuration_interrupt_line_41), .d(n_3295), .o(n_3294) );
ao22f02 g64049_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_491), .c(n_16791), .d(pciu_bar0_in_369), .o(n_2917) );
ao22f02 g64050_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_476), .c(configuration_interrupt_line_42), .d(n_3295), .o(n_3393) );
in01f02 g64051_u0 ( .a(n_2916), .o(n_3114) );
ao22f04 g64052_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_500), .c(n_3252), .d(configuration_pci_err_cs_bit_469), .o(n_2916) );
na04f04 TIMEBOOST_cell_24211 ( .a(n_9519), .b(g57420_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q), .d(FE_OFN1419_n_8567), .o(n_11318) );
ao22f02 g64055_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_490), .c(n_16791), .d(pciu_bar0_in_368), .o(n_2913) );
na02f06 TIMEBOOST_cell_18550 ( .a(TIMEBOOST_net_5638), .b(n_2957), .o(n_4875) );
in01f02 g64060_u0 ( .a(n_2910), .o(n_3112) );
ao22f02 g64061_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_497), .c(n_3252), .d(configuration_pci_err_cs_bit_466), .o(n_2910) );
in01f02 g64062_u0 ( .a(n_2909), .o(n_3111) );
ao22f02 g64063_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_498), .c(n_3252), .d(configuration_pci_err_cs_bit_467), .o(n_2909) );
ao22f04 g64064_u0 ( .a(n_2699), .b(wbu_map_in_131), .c(n_2698), .d(wbu_map_in_132), .o(n_2700) );
ao22f02 g64065_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr), .c(configuration_wb_err_addr), .d(n_15445), .o(n_15435) );
ao22s02 g64066_u0 ( .a(n_2699), .b(wbu_pref_en_in_136), .c(n_2698), .d(wbu_pref_en_in_137), .o(n_2697) );
in01f02 g64067_u0 ( .a(n_2907), .o(n_3110) );
ao22f02 g64068_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_499), .c(n_3252), .d(configuration_pci_err_cs_bit_468), .o(n_2907) );
ao22f02 g64069_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_472), .c(configuration_interrupt_line_38), .d(n_3295), .o(n_3293) );
ao22f01 g64070_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_481), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_245), .o(n_2906) );
ao22s02 g64071_u0 ( .a(n_2699), .b(wbu_mrl_en_in_141), .c(n_2698), .d(wbu_mrl_en_in_142), .o(n_2696) );
ao22f04 g64072_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_482), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_246), .o(n_2905) );
ao22f02 g64073_u0 ( .a(n_3115), .b(configuration_icr_bit_2967), .c(configuration_wb_err_addr_534), .d(n_15444), .o(n_3109) );
ao22f01 g64074_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_483), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_247), .o(n_2904) );
ao22f01 g64075_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_484), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_248), .o(n_15434) );
ao22f02 g64076_u0 ( .a(FE_OFN1005_n_16288), .b(configuration_pci_err_addr_496), .c(n_3252), .d(configuration_pci_err_cs_bit_465), .o(n_2902) );
ao22f02 g64077_u0 ( .a(FE_OFN1006_n_16288), .b(configuration_pci_err_addr_485), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_249), .o(n_16852) );
in01m01 g64078_u0 ( .a(FE_OFN1077_n_4740), .o(g64078_sb) );
na02m01 TIMEBOOST_cell_68636 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q), .b(FE_OFN667_n_4495), .o(TIMEBOOST_net_21526) );
na02f01 g64078_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q), .b(FE_OFN1077_n_4740), .o(g64078_db) );
na03f10 TIMEBOOST_cell_68092 ( .a(n_2557), .b(wbs_stb_i), .c(n_3083), .o(TIMEBOOST_net_21254) );
in01m01 g64079_u0 ( .a(FE_OFN1046_n_16657), .o(g64079_sb) );
na02m01 TIMEBOOST_cell_53377 ( .a(n_2499), .b(pci_target_unit_pcit_if_strd_addr_in_688), .o(TIMEBOOST_net_16906) );
na02f01 g64079_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q), .b(FE_OFN1046_n_16657), .o(g64079_db) );
na02m10 TIMEBOOST_cell_45819 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q), .o(TIMEBOOST_net_13804) );
in01m04 g64080_u0 ( .a(FE_OFN1077_n_4740), .o(g64080_sb) );
na03f02 TIMEBOOST_cell_47296 ( .a(FE_OFN1736_n_16317), .b(FE_OFN1742_n_11019), .c(TIMEBOOST_net_13574), .o(n_12487) );
na03f02 TIMEBOOST_cell_47297 ( .a(FE_OFN1736_n_16317), .b(TIMEBOOST_net_13575), .c(FE_OFN1742_n_11019), .o(n_12492) );
in01m01 g64081_u0 ( .a(FE_OFN1075_n_4740), .o(g64081_sb) );
na02s02 TIMEBOOST_cell_48162 ( .a(TIMEBOOST_net_14298), .b(g58189_sb), .o(TIMEBOOST_net_10527) );
na02s01 TIMEBOOST_cell_31829 ( .a(n_16945), .b(n_4078), .o(TIMEBOOST_net_10019) );
in01f02 g64082_u0 ( .a(FE_OFN1077_n_4740), .o(g64082_sb) );
na02f02 TIMEBOOST_cell_49466 ( .a(TIMEBOOST_net_14950), .b(g63063_db), .o(TIMEBOOST_net_11362) );
na03f02 TIMEBOOST_cell_64476 ( .a(n_1802), .b(n_3334), .c(n_2410), .o(TIMEBOOST_net_276) );
in01m01 g64083_u0 ( .a(FE_OFN1076_n_4740), .o(g64083_sb) );
na02m02 TIMEBOOST_cell_29325 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q), .b(g64311_sb), .o(TIMEBOOST_net_8767) );
na02f01 g64083_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q), .b(FE_OFN1076_n_4740), .o(g64083_db) );
na02f02 TIMEBOOST_cell_44588 ( .a(TIMEBOOST_net_13188), .b(g63062_sb), .o(n_5126) );
in01m01 g64084_u0 ( .a(FE_OFN1077_n_4740), .o(g64084_sb) );
in01m01 g64085_u0 ( .a(FE_OFN906_n_4736), .o(g64085_sb) );
na02m01 g64085_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q), .b(FE_OFN906_n_4736), .o(g64085_db) );
na02f02 TIMEBOOST_cell_71445 ( .a(TIMEBOOST_net_22930), .b(n_3438), .o(n_4877) );
in01m01 g64086_u0 ( .a(FE_OFN1075_n_4740), .o(g64086_sb) );
na03f02 TIMEBOOST_cell_73519 ( .a(TIMEBOOST_net_13378), .b(n_6431), .c(g62363_sb), .o(n_6875) );
na02m02 TIMEBOOST_cell_71909 ( .a(TIMEBOOST_net_23162), .b(g65738_sb), .o(n_2056) );
in01m01 g64087_u0 ( .a(FE_OFN906_n_4736), .o(g64087_sb) );
na02m01 TIMEBOOST_cell_52443 ( .a(configuration_pci_err_data_509), .b(wbm_dat_o_8_), .o(TIMEBOOST_net_16439) );
na03f40 TIMEBOOST_cell_22024 ( .a(n_15735), .b(n_15736), .c(n_15739), .o(n_16486) );
in01m02 g64088_u0 ( .a(FE_OFN1075_n_4740), .o(g64088_sb) );
in01m06 g64089_u0 ( .a(FE_OFN1077_n_4740), .o(g64089_sb) );
na02s01 TIMEBOOST_cell_38988 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q), .b(g58328_sb), .o(TIMEBOOST_net_11106) );
in01s01 g64090_u0 ( .a(FE_OFN1046_n_16657), .o(g64090_sb) );
na02s01 TIMEBOOST_cell_53379 ( .a(n_2544), .b(pci_target_unit_pcit_if_strd_addr_in_690), .o(TIMEBOOST_net_16907) );
na02s01 g64090_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q), .b(FE_OFN1046_n_16657), .o(g64090_db) );
na03s06 TIMEBOOST_cell_70234 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q), .b(TIMEBOOST_net_16200), .c(g65800_sb), .o(TIMEBOOST_net_22325) );
in01m01 g64091_u0 ( .a(FE_OFN1051_n_16657), .o(g64091_sb) );
na03m02 TIMEBOOST_cell_72753 ( .a(TIMEBOOST_net_16203), .b(g65676_sb), .c(TIMEBOOST_net_22043), .o(TIMEBOOST_net_14802) );
na02s02 TIMEBOOST_cell_38549 ( .a(TIMEBOOST_net_10886), .b(g58197_db), .o(n_9589) );
na02m01 TIMEBOOST_cell_47807 ( .a(n_3747), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q), .o(TIMEBOOST_net_14121) );
in01m02 g64092_u0 ( .a(FE_OFN1075_n_4740), .o(g64092_sb) );
na03s02 TIMEBOOST_cell_65031 ( .a(g65733_db), .b(TIMEBOOST_net_6913), .c(TIMEBOOST_net_8197), .o(n_8417) );
na02s01 TIMEBOOST_cell_63840 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q), .o(TIMEBOOST_net_20906) );
na03m02 TIMEBOOST_cell_65479 ( .a(TIMEBOOST_net_20323), .b(g64168_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_13091) );
in01f01 g64093_u0 ( .a(FE_OFN1049_n_16657), .o(g64093_sb) );
na03m02 TIMEBOOST_cell_65603 ( .a(g64264_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q), .c(TIMEBOOST_net_12841), .o(TIMEBOOST_net_13050) );
na03f02 TIMEBOOST_cell_35061 ( .a(TIMEBOOST_net_10019), .b(FE_OFN1438_n_9372), .c(g58842_sb), .o(n_8672) );
na04m02 TIMEBOOST_cell_67320 ( .a(TIMEBOOST_net_12420), .b(n_4452), .c(g64828_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q), .o(TIMEBOOST_net_17537) );
in01f08 g64094_u0 ( .a(FE_OFN1074_n_4740), .o(g64094_sb) );
na02s02 TIMEBOOST_cell_49298 ( .a(TIMEBOOST_net_14866), .b(TIMEBOOST_net_12763), .o(TIMEBOOST_net_9421) );
na02f01 TIMEBOOST_cell_50006 ( .a(TIMEBOOST_net_15220), .b(n_4637), .o(n_4639) );
in01m04 g64095_u0 ( .a(FE_OFN905_n_4736), .o(g64095_sb) );
na02m08 TIMEBOOST_cell_45457 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q), .o(TIMEBOOST_net_13623) );
na02s02 TIMEBOOST_cell_39710 ( .a(g58447_sb), .b(FE_OFN203_n_9228), .o(TIMEBOOST_net_11467) );
in01m02 g64096_u0 ( .a(FE_OFN905_n_4736), .o(g64096_sb) );
na02f02 TIMEBOOST_cell_71621 ( .a(TIMEBOOST_net_23018), .b(FE_OFN1552_n_12104), .o(n_12784) );
na02s02 TIMEBOOST_cell_39712 ( .a(FE_OFN201_n_9230), .b(g58415_sb), .o(TIMEBOOST_net_11468) );
na02m01 TIMEBOOST_cell_62427 ( .a(TIMEBOOST_net_20160), .b(n_4730), .o(TIMEBOOST_net_14126) );
in01m01 g64097_u0 ( .a(FE_OFN1049_n_16657), .o(g64097_sb) );
na03f02 TIMEBOOST_cell_73520 ( .a(TIMEBOOST_net_17056), .b(n_6287), .c(g62905_sb), .o(n_6067) );
na02f02 TIMEBOOST_cell_54306 ( .a(TIMEBOOST_net_17370), .b(FE_OFN1194_n_6935), .o(TIMEBOOST_net_15434) );
in01m01 g64098_u0 ( .a(FE_OFN1049_n_16657), .o(g64098_sb) );
na04f02 TIMEBOOST_cell_67590 ( .a(TIMEBOOST_net_13837), .b(g62118_sb), .c(configuration_wb_err_addr_549), .d(FE_OFN1170_n_5592), .o(n_5578) );
in01s01 TIMEBOOST_cell_73987 ( .a(TIMEBOOST_net_23551), .o(TIMEBOOST_net_23552) );
in01m02 g64099_u0 ( .a(FE_OFN1049_n_16657), .o(g64099_sb) );
na02m02 TIMEBOOST_cell_49764 ( .a(TIMEBOOST_net_15099), .b(g61917_sb), .o(n_7987) );
na02m04 TIMEBOOST_cell_68681 ( .a(TIMEBOOST_net_21548), .b(TIMEBOOST_net_14292), .o(TIMEBOOST_net_13361) );
na02m02 TIMEBOOST_cell_54710 ( .a(TIMEBOOST_net_17572), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_15367) );
in01m01 g64100_u0 ( .a(FE_OFN1076_n_4740), .o(g64100_sb) );
na03f02 TIMEBOOST_cell_73730 ( .a(TIMEBOOST_net_13614), .b(FE_OFN2209_n_11027), .c(FE_OFN1752_n_12086), .o(n_12766) );
na03f02 TIMEBOOST_cell_68038 ( .a(FE_OFN1774_n_13800), .b(TIMEBOOST_net_13708), .c(FE_OFN1770_n_14054), .o(n_14479) );
oa12m02 g64101_u0 ( .a(n_1815), .b(FE_OFN923_n_4740), .c(pci_target_unit_fifos_pciw_control_in), .o(n_4528) );
in01m02 g64102_u0 ( .a(FE_OFN905_n_4736), .o(g64102_sb) );
na02s02 TIMEBOOST_cell_39714 ( .a(FE_OFN203_n_9228), .b(g58416_sb), .o(TIMEBOOST_net_11469) );
na03f02 TIMEBOOST_cell_66472 ( .a(TIMEBOOST_net_20588), .b(FE_OFN1274_n_4096), .c(g62557_sb), .o(n_6448) );
na02m01 TIMEBOOST_cell_70336 ( .a(TIMEBOOST_net_17290), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_22376) );
in01m04 g64103_u0 ( .a(FE_OFN1076_n_4740), .o(g64103_sb) );
na03f02 TIMEBOOST_cell_67950 ( .a(TIMEBOOST_net_13107), .b(FE_OFN1132_g64577_p), .c(g63169_sb), .o(n_4955) );
na03f02 TIMEBOOST_cell_66214 ( .a(TIMEBOOST_net_13235), .b(FE_OFN1224_n_6391), .c(g62583_sb), .o(n_6386) );
na02s01 TIMEBOOST_cell_70870 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q), .o(TIMEBOOST_net_22643) );
oa12f01 g64104_u0 ( .a(n_1795), .b(FE_OFN1046_n_16657), .c(pci_target_unit_fifos_pciw_control_in), .o(n_4527) );
in01m01 g64105_u0 ( .a(FE_OFN904_n_4736), .o(g64105_sb) );
na02s02 TIMEBOOST_cell_39716 ( .a(g58412_sb), .b(FE_OFN201_n_9230), .o(TIMEBOOST_net_11470) );
na03f02 TIMEBOOST_cell_34801 ( .a(TIMEBOOST_net_9551), .b(FE_OFN1381_n_8567), .c(g57279_sb), .o(n_10413) );
in01m01 g64106_u0 ( .a(FE_OFN1046_n_16657), .o(g64106_sb) );
na02m02 TIMEBOOST_cell_50300 ( .a(TIMEBOOST_net_15367), .b(g62602_sb), .o(n_6347) );
na02m02 g64106_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q), .b(FE_OFN1046_n_16657), .o(g64106_db) );
na02f02 TIMEBOOST_cell_54708 ( .a(TIMEBOOST_net_17571), .b(FE_OFN1261_n_4143), .o(TIMEBOOST_net_15501) );
in01m02 g64107_u0 ( .a(FE_OFN1049_n_16657), .o(g64107_sb) );
na02m02 TIMEBOOST_cell_63919 ( .a(TIMEBOOST_net_20945), .b(g58365_sb), .o(n_9210) );
na03s01 TIMEBOOST_cell_35790 ( .a(g58330_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q), .c(g58330_db), .o(n_9215) );
na02m01 TIMEBOOST_cell_53978 ( .a(TIMEBOOST_net_17206), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_14175) );
in01m08 g64108_u0 ( .a(FE_OFN1046_n_16657), .o(g64108_sb) );
in01s01 TIMEBOOST_cell_45933 ( .a(TIMEBOOST_net_13955), .o(TIMEBOOST_net_13894) );
na03f02 TIMEBOOST_cell_73128 ( .a(TIMEBOOST_net_12854), .b(g64079_sb), .c(g64079_db), .o(TIMEBOOST_net_15176) );
in01s01 TIMEBOOST_cell_45934 ( .a(TIMEBOOST_net_13894), .o(TIMEBOOST_net_13895) );
in01m01 g64109_u0 ( .a(FE_OFN1076_n_4740), .o(g64109_sb) );
na02f02 TIMEBOOST_cell_40831 ( .a(TIMEBOOST_net_12027), .b(FE_OFN1575_n_12028), .o(n_12720) );
na02f02 TIMEBOOST_cell_71044 ( .a(FE_OFN1265_n_4095), .b(TIMEBOOST_net_17010), .o(TIMEBOOST_net_22730) );
na02s01 TIMEBOOST_cell_68508 ( .a(n_2526), .b(g66398_sb), .o(TIMEBOOST_net_21462) );
in01m08 g64110_u0 ( .a(FE_OFN1046_n_16657), .o(g64110_sb) );
no02f08 TIMEBOOST_cell_29461 ( .a(FE_OFN969_n_13784), .b(FE_RN_559_0), .o(TIMEBOOST_net_8835) );
na03f02 TIMEBOOST_cell_72864 ( .a(TIMEBOOST_net_21720), .b(g65400_sb), .c(TIMEBOOST_net_22104), .o(TIMEBOOST_net_20519) );
in01f08 g64111_u0 ( .a(FE_OFN1074_n_4740), .o(g64111_sb) );
na02m04 TIMEBOOST_cell_69030 ( .a(g65319_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q), .o(TIMEBOOST_net_21723) );
na02s02 TIMEBOOST_cell_68908 ( .a(g65743_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q), .o(TIMEBOOST_net_21662) );
in01m04 g64112_u0 ( .a(FE_OFN1077_n_4740), .o(g64112_sb) );
na02m02 TIMEBOOST_cell_49172 ( .a(TIMEBOOST_net_14803), .b(g61774_sb), .o(n_8260) );
na04f04 TIMEBOOST_cell_73063 ( .a(n_1895), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q), .c(FE_OFN710_n_8232), .d(g61876_sb), .o(n_8079) );
in01m01 g64113_u0 ( .a(FE_OFN1046_n_16657), .o(g64113_sb) );
na02s02 TIMEBOOST_cell_48874 ( .a(TIMEBOOST_net_14654), .b(g58136_sb), .o(TIMEBOOST_net_10856) );
na02m01 TIMEBOOST_cell_68331 ( .a(TIMEBOOST_net_21373), .b(g65377_sb), .o(TIMEBOOST_net_12347) );
na02s02 TIMEBOOST_cell_37245 ( .a(TIMEBOOST_net_10234), .b(g65719_sb), .o(n_2066) );
in01m02 g64114_u0 ( .a(FE_OFN937_n_2292), .o(g64114_sb) );
na03f02 TIMEBOOST_cell_34861 ( .a(TIMEBOOST_net_9510), .b(FE_OFN1383_n_8567), .c(g57416_sb), .o(n_11326) );
na03f02 TIMEBOOST_cell_66307 ( .a(TIMEBOOST_net_13375), .b(n_6232), .c(g62978_sb), .o(n_5926) );
in01m06 g64115_u0 ( .a(FE_OFN1076_n_4740), .o(g64115_sb) );
na02f02 TIMEBOOST_cell_70631 ( .a(TIMEBOOST_net_22523), .b(g63068_sb), .o(n_5114) );
na04m02 TIMEBOOST_cell_67866 ( .a(n_3744), .b(g65087_sb), .c(FE_OFN662_n_4392), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q), .o(n_3598) );
na02s02 TIMEBOOST_cell_71421 ( .a(TIMEBOOST_net_22918), .b(TIMEBOOST_net_20514), .o(TIMEBOOST_net_14532) );
in01m01 g64116_u0 ( .a(FE_OFN1049_n_16657), .o(g64116_sb) );
na02m10 TIMEBOOST_cell_29465 ( .a(configuration_pci_err_data_507), .b(wbm_dat_o_6_), .o(TIMEBOOST_net_8837) );
na02f01 g64116_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN1049_n_16657), .o(g64116_db) );
na02f01 TIMEBOOST_cell_48016 ( .a(TIMEBOOST_net_14225), .b(FE_OFN1010_n_4734), .o(TIMEBOOST_net_12613) );
in01f02 g64117_u0 ( .a(FE_OFN1075_n_4740), .o(g64117_sb) );
in01m01 g64118_u0 ( .a(FE_OFN908_n_4734), .o(g64118_sb) );
na03m04 TIMEBOOST_cell_72845 ( .a(g65062_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q), .c(TIMEBOOST_net_16243), .o(TIMEBOOST_net_20974) );
na02s02 TIMEBOOST_cell_62466 ( .a(g58123_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q), .o(TIMEBOOST_net_20180) );
in01m02 g64119_u0 ( .a(FE_OFN906_n_4736), .o(g64119_sb) );
na03f02 TIMEBOOST_cell_66915 ( .a(FE_OFN1733_n_16317), .b(TIMEBOOST_net_16488), .c(FE_OFN1738_n_11019), .o(n_12634) );
na02f02 TIMEBOOST_cell_71017 ( .a(TIMEBOOST_net_22716), .b(g62375_sb), .o(n_6853) );
na02s01 TIMEBOOST_cell_39720 ( .a(FE_OFN201_n_9230), .b(g58410_sb), .o(TIMEBOOST_net_11472) );
in01m01 g64120_u0 ( .a(FE_OFN904_n_4736), .o(g64120_sb) );
na03f02 TIMEBOOST_cell_34847 ( .a(TIMEBOOST_net_9428), .b(FE_OFN1390_n_8567), .c(g57355_sb), .o(n_11393) );
na02f02 TIMEBOOST_cell_70099 ( .a(TIMEBOOST_net_22257), .b(FE_OFN1092_g64577_p), .o(TIMEBOOST_net_15192) );
oa12m02 g64121_u0 ( .a(n_1804), .b(FE_OFN903_n_4736), .c(pci_target_unit_fifos_pciw_control_in), .o(n_4524) );
in01m02 g64122_u0 ( .a(FE_OFN902_n_4736), .o(g64122_sb) );
na03f02 TIMEBOOST_cell_35131 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q), .b(n_13617), .c(g54489_da), .o(n_13607) );
na03m04 TIMEBOOST_cell_72490 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q), .b(n_3749), .c(TIMEBOOST_net_22073), .o(TIMEBOOST_net_17079) );
in01m02 g64123_u0 ( .a(FE_OFN904_n_4736), .o(g64123_sb) );
na02s01 TIMEBOOST_cell_39722 ( .a(FE_OFN203_n_9228), .b(g58411_sb), .o(TIMEBOOST_net_11473) );
na02m02 TIMEBOOST_cell_50404 ( .a(TIMEBOOST_net_15419), .b(g63149_sb), .o(n_5842) );
no02m04 g64124_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .b(n_1176), .o(g64124_p) );
ao12m02 g64124_u1 ( .a(g64124_p), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .c(n_1176), .o(n_1750) );
in01m04 g64125_u0 ( .a(FE_OFN923_n_4740), .o(g64125_sb) );
na03f02 TIMEBOOST_cell_73703 ( .a(TIMEBOOST_net_13511), .b(FE_OFN1762_n_10780), .c(FE_OFN1583_n_12306), .o(n_12625) );
na03f02 TIMEBOOST_cell_69032 ( .a(TIMEBOOST_net_20251), .b(FE_OFN1012_n_4734), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q), .o(TIMEBOOST_net_21724) );
in01m02 g64126_u0 ( .a(FE_OFN905_n_4736), .o(g64126_sb) );
na02s02 TIMEBOOST_cell_39724 ( .a(g57906_sb), .b(FE_OFN201_n_9230), .o(TIMEBOOST_net_11474) );
in01s01 TIMEBOOST_cell_67719 ( .a(pci_target_unit_fifos_pcir_data_in_159), .o(TIMEBOOST_net_21146) );
na03s02 TIMEBOOST_cell_66253 ( .a(TIMEBOOST_net_14167), .b(n_8272), .c(g61930_sb), .o(n_7963) );
in01m01 g64127_u0 ( .a(FE_OFN1049_n_16657), .o(g64127_sb) );
na02f03 TIMEBOOST_cell_29467 ( .a(configuration_pci_err_data_502), .b(wbm_dat_o_1_), .o(TIMEBOOST_net_8838) );
na02f01 TIMEBOOST_cell_48018 ( .a(TIMEBOOST_net_14226), .b(FE_OFN1011_n_4734), .o(TIMEBOOST_net_10569) );
in01m01 g64128_u0 ( .a(FE_OFN905_n_4736), .o(g64128_sb) );
na02s02 TIMEBOOST_cell_39726 ( .a(g57907_sb), .b(FE_OFN203_n_9228), .o(TIMEBOOST_net_11475) );
na03f08 TIMEBOOST_cell_65315 ( .a(TIMEBOOST_net_14564), .b(n_3335), .c(n_8566), .o(n_8819) );
na02s01 TIMEBOOST_cell_30993 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_0__Q), .b(FE_OFN207_n_9865), .o(TIMEBOOST_net_9601) );
in01m02 g64129_u0 ( .a(FE_OFN1010_n_4734), .o(g64129_sb) );
na02s01 TIMEBOOST_cell_39728 ( .a(g57901_sb), .b(FE_OFN203_n_9228), .o(TIMEBOOST_net_11476) );
no03f08 TIMEBOOST_cell_22388 ( .a(n_4165), .b(n_16168), .c(TIMEBOOST_net_583), .o(n_5722) );
na02m10 TIMEBOOST_cell_45801 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q), .o(TIMEBOOST_net_13795) );
in01m04 g64130_u0 ( .a(FE_OFN1013_n_4734), .o(g64130_sb) );
na03f02 TIMEBOOST_cell_66730 ( .a(TIMEBOOST_net_16829), .b(FE_OFN1305_n_13124), .c(g54360_sb), .o(n_13082) );
na02f01 TIMEBOOST_cell_62465 ( .a(TIMEBOOST_net_20179), .b(FE_OFN905_n_4736), .o(TIMEBOOST_net_14141) );
na02f01 TIMEBOOST_cell_43913 ( .a(TIMEBOOST_net_10977), .b(n_12595), .o(TIMEBOOST_net_12851) );
in01m10 g64131_u0 ( .a(FE_OFN1046_n_16657), .o(g64131_sb) );
na02f03 TIMEBOOST_cell_29469 ( .a(configuration_pci_err_data_503), .b(wbm_dat_o_2_), .o(TIMEBOOST_net_8839) );
na02s02 TIMEBOOST_cell_49490 ( .a(TIMEBOOST_net_14962), .b(FE_OFN580_n_9531), .o(TIMEBOOST_net_11197) );
na02f01 TIMEBOOST_cell_48020 ( .a(TIMEBOOST_net_14227), .b(FE_OFN1011_n_4734), .o(TIMEBOOST_net_10571) );
in01m01 g64132_u0 ( .a(FE_OFN908_n_4734), .o(g64132_sb) );
na02m01 TIMEBOOST_cell_42904 ( .a(TIMEBOOST_net_12346), .b(g60689_sb), .o(n_3815) );
in01m01 g64133_u0 ( .a(FE_OFN1046_n_16657), .o(g64133_sb) );
na02f03 TIMEBOOST_cell_29471 ( .a(configuration_pci_err_addr_471), .b(wbm_adr_o_1_), .o(TIMEBOOST_net_8840) );
na02s01 TIMEBOOST_cell_68182 ( .a(TIMEBOOST_net_10153), .b(n_2299), .o(TIMEBOOST_net_21299) );
na02s02 TIMEBOOST_cell_48022 ( .a(TIMEBOOST_net_14228), .b(g58167_sb), .o(TIMEBOOST_net_10381) );
in01f01 g64134_u0 ( .a(FE_OFN1049_n_16657), .o(g64134_sb) );
na03m04 TIMEBOOST_cell_72848 ( .a(g64868_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q), .c(TIMEBOOST_net_10581), .o(TIMEBOOST_net_17072) );
na02f01 g64134_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q), .b(FE_OFN1049_n_16657), .o(g64134_db) );
na02m01 TIMEBOOST_cell_48201 ( .a(n_26), .b(FE_OFN662_n_4392), .o(TIMEBOOST_net_14318) );
in01m01 g64135_u0 ( .a(FE_OFN906_n_4736), .o(g64135_sb) );
na02f01 g64135_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q), .b(FE_OFN906_n_4736), .o(g64135_db) );
na02f01 TIMEBOOST_cell_47575 ( .a(n_1679), .b(n_1415), .o(TIMEBOOST_net_14005) );
in01m02 g64136_u0 ( .a(FE_OFN1076_n_4740), .o(g64136_sb) );
na03m02 TIMEBOOST_cell_69044 ( .a(FE_OFN1640_n_4671), .b(g65323_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q), .o(TIMEBOOST_net_21730) );
na02s02 TIMEBOOST_cell_38809 ( .a(TIMEBOOST_net_11016), .b(g65892_sb), .o(n_2582) );
in01m04 g64137_u0 ( .a(FE_OFN1049_n_16657), .o(g64137_sb) );
na02m80 TIMEBOOST_cell_29473 ( .a(configuration_pci_err_cs_bit31_24), .b(pci_target_unit_wishbone_master_bc_register_reg_0__Q), .o(TIMEBOOST_net_8841) );
na02f02 TIMEBOOST_cell_49160 ( .a(TIMEBOOST_net_14797), .b(g61944_sb), .o(n_7937) );
in01s01 g64138_u0 ( .a(FE_OFN904_n_4736), .o(g64138_sb) );
na02m01 TIMEBOOST_cell_53455 ( .a(TIMEBOOST_net_12852), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q), .o(TIMEBOOST_net_16945) );
na02s01 TIMEBOOST_cell_45407 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q), .o(TIMEBOOST_net_13598) );
na02s02 TIMEBOOST_cell_39730 ( .a(g57898_sb), .b(FE_OFN203_n_9228), .o(TIMEBOOST_net_11477) );
in01m01 g64139_u0 ( .a(FE_OFN905_n_4736), .o(g64139_sb) );
na02m10 TIMEBOOST_cell_52269 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_138), .o(TIMEBOOST_net_16352) );
na02f01 g64139_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q), .b(FE_OFN905_n_4736), .o(g64139_db) );
in01m02 g64140_u0 ( .a(FE_OFN923_n_4740), .o(g64140_sb) );
na02m04 TIMEBOOST_cell_68992 ( .a(FE_OFN653_n_4508), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q), .o(TIMEBOOST_net_21704) );
na02s02 TIMEBOOST_cell_38795 ( .a(TIMEBOOST_net_11009), .b(g65892_sb), .o(n_2587) );
in01m02 g64141_u0 ( .a(FE_OFN906_n_4736), .o(g64141_sb) );
na03f02 TIMEBOOST_cell_34930 ( .a(TIMEBOOST_net_9520), .b(FE_OFN1368_n_8567), .c(g57330_sb), .o(n_10397) );
na03f06 TIMEBOOST_cell_73704 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q), .b(FE_OFN1747_n_12004), .c(TIMEBOOST_net_20691), .o(TIMEBOOST_net_478) );
in01s02 g64142_u0 ( .a(FE_OFN953_n_2055), .o(g64142_sb) );
na02m01 TIMEBOOST_cell_62464 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_130), .o(TIMEBOOST_net_20179) );
na02m02 TIMEBOOST_cell_68645 ( .a(TIMEBOOST_net_21530), .b(g64791_sb), .o(TIMEBOOST_net_8679) );
in01m02 g64143_u0 ( .a(FE_OFN908_n_4734), .o(g64143_sb) );
na02m01 TIMEBOOST_cell_71966 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q), .o(TIMEBOOST_net_23191) );
na03m08 TIMEBOOST_cell_72534 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q), .b(g58022_sb), .c(TIMEBOOST_net_10616), .o(TIMEBOOST_net_16842) );
in01m01 g64144_u0 ( .a(FE_OFN1013_n_4734), .o(g64144_sb) );
na02f02 TIMEBOOST_cell_71748 ( .a(TIMEBOOST_net_13792), .b(n_13903), .o(TIMEBOOST_net_23082) );
in01s01 g64145_u0 ( .a(FE_OFN2109_n_2047), .o(g64145_sb) );
na02s02 TIMEBOOST_cell_49289 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q), .b(FE_OFN526_n_9899), .o(TIMEBOOST_net_14862) );
na03f02 TIMEBOOST_cell_73633 ( .a(TIMEBOOST_net_20521), .b(FE_OFN1216_n_4151), .c(g63150_sb), .o(n_5840) );
na02s06 TIMEBOOST_cell_43091 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q), .b(pci_target_unit_fifos_pcir_data_in_188), .o(TIMEBOOST_net_12440) );
in01f01 g64146_u0 ( .a(FE_OFN1010_n_4734), .o(g64146_sb) );
in01m02 g64147_u0 ( .a(FE_OFN906_n_4736), .o(g64147_sb) );
na03f06 TIMEBOOST_cell_73577 ( .a(TIMEBOOST_net_7607), .b(FE_OFN1085_n_13221), .c(g54176_da), .o(TIMEBOOST_net_22879) );
na03s02 TIMEBOOST_cell_72640 ( .a(TIMEBOOST_net_21416), .b(n_8272), .c(g61949_sb), .o(n_7927) );
in01m01 g64148_u0 ( .a(FE_OFN906_n_4736), .o(g64148_sb) );
na02m10 TIMEBOOST_cell_52657 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q), .o(TIMEBOOST_net_16546) );
na03f02 TIMEBOOST_cell_34931 ( .a(TIMEBOOST_net_9491), .b(FE_OFN1413_n_8567), .c(g57266_sb), .o(n_10418) );
in01m01 g64149_u0 ( .a(FE_OFN1074_n_4740), .o(g64149_sb) );
na02m02 TIMEBOOST_cell_53973 ( .a(pci_target_unit_fifos_pciw_cbe_in_153), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q), .o(TIMEBOOST_net_17204) );
na02s01 TIMEBOOST_cell_53530 ( .a(TIMEBOOST_net_16982), .b(TIMEBOOST_net_12480), .o(TIMEBOOST_net_9325) );
in01f01 g64150_u0 ( .a(FE_OFN1011_n_4734), .o(g64150_sb) );
na02m02 TIMEBOOST_cell_68957 ( .a(TIMEBOOST_net_21686), .b(TIMEBOOST_net_16239), .o(TIMEBOOST_net_17446) );
na03f02 TIMEBOOST_cell_34824 ( .a(TIMEBOOST_net_9345), .b(FE_OFN1407_n_8567), .c(g57288_sb), .o(n_11464) );
na03f10 TIMEBOOST_cell_32069 ( .a(n_2458), .b(n_2982), .c(n_2457), .o(n_2459) );
in01f01 g64151_u0 ( .a(FE_OFN1011_n_4734), .o(g64151_sb) );
na02m01 TIMEBOOST_cell_38044 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q), .b(FE_OFN1660_n_4490), .o(TIMEBOOST_net_10634) );
na02f01 g64151_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q), .b(FE_OFN1011_n_4734), .o(g64151_db) );
in01m01 g64152_u0 ( .a(FE_OFN1010_n_4734), .o(g64152_sb) );
na02m02 TIMEBOOST_cell_69218 ( .a(g65398_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q), .o(TIMEBOOST_net_21817) );
na02s01 TIMEBOOST_cell_45361 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q), .o(TIMEBOOST_net_13575) );
in01m01 g64153_u0 ( .a(FE_OFN1013_n_4734), .o(g64153_sb) );
na03m04 TIMEBOOST_cell_72927 ( .a(g65282_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q), .c(TIMEBOOST_net_16293), .o(TIMEBOOST_net_20521) );
na03f02 TIMEBOOST_cell_34826 ( .a(TIMEBOOST_net_9346), .b(FE_OFN1383_n_8567), .c(g57157_sb), .o(n_11593) );
na04f02 TIMEBOOST_cell_67924 ( .a(n_9), .b(g60409_sb), .c(n_2234), .d(n_7078), .o(n_4859) );
in01f01 g64154_u0 ( .a(FE_OFN1010_n_4734), .o(g64154_sb) );
na02s02 TIMEBOOST_cell_49994 ( .a(TIMEBOOST_net_15214), .b(g58442_sb), .o(n_8993) );
na04f02 TIMEBOOST_cell_66093 ( .a(n_3390), .b(n_3052), .c(n_3259), .d(n_3229), .o(n_4786) );
na02s01 TIMEBOOST_cell_48715 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q), .b(FE_OFN587_n_9692), .o(TIMEBOOST_net_14575) );
in01f02 g64155_u0 ( .a(FE_OFN1010_n_4734), .o(g64155_sb) );
na02m02 TIMEBOOST_cell_30857 ( .a(n_9490), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q), .o(TIMEBOOST_net_9533) );
na03f02 TIMEBOOST_cell_70774 ( .a(n_2271), .b(FE_OFN1697_n_5751), .c(wbm_adr_o_5_), .o(TIMEBOOST_net_22595) );
in01m01 g64156_u0 ( .a(FE_OFN1012_n_4734), .o(g64156_sb) );
na03f02 TIMEBOOST_cell_44347 ( .a(g65905_da), .b(g65905_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q), .o(TIMEBOOST_net_13068) );
in01m01 g64157_u0 ( .a(FE_OFN1075_n_4740), .o(g64157_sb) );
na03s01 TIMEBOOST_cell_41746 ( .a(g58336_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q), .c(g58336_db), .o(n_9020) );
in01m01 g64158_u0 ( .a(FE_OFN1011_n_4734), .o(g64158_sb) );
na02f10 TIMEBOOST_cell_49067 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_780), .o(TIMEBOOST_net_14751) );
na03f02 TIMEBOOST_cell_34828 ( .a(TIMEBOOST_net_9338), .b(FE_OFN1420_n_8567), .c(g57514_sb), .o(n_11228) );
in01f01 g64159_u0 ( .a(FE_OFN1013_n_4734), .o(g64159_sb) );
na02f02 TIMEBOOST_cell_71003 ( .a(TIMEBOOST_net_22709), .b(g62515_sb), .o(n_6548) );
na02m02 TIMEBOOST_cell_48792 ( .a(TIMEBOOST_net_14613), .b(TIMEBOOST_net_11081), .o(TIMEBOOST_net_9375) );
na02f02 TIMEBOOST_cell_38269 ( .a(TIMEBOOST_net_10746), .b(g65972_sb), .o(n_2152) );
in01f01 g64160_u0 ( .a(FE_OFN1010_n_4734), .o(g64160_sb) );
na02f01 g64160_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q), .b(FE_OFN1010_n_4734), .o(g64160_db) );
na04f04 TIMEBOOST_cell_23322 ( .a(wbm_adr_o_9_), .b(g59800_sb), .c(g59800_db), .d(g52455_sb), .o(g52455_da) );
in01m01 g64161_u0 ( .a(FE_OFN1011_n_4734), .o(g64161_sb) );
na03f02 TIMEBOOST_cell_73634 ( .a(TIMEBOOST_net_17482), .b(n_6645), .c(g62540_sb), .o(n_6488) );
in01f01 g64162_u0 ( .a(FE_OFN908_n_4734), .o(g64162_sb) );
na03f02 TIMEBOOST_cell_69966 ( .a(FE_OCPUNCON1952_FE_OFN697_n_16760), .b(pci_target_unit_pcit_if_strd_addr_in_711), .c(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75), .o(TIMEBOOST_net_22191) );
na02m01 g52463_u1 ( .a(wbs_adr_i_17_), .b(g52463_sb), .o(g52463_da) );
na02m10 TIMEBOOST_cell_52987 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q), .b(wishbone_slave_unit_pcim_sm_data_in_639), .o(TIMEBOOST_net_16711) );
in01f02 g64163_u0 ( .a(FE_OFN1011_n_4734), .o(g64163_sb) );
na02f02 TIMEBOOST_cell_54318 ( .a(TIMEBOOST_net_17376), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_15706) );
na02m02 TIMEBOOST_cell_54731 ( .a(g58127_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q), .o(TIMEBOOST_net_17583) );
in01m01 g64164_u0 ( .a(FE_OFN1010_n_4734), .o(g64164_sb) );
na03f02 TIMEBOOST_cell_34830 ( .a(TIMEBOOST_net_9339), .b(FE_OFN1404_n_8567), .c(g57393_sb), .o(n_11349) );
in01m01 g64165_u0 ( .a(FE_OFN1074_n_4740), .o(g64165_sb) );
na02s02 TIMEBOOST_cell_49444 ( .a(TIMEBOOST_net_14939), .b(g58147_db), .o(n_9647) );
na02s01 TIMEBOOST_cell_51669 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q), .o(TIMEBOOST_net_16052) );
in01s01 TIMEBOOST_cell_45942 ( .a(TIMEBOOST_net_13902), .o(TIMEBOOST_net_13903) );
in01m02 g64166_u0 ( .a(FE_OFN1013_n_4734), .o(g64166_sb) );
na04f04 TIMEBOOST_cell_67690 ( .a(TIMEBOOST_net_16858), .b(FE_OFN2198_n_10256), .c(g52595_sb), .d(TIMEBOOST_net_702), .o(n_11878) );
na03f02 TIMEBOOST_cell_34832 ( .a(TIMEBOOST_net_9384), .b(FE_OFN1381_n_8567), .c(g57375_sb), .o(n_10380) );
na02s01 TIMEBOOST_cell_45265 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q), .o(TIMEBOOST_net_13527) );
in01m01 g64167_u0 ( .a(FE_OFN905_n_4736), .o(g64167_sb) );
na02s02 TIMEBOOST_cell_52229 ( .a(g58118_sb), .b(FE_OFN221_n_9846), .o(TIMEBOOST_net_16332) );
na02m01 g64167_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q), .b(FE_OFN905_n_4736), .o(g64167_db) );
in01s01 TIMEBOOST_cell_73859 ( .a(TIMEBOOST_net_23423), .o(TIMEBOOST_net_23424) );
in01m01 g64168_u0 ( .a(FE_OFN1012_n_4734), .o(g64168_sb) );
na02s01 TIMEBOOST_cell_43165 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q), .o(TIMEBOOST_net_12477) );
na03f02 TIMEBOOST_cell_72870 ( .a(n_2566), .b(FE_OFN989_n_574), .c(TIMEBOOST_net_8654), .o(n_2567) );
in01m01 g64169_u0 ( .a(FE_OFN906_n_4736), .o(g64169_sb) );
na02s01 TIMEBOOST_cell_62536 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q), .o(TIMEBOOST_net_20215) );
na04f04 TIMEBOOST_cell_68005 ( .a(g54180_db), .b(FE_OFN1000_n_15978), .c(TIMEBOOST_net_13391), .d(g54180_sb), .o(TIMEBOOST_net_20594) );
in01m02 g64170_u0 ( .a(FE_OFN923_n_4740), .o(g64170_sb) );
na04f01 TIMEBOOST_cell_67811 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q), .b(FE_OFN601_n_9687), .c(FE_OFN211_n_9858), .d(g58110_sb), .o(n_9684) );
in01f01 g64171_u0 ( .a(FE_OFN1010_n_4734), .o(g64171_sb) );
na02s02 TIMEBOOST_cell_39732 ( .a(FE_OFN203_n_9228), .b(g57895_sb), .o(TIMEBOOST_net_11478) );
na02m10 TIMEBOOST_cell_45805 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q), .o(TIMEBOOST_net_13797) );
in01s01 g64172_u0 ( .a(FE_OFN904_n_4736), .o(g64172_sb) );
na03s02 TIMEBOOST_cell_67826 ( .a(FE_OFN525_n_9899), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q), .c(g58011_sb), .o(TIMEBOOST_net_14533) );
na02m10 TIMEBOOST_cell_53021 ( .a(configuration_pci_err_data_521), .b(wbm_dat_o_20_), .o(TIMEBOOST_net_16728) );
na03f06 TIMEBOOST_cell_22054 ( .a(n_15908), .b(FE_OCP_RBN2221_n_15347), .c(n_319), .o(g74563_p) );
in01m01 g64173_u0 ( .a(FE_OFN1050_n_16657), .o(g64173_sb) );
na02f03 TIMEBOOST_cell_29475 ( .a(configuration_pci_err_addr), .b(wbm_adr_o_0_), .o(TIMEBOOST_net_8842) );
na02f02 TIMEBOOST_cell_71387 ( .a(TIMEBOOST_net_22901), .b(g59111_sb), .o(n_8707) );
oa12f01 g64174_u0 ( .a(n_1803), .b(FE_OFN1012_n_4734), .c(pci_target_unit_fifos_pciw_control_in), .o(n_4521) );
in01m02 g64175_u0 ( .a(FE_OFN1013_n_4734), .o(g64175_sb) );
na03f02 TIMEBOOST_cell_73440 ( .a(TIMEBOOST_net_20967), .b(FE_OFN1294_n_4098), .c(g62897_sb), .o(n_6083) );
in01m02 g64176_u0 ( .a(FE_OFN1012_n_4734), .o(g64176_sb) );
na02f02 TIMEBOOST_cell_63989 ( .a(TIMEBOOST_net_20980), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_15689) );
na03f02 TIMEBOOST_cell_34932 ( .a(TIMEBOOST_net_9521), .b(FE_OFN1400_n_8567), .c(g57136_sb), .o(n_11614) );
in01m02 g64177_u0 ( .a(FE_OFN906_n_4736), .o(g64177_sb) );
na03m02 TIMEBOOST_cell_68010 ( .a(TIMEBOOST_net_14947), .b(FE_OFN272_n_9828), .c(TIMEBOOST_net_15085), .o(TIMEBOOST_net_9410) );
in01m01 g64178_u0 ( .a(FE_OFN908_n_4734), .o(g64178_sb) );
na03f02 TIMEBOOST_cell_66595 ( .a(TIMEBOOST_net_16786), .b(FE_OFN1315_n_6624), .c(g62635_sb), .o(n_6281) );
na02f02 TIMEBOOST_cell_53868 ( .a(TIMEBOOST_net_17151), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_15502) );
na02m08 TIMEBOOST_cell_52877 ( .a(wbs_dat_i_22_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q), .o(TIMEBOOST_net_16656) );
in01m02 g64179_u0 ( .a(FE_OFN1049_n_16657), .o(g64179_sb) );
na02s02 TIMEBOOST_cell_52474 ( .a(TIMEBOOST_net_16454), .b(g58156_sb), .o(TIMEBOOST_net_9558) );
in01s01 TIMEBOOST_cell_73988 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .o(TIMEBOOST_net_23553) );
na03m02 TIMEBOOST_cell_67411 ( .a(g58293_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q), .c(TIMEBOOST_net_10804), .o(TIMEBOOST_net_9394) );
in01f01 g64180_u0 ( .a(FE_OFN1011_n_4734), .o(g64180_sb) );
na02m10 TIMEBOOST_cell_45551 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q), .o(TIMEBOOST_net_13670) );
na03m02 TIMEBOOST_cell_65900 ( .a(n_4618), .b(g61837_sb), .c(g61837_db), .o(n_6973) );
in01m01 g64181_u0 ( .a(FE_OFN908_n_4734), .o(g64181_sb) );
na03s02 TIMEBOOST_cell_32083 ( .a(g58108_sb), .b(g58137_db), .c(FE_OFN254_n_9825), .o(n_9659) );
na02m04 TIMEBOOST_cell_53123 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_403), .b(FE_OFN2072_n_15978), .o(TIMEBOOST_net_16779) );
in01f01 g64182_u0 ( .a(FE_OFN1011_n_4734), .o(g64182_sb) );
na02m02 TIMEBOOST_cell_44231 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q), .b(g58371_sb), .o(TIMEBOOST_net_13010) );
na03f02 TIMEBOOST_cell_34834 ( .a(TIMEBOOST_net_9559), .b(FE_OFN1422_n_8567), .c(g57211_sb), .o(n_11545) );
na02f02 TIMEBOOST_cell_53310 ( .a(TIMEBOOST_net_16872), .b(FE_RN_715_0), .o(n_12148) );
in01m02 g64183_u0 ( .a(FE_OFN1049_n_16657), .o(g64183_sb) );
na02f01 TIMEBOOST_cell_37462 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(g65691_sb), .o(TIMEBOOST_net_10343) );
na02s01 TIMEBOOST_cell_37463 ( .a(TIMEBOOST_net_10343), .b(g65765_db), .o(n_1916) );
in01f01 g64184_u0 ( .a(FE_OFN1011_n_4734), .o(g64184_sb) );
na03m02 TIMEBOOST_cell_66479 ( .a(TIMEBOOST_net_10728), .b(g64957_sb), .c(n_40), .o(TIMEBOOST_net_20623) );
na02f01 g64184_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN1011_n_4734), .o(g64184_db) );
in01m01 g64185_u0 ( .a(FE_OFN908_n_4734), .o(g64185_sb) );
na02m02 TIMEBOOST_cell_63377 ( .a(TIMEBOOST_net_20635), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_15798) );
na02m06 TIMEBOOST_cell_68296 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q), .b(n_4677), .o(TIMEBOOST_net_21356) );
in01m02 g64186_u0 ( .a(FE_OFN1013_n_4734), .o(g64186_sb) );
na03s02 TIMEBOOST_cell_73677 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q), .b(g58229_db), .c(FE_OFN260_n_9860), .o(TIMEBOOST_net_20601) );
na02m01 TIMEBOOST_cell_62534 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_147), .o(TIMEBOOST_net_20214) );
in01m01 g64187_u0 ( .a(FE_OFN1051_n_16657), .o(g64187_sb) );
na02f02 TIMEBOOST_cell_50568 ( .a(TIMEBOOST_net_15501), .b(g62442_sb), .o(n_6712) );
na02m02 g64187_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q), .b(FE_OFN1051_n_16657), .o(g64187_db) );
in01s01 TIMEBOOST_cell_35487 ( .a(TIMEBOOST_net_10078), .o(TIMEBOOST_net_10077) );
in01m01 g64188_u0 ( .a(FE_OFN906_n_4736), .o(g64188_sb) );
na02m01 TIMEBOOST_cell_62984 ( .a(configuration_wb_err_addr_556), .b(conf_wb_err_addr_in_965), .o(TIMEBOOST_net_20439) );
na03f02 TIMEBOOST_cell_72680 ( .a(TIMEBOOST_net_16186), .b(FE_OFN786_n_2678), .c(g65211_sb), .o(n_2677) );
na02f01 TIMEBOOST_cell_49688 ( .a(TIMEBOOST_net_15061), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_13165) );
in01f01 g64189_u0 ( .a(FE_OFN905_n_4736), .o(g64189_sb) );
na02m04 TIMEBOOST_cell_42851 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_122), .o(TIMEBOOST_net_12320) );
na03m04 TIMEBOOST_cell_72847 ( .a(g65055_sb), .b(n_36), .c(TIMEBOOST_net_10641), .o(TIMEBOOST_net_17084) );
in01m01 g64190_u0 ( .a(FE_OFN1785_n_1699), .o(g64190_sb) );
na02s01 TIMEBOOST_cell_43425 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q), .o(TIMEBOOST_net_12607) );
na02m02 TIMEBOOST_cell_43423 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q), .b(g65315_sb), .o(TIMEBOOST_net_12606) );
in01m02 g64191_u0 ( .a(FE_OFN905_n_4736), .o(g64191_sb) );
na02s01 TIMEBOOST_cell_45409 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q), .o(TIMEBOOST_net_13599) );
na02f01 TIMEBOOST_cell_63053 ( .a(TIMEBOOST_net_20473), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_15558) );
in01m04 g64192_u0 ( .a(FE_OFN1051_n_16657), .o(g64192_sb) );
na03m01 TIMEBOOST_cell_41897 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q), .b(g58272_sb), .c(TIMEBOOST_net_9884), .o(n_9529) );
na03f02 TIMEBOOST_cell_66884 ( .a(FE_OFN1748_n_12004), .b(n_12010), .c(TIMEBOOST_net_13560), .o(n_12732) );
in01m02 g64193_u0 ( .a(FE_OFN1051_n_16657), .o(g64193_sb) );
na04f04 TIMEBOOST_cell_24778 ( .a(wbu_addr_in_271), .b(g52606_sb), .c(g52606_db), .d(TIMEBOOST_net_748), .o(n_11865) );
na03s02 TIMEBOOST_cell_41899 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q), .b(TIMEBOOST_net_9883), .c(g58342_sb), .o(n_9478) );
no02f01 g64194_u0 ( .a(n_1437), .b(pci_target_unit_wishbone_master_rty_counter_3_), .o(g64194_p) );
ao12f01 g64194_u1 ( .a(g64194_p), .b(pci_target_unit_wishbone_master_rty_counter_3_), .c(n_1437), .o(n_1662) );
in01m02 g64195_u0 ( .a(FE_OFN1051_n_16657), .o(g64195_sb) );
in01f04 TIMEBOOST_cell_35475 ( .a(TIMEBOOST_net_10066), .o(TIMEBOOST_net_10065) );
in01m02 g64196_u0 ( .a(FE_OFN903_n_4736), .o(g64196_sb) );
na02f01 TIMEBOOST_cell_44392 ( .a(TIMEBOOST_net_13090), .b(FE_OFN1115_g64577_p), .o(TIMEBOOST_net_11425) );
na02m10 TIMEBOOST_cell_41064 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q), .o(TIMEBOOST_net_12144) );
in01m01 g64197_u0 ( .a(FE_OFN906_n_4736), .o(g64197_sb) );
na03s01 TIMEBOOST_cell_72436 ( .a(pci_target_unit_del_sync_addr_in_230), .b(g66399_db), .c(g66399_sb), .o(n_2543) );
na03m02 TIMEBOOST_cell_73110 ( .a(TIMEBOOST_net_22075), .b(g65381_sb), .c(TIMEBOOST_net_22171), .o(TIMEBOOST_net_17060) );
in01f01 g64198_u0 ( .a(FE_OFN1011_n_4734), .o(g64198_sb) );
na03f02 TIMEBOOST_cell_44433 ( .a(TIMEBOOST_net_10318), .b(g60677_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q), .o(TIMEBOOST_net_13111) );
na03f02 TIMEBOOST_cell_73808 ( .a(TIMEBOOST_net_13782), .b(FE_OFN1775_n_13800), .c(FE_OFN1768_n_14054), .o(n_14508) );
na02f02 TIMEBOOST_cell_44434 ( .a(TIMEBOOST_net_13111), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_11408) );
in01m01 g64199_u0 ( .a(FE_OFN906_n_4736), .o(g64199_sb) );
na03f02 TIMEBOOST_cell_73521 ( .a(TIMEBOOST_net_13361), .b(n_6554), .c(g62434_sb), .o(n_6729) );
na02m01 g64199_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q), .b(FE_OFN906_n_4736), .o(g64199_db) );
in01s01 g64200_u0 ( .a(FE_OFN1051_n_16657), .o(g64200_sb) );
na03f02 TIMEBOOST_cell_73664 ( .a(TIMEBOOST_net_21062), .b(FE_OFN1135_g64577_p), .c(g62845_sb), .o(n_5281) );
na02m01 g64200_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q), .b(FE_OFN1051_n_16657), .o(g64200_db) );
na02s01 TIMEBOOST_cell_48875 ( .a(g57968_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q), .o(TIMEBOOST_net_14655) );
in01f02 g64201_u0 ( .a(FE_OFN906_n_4736), .o(g64201_sb) );
in01m01 g64202_u0 ( .a(FE_OFN905_n_4736), .o(g64202_sb) );
na02s02 TIMEBOOST_cell_39734 ( .a(FE_OFN203_n_9228), .b(g57892_sb), .o(TIMEBOOST_net_11479) );
na03m02 TIMEBOOST_cell_66095 ( .a(pci_target_unit_wishbone_master_bc_register_reg_3__Q), .b(g52593_sb), .c(TIMEBOOST_net_5510), .o(n_14683) );
na03s02 TIMEBOOST_cell_72552 ( .a(TIMEBOOST_net_13911), .b(g65679_sb), .c(g65679_db), .o(n_1956) );
in01m01 g64203_u0 ( .a(FE_OFN906_n_4736), .o(g64203_sb) );
na02m10 TIMEBOOST_cell_52663 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q), .o(TIMEBOOST_net_16549) );
na03f02 TIMEBOOST_cell_67582 ( .a(TIMEBOOST_net_13073), .b(FE_OFN1128_g64577_p), .c(g62756_sb), .o(n_6125) );
in01s01 g64204_u0 ( .a(FE_OFN1051_n_16657), .o(g64204_sb) );
na02s02 TIMEBOOST_cell_48119 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q), .b(FE_OFN1785_n_1699), .o(TIMEBOOST_net_14277) );
na02f01 TIMEBOOST_cell_49696 ( .a(TIMEBOOST_net_15065), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_13171) );
na04f04 TIMEBOOST_cell_24781 ( .a(n_10554), .b(n_9968), .c(n_10556), .d(n_9971), .o(n_12132) );
in01f01 g64205_u0 ( .a(FE_OFN1075_n_4740), .o(g64205_sb) );
in01m01 g64206_u0 ( .a(FE_OFN1049_n_16657), .o(g64206_sb) );
na02m01 TIMEBOOST_cell_54185 ( .a(conf_wb_err_addr_in_952), .b(configuration_wb_err_addr_543), .o(TIMEBOOST_net_17310) );
na02f01 g64206_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q), .b(FE_OFN1049_n_16657), .o(g64206_db) );
na02s01 TIMEBOOST_cell_62428 ( .a(g58779_sb), .b(FE_OFN2054_n_8831), .o(TIMEBOOST_net_20161) );
in01m02 g64207_u0 ( .a(FE_OFN905_n_4736), .o(g64207_sb) );
na02s01 TIMEBOOST_cell_39736 ( .a(FE_OFN201_n_9230), .b(g57894_sb), .o(TIMEBOOST_net_11480) );
na03f02 TIMEBOOST_cell_34849 ( .a(TIMEBOOST_net_9370), .b(FE_OFN1398_n_8567), .c(g58597_sb), .o(n_9189) );
na02s01 TIMEBOOST_cell_42775 ( .a(n_1218), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(TIMEBOOST_net_12282) );
in01m02 g64208_u0 ( .a(FE_OFN1049_n_16657), .o(g64208_sb) );
na03f02 TIMEBOOST_cell_73731 ( .a(TIMEBOOST_net_8603), .b(FE_OFN1572_n_11027), .c(n_12362), .o(n_12788) );
na02m08 TIMEBOOST_cell_45473 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q), .o(TIMEBOOST_net_13631) );
na02m08 TIMEBOOST_cell_37336 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q), .o(TIMEBOOST_net_10280) );
in01f02 g64209_u0 ( .a(FE_OFN1075_n_4740), .o(g64209_sb) );
na04f04 TIMEBOOST_cell_25168 ( .a(n_12341), .b(n_12195), .c(n_12196), .d(n_12112), .o(n_12868) );
na02f02 TIMEBOOST_cell_68291 ( .a(TIMEBOOST_net_21353), .b(n_969), .o(TIMEBOOST_net_20668) );
in01m02 g64210_u0 ( .a(FE_OFN1051_n_16657), .o(g64210_sb) );
na04f04 TIMEBOOST_cell_24782 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q), .b(g58820_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q), .d(FE_OFN2158_n_16439), .o(n_8621) );
na04f04 TIMEBOOST_cell_24783 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q), .b(g58819_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q), .d(FE_OFN2158_n_16439), .o(n_8622) );
in01m04 g64211_u0 ( .a(FE_OFN1077_n_4740), .o(g64211_sb) );
na02s02 TIMEBOOST_cell_48830 ( .a(TIMEBOOST_net_14632), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_10843) );
na03m02 TIMEBOOST_cell_68007 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_31__Q), .b(FE_OFN1082_n_13221), .c(FE_OFN1001_n_15978), .o(TIMEBOOST_net_655) );
in01m04 g64212_u0 ( .a(FE_OFN923_n_4740), .o(g64212_sb) );
in01m02 g64213_u0 ( .a(FE_OFN1051_n_16657), .o(g64213_sb) );
na02m02 TIMEBOOST_cell_69101 ( .a(TIMEBOOST_net_21758), .b(TIMEBOOST_net_20236), .o(TIMEBOOST_net_17465) );
na02f01 TIMEBOOST_cell_72254 ( .a(TIMEBOOST_net_16733), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_23335) );
in01m06 g64214_u0 ( .a(FE_OFN1076_n_4740), .o(g64214_sb) );
na02f02 TIMEBOOST_cell_70763 ( .a(TIMEBOOST_net_22589), .b(g52403_sb), .o(TIMEBOOST_net_684) );
na02s01 TIMEBOOST_cell_38777 ( .a(TIMEBOOST_net_11000), .b(g65813_sb), .o(n_2595) );
in01m06 g64215_u0 ( .a(FE_OFN1050_n_16657), .o(g64215_sb) );
na03f02 TIMEBOOST_cell_68009 ( .a(TIMEBOOST_net_17470), .b(FE_OFN1260_n_4143), .c(g62398_sb), .o(n_6804) );
na02f01 TIMEBOOST_cell_71074 ( .a(TIMEBOOST_net_17404), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_22745) );
na02s01 TIMEBOOST_cell_48172 ( .a(TIMEBOOST_net_14303), .b(g58172_sb), .o(TIMEBOOST_net_12480) );
in01m02 g64216_u0 ( .a(FE_OFN905_n_4736), .o(g64216_sb) );
na04f02 TIMEBOOST_cell_33560 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q), .b(FE_OCPN1909_n_16497), .c(pci_target_unit_pcit_if_pcir_fifo_data_in_768), .d(g54322_sb), .o(n_12998) );
na02s02 TIMEBOOST_cell_62955 ( .a(TIMEBOOST_net_20424), .b(g58117_sb), .o(TIMEBOOST_net_9407) );
na04f02 TIMEBOOST_cell_33561 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q), .b(FE_OCPN1909_n_16497), .c(pci_target_unit_pcit_if_pcir_fifo_data_in_770), .d(g54324_sb), .o(n_12994) );
in01m01 g64217_u0 ( .a(FE_OFN1051_n_16657), .o(g64217_sb) );
na04f04 TIMEBOOST_cell_24784 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q), .b(g58818_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q), .d(FE_OFN2157_n_16439), .o(n_8623) );
na04f04 TIMEBOOST_cell_24785 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q), .b(g58817_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q), .d(FE_OFN2156_n_16439), .o(n_8624) );
in01m01 g64218_u0 ( .a(FE_OFN1077_n_4740), .o(g64218_sb) );
na03f02 TIMEBOOST_cell_73412 ( .a(TIMEBOOST_net_17365), .b(FE_OFN1248_n_4093), .c(g62525_sb), .o(n_6526) );
na02m02 TIMEBOOST_cell_71921 ( .a(TIMEBOOST_net_23168), .b(g64849_db), .o(TIMEBOOST_net_17415) );
na02f02 TIMEBOOST_cell_52920 ( .a(TIMEBOOST_net_16677), .b(g63554_sb), .o(n_4603) );
in01m02 g64219_u0 ( .a(FE_OFN903_n_4736), .o(g64219_sb) );
na02m04 TIMEBOOST_cell_68702 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q), .b(FE_OFN687_n_4417), .o(TIMEBOOST_net_21559) );
na02m04 TIMEBOOST_cell_69906 ( .a(g65000_sb), .b(n_27), .o(TIMEBOOST_net_22161) );
na03s08 TIMEBOOST_cell_72423 ( .a(FE_OFN2054_n_8831), .b(n_8832), .c(wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q), .o(n_9230) );
in01f01 g64220_u0 ( .a(FE_OFN1076_n_4740), .o(g64220_sb) );
in01s01 TIMEBOOST_cell_45956 ( .a(TIMEBOOST_net_13917), .o(TIMEBOOST_net_13916) );
in01m01 g64221_u0 ( .a(FE_OFN1076_n_4740), .o(g64221_sb) );
na02f01 TIMEBOOST_cell_52834 ( .a(TIMEBOOST_net_16634), .b(FE_OFN1075_n_4740), .o(TIMEBOOST_net_14887) );
na02f02 TIMEBOOST_cell_71923 ( .a(TIMEBOOST_net_23169), .b(g64353_sb), .o(TIMEBOOST_net_13106) );
na03f02 TIMEBOOST_cell_66917 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_16495), .c(FE_OFN1513_n_14987), .o(n_12738) );
in01m02 g64222_u0 ( .a(FE_OFN1074_n_4740), .o(g64222_sb) );
na02s01 TIMEBOOST_cell_68176 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_408), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q), .o(TIMEBOOST_net_21296) );
na02m02 TIMEBOOST_cell_71925 ( .a(TIMEBOOST_net_23170), .b(TIMEBOOST_net_14213), .o(TIMEBOOST_net_17360) );
in01m01 g64223_u0 ( .a(FE_OFN1051_n_16657), .o(g64223_sb) );
na04f04 TIMEBOOST_cell_24786 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q), .b(g58816_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q), .d(FE_OFN2158_n_16439), .o(n_8625) );
na02m02 TIMEBOOST_cell_71434 ( .a(FE_OFN1186_n_3476), .b(configuration_pci_err_cs_bit9), .o(TIMEBOOST_net_22925) );
na04f04 TIMEBOOST_cell_24787 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q), .b(g58815_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q), .d(FE_OFN2153_n_16439), .o(n_8626) );
in01s01 g64224_u0 ( .a(FE_OFN1016_n_2053), .o(g64224_sb) );
na02f02 TIMEBOOST_cell_50614 ( .a(TIMEBOOST_net_15524), .b(g62993_sb), .o(n_5896) );
na03f02 TIMEBOOST_cell_66697 ( .a(TIMEBOOST_net_17123), .b(FE_OFN1316_n_6624), .c(g62902_sb), .o(n_6073) );
na02f01 TIMEBOOST_cell_43947 ( .a(TIMEBOOST_net_7109), .b(FE_OFN1031_n_4732), .o(TIMEBOOST_net_12868) );
in01s01 g64225_u0 ( .a(FE_OFN2111_n_2248), .o(g64225_sb) );
na02m01 TIMEBOOST_cell_71885 ( .a(TIMEBOOST_net_23150), .b(FE_OFN686_n_4417), .o(TIMEBOOST_net_10506) );
na02m02 TIMEBOOST_cell_68197 ( .a(TIMEBOOST_net_21306), .b(g65835_sb), .o(n_2185) );
in01s01 g64226_u0 ( .a(FE_OFN1042_n_2037), .o(g64226_sb) );
na04f04 TIMEBOOST_cell_24296 ( .a(n_9623), .b(g57307_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q), .d(FE_OFN1425_n_8567), .o(n_11443) );
na03f02 TIMEBOOST_cell_73635 ( .a(TIMEBOOST_net_17366), .b(FE_OFN1246_n_4093), .c(g62361_sb), .o(n_6876) );
in01s01 g64227_u0 ( .a(FE_OFN918_n_4725), .o(g64227_sb) );
na03f02 TIMEBOOST_cell_66288 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q), .b(g62326_sb), .c(g62326_db), .o(n_6937) );
in01s01 TIMEBOOST_cell_67721 ( .a(pci_target_unit_fifos_pcir_data_in_166), .o(TIMEBOOST_net_21148) );
in01s01 TIMEBOOST_cell_67780 ( .a(TIMEBOOST_net_21207), .o(TIMEBOOST_net_21206) );
in01m01 g64228_u0 ( .a(FE_OFN912_n_4727), .o(g64228_sb) );
na02m01 TIMEBOOST_cell_29545 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_404), .b(FE_OFN1000_n_15978), .o(TIMEBOOST_net_8877) );
na03m04 TIMEBOOST_cell_68400 ( .a(FE_OFN1001_n_15978), .b(conf_wb_err_bc_in_846), .c(wishbone_slave_unit_del_sync_bc_out_reg_1__Q), .o(TIMEBOOST_net_21408) );
in01m01 g64229_u0 ( .a(FE_OFN1056_n_4727), .o(g64229_sb) );
na04m04 TIMEBOOST_cell_67506 ( .a(n_1876), .b(FE_OFN704_n_8069), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q), .d(g61916_sb), .o(n_7989) );
na02s01 TIMEBOOST_cell_37601 ( .a(TIMEBOOST_net_10412), .b(g58046_db), .o(n_9744) );
in01m02 g64230_u0 ( .a(FE_OFN1056_n_4727), .o(g64230_sb) );
no02f02 TIMEBOOST_cell_51521 ( .a(TIMEBOOST_net_7529), .b(FE_RN_377_0), .o(TIMEBOOST_net_15978) );
in01m02 g64231_u0 ( .a(FE_OFN1035_n_4732), .o(g64231_sb) );
na02f08 TIMEBOOST_cell_42726 ( .a(TIMEBOOST_net_12257), .b(n_1409), .o(n_1410) );
na02s02 TIMEBOOST_cell_49450 ( .a(TIMEBOOST_net_14942), .b(g58237_sb), .o(n_9554) );
na02m10 TIMEBOOST_cell_51673 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q), .o(TIMEBOOST_net_16054) );
in01f01 g64232_u0 ( .a(FE_OFN1055_n_4727), .o(g64232_sb) );
in01s01 TIMEBOOST_cell_73830 ( .a(n_1545), .o(TIMEBOOST_net_23395) );
in01f01 g64233_u0 ( .a(FE_OFN1055_n_4727), .o(g64233_sb) );
na02m01 TIMEBOOST_cell_62450 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q), .o(TIMEBOOST_net_20172) );
na02m01 TIMEBOOST_cell_62816 ( .a(n_4645), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q), .o(TIMEBOOST_net_20355) );
na03m06 TIMEBOOST_cell_64762 ( .a(n_3749), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q), .c(FE_OFN1663_n_4490), .o(TIMEBOOST_net_16243) );
in01m01 g64234_u0 ( .a(FE_OFN1056_n_4727), .o(g64234_sb) );
na02s01 TIMEBOOST_cell_37586 ( .a(g58023_sb), .b(FE_OFN227_n_9841), .o(TIMEBOOST_net_10405) );
na02m01 TIMEBOOST_cell_49386 ( .a(TIMEBOOST_net_14910), .b(TIMEBOOST_net_569), .o(n_2577) );
in01m01 g64235_u0 ( .a(FE_OFN1034_n_4732), .o(g64235_sb) );
na03f02 TIMEBOOST_cell_34872 ( .a(TIMEBOOST_net_9394), .b(FE_OFN1368_n_8567), .c(g57430_sb), .o(n_10359) );
na03f02 TIMEBOOST_cell_73327 ( .a(TIMEBOOST_net_13112), .b(FE_OFN1135_g64577_p), .c(g62770_sb), .o(n_5454) );
na02s01 TIMEBOOST_cell_70118 ( .a(TIMEBOOST_net_12775), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q), .o(TIMEBOOST_net_22267) );
in01m01 g64236_u0 ( .a(FE_OFN1033_n_4732), .o(g64236_sb) );
na03s02 TIMEBOOST_cell_41618 ( .a(g58077_sb), .b(FE_OFN219_n_9853), .c(g58077_db), .o(n_9717) );
in01f01 g64237_u0 ( .a(FE_OFN1055_n_4727), .o(g64237_sb) );
na02f01 g64237_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(FE_OFN1055_n_4727), .o(g64237_db) );
in01f01 g64238_u0 ( .a(FE_OFN1056_n_4727), .o(g64238_sb) );
na03m02 TIMEBOOST_cell_72684 ( .a(TIMEBOOST_net_21454), .b(TIMEBOOST_net_16183), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q), .o(TIMEBOOST_net_16782) );
na02s02 TIMEBOOST_cell_48178 ( .a(TIMEBOOST_net_14306), .b(FE_OFN2109_n_2047), .o(TIMEBOOST_net_12696) );
in01m02 g64239_u0 ( .a(FE_OFN1032_n_4732), .o(g64239_sb) );
na04f04 TIMEBOOST_cell_24822 ( .a(n_10048), .b(n_9265), .c(n_16834), .d(n_16835), .o(n_12145) );
na04f02 TIMEBOOST_cell_24823 ( .a(n_10627), .b(n_10922), .c(n_10630), .d(n_12573), .o(n_12835) );
in01m01 g64240_u0 ( .a(FE_OFN1055_n_4727), .o(g64240_sb) );
na04f04 TIMEBOOST_cell_73328 ( .a(n_3925), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q), .c(FE_OFN1140_g64577_p), .d(g63104_sb), .o(n_5046) );
na02s01 TIMEBOOST_cell_48180 ( .a(TIMEBOOST_net_14307), .b(FE_OFN2108_n_2047), .o(TIMEBOOST_net_12699) );
in01m01 g64241_u0 ( .a(FE_OFN917_n_4725), .o(g64241_sb) );
na02s01 TIMEBOOST_cell_53059 ( .a(wbm_adr_o_2_), .b(configuration_pci_err_addr_472), .o(TIMEBOOST_net_16747) );
na03m02 TIMEBOOST_cell_69138 ( .a(n_3744), .b(g64963_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q), .o(TIMEBOOST_net_21777) );
na02m02 TIMEBOOST_cell_72333 ( .a(TIMEBOOST_net_23374), .b(g58281_sb), .o(TIMEBOOST_net_9340) );
in01m06 g64242_u0 ( .a(FE_OFN1056_n_4727), .o(g64242_sb) );
na02m10 TIMEBOOST_cell_51675 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q), .o(TIMEBOOST_net_16055) );
na02m02 g64242_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(FE_OFN1056_n_4727), .o(g64242_db) );
in01m04 g64243_u0 ( .a(FE_OFN1056_n_4727), .o(g64243_sb) );
na02f01 TIMEBOOST_cell_69922 ( .a(TIMEBOOST_net_12866), .b(n_16791), .o(TIMEBOOST_net_22169) );
na02m01 TIMEBOOST_cell_48184 ( .a(TIMEBOOST_net_14309), .b(FE_OFN2109_n_2047), .o(TIMEBOOST_net_12697) );
in01f01 g64244_u0 ( .a(FE_OFN1055_n_4727), .o(g64244_sb) );
na02f02 TIMEBOOST_cell_72315 ( .a(TIMEBOOST_net_23365), .b(g54170_sb), .o(n_13500) );
na02f01 g64244_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_143), .b(FE_OFN1055_n_4727), .o(g64244_db) );
na03m02 TIMEBOOST_cell_67164 ( .a(n_3792), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q), .c(FE_OFN687_n_4417), .o(TIMEBOOST_net_10455) );
in01m01 g64245_u0 ( .a(FE_OFN1057_n_4727), .o(g64245_sb) );
na02s01 TIMEBOOST_cell_70492 ( .a(TIMEBOOST_net_20449), .b(FE_OFN525_n_9899), .o(TIMEBOOST_net_22454) );
na03s03 TIMEBOOST_cell_64471 ( .a(TIMEBOOST_net_21177), .b(g65803_sb), .c(TIMEBOOST_net_14159), .o(n_2187) );
na02s02 TIMEBOOST_cell_53873 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q), .b(g58343_sb), .o(TIMEBOOST_net_17154) );
in01m02 g64246_u0 ( .a(FE_OFN1055_n_4727), .o(g64246_sb) );
na03f02 TIMEBOOST_cell_42039 ( .a(TIMEBOOST_net_5269), .b(g62114_sb), .c(g62114_db), .o(n_5582) );
na03f02 TIMEBOOST_cell_66864 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_16478), .c(FE_OFN1584_n_12306), .o(n_12485) );
in01m02 g64247_u0 ( .a(FE_OFN1032_n_4732), .o(g64247_sb) );
na04f04 TIMEBOOST_cell_24824 ( .a(g55853_sb), .b(pci_target_unit_pci_target_sm_n_3), .c(n_9177), .d(n_9175), .o(n_9176) );
in01s01 TIMEBOOST_cell_73897 ( .a(TIMEBOOST_net_23461), .o(TIMEBOOST_net_23462) );
na04f04 TIMEBOOST_cell_24825 ( .a(g55852_sb), .b(pci_target_unit_pci_target_sm_n_2), .c(n_9177), .d(n_9178), .o(n_9179) );
in01m01 g64248_u0 ( .a(FE_OFN1056_n_4727), .o(g64248_sb) );
in01s01 TIMEBOOST_cell_67783 ( .a(TIMEBOOST_net_21221), .o(TIMEBOOST_net_21210) );
oa12m02 g64249_u0 ( .a(n_3805), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_2__231), .c(FE_OFN1036_n_4732), .o(n_4733) );
in01m06 g64250_u0 ( .a(FE_OFN912_n_4727), .o(g64250_sb) );
na03f10 TIMEBOOST_cell_31948 ( .a(n_696), .b(n_15331), .c(n_16936), .o(n_2687) );
na02m04 g64250_u2 ( .a(FE_OFN912_n_4727), .b(pci_target_unit_fifos_pciw_addr_data_in_148), .o(g64250_db) );
na02f02 TIMEBOOST_cell_51835 ( .a(FE_OFN1589_n_13736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q), .o(TIMEBOOST_net_16135) );
in01m02 g64251_u0 ( .a(FE_OFN1057_n_4727), .o(g64251_sb) );
na03f02 TIMEBOOST_cell_72617 ( .a(TIMEBOOST_net_16899), .b(FE_OFN908_n_4734), .c(g64162_sb), .o(TIMEBOOST_net_13047) );
na03m02 TIMEBOOST_cell_70360 ( .a(FE_OFN2022_n_4778), .b(TIMEBOOST_net_16655), .c(TIMEBOOST_net_635), .o(TIMEBOOST_net_22388) );
in01m01 g64252_u0 ( .a(FE_OFN912_n_4727), .o(g64252_sb) );
na02m01 g64252_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(FE_OFN912_n_4727), .o(g64252_db) );
na03m02 TIMEBOOST_cell_72862 ( .a(TIMEBOOST_net_21712), .b(g65414_sb), .c(TIMEBOOST_net_21944), .o(TIMEBOOST_net_17018) );
in01f01 g64253_u0 ( .a(FE_OFN1033_n_4732), .o(g64253_sb) );
na02m02 TIMEBOOST_cell_48186 ( .a(TIMEBOOST_net_14310), .b(FE_OFN1797_n_2299), .o(TIMEBOOST_net_12695) );
na03f02 TIMEBOOST_cell_32958 ( .a(TIMEBOOST_net_8278), .b(n_5633), .c(g62072_sb), .o(n_5639) );
na02m01 TIMEBOOST_cell_48393 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q), .b(FE_OFN654_n_4508), .o(TIMEBOOST_net_14414) );
in01m01 g64254_u0 ( .a(FE_OFN918_n_4725), .o(g64254_sb) );
na03s02 TIMEBOOST_cell_72522 ( .a(TIMEBOOST_net_14155), .b(g65756_sb), .c(g65756_db), .o(TIMEBOOST_net_7113) );
na03f08 TIMEBOOST_cell_67846 ( .a(n_1966), .b(n_1965), .c(n_2914), .o(TIMEBOOST_net_20827) );
na02s01 TIMEBOOST_cell_52445 ( .a(configuration_pci_err_addr_491), .b(wbm_adr_o_21_), .o(TIMEBOOST_net_16440) );
in01m01 g64255_u0 ( .a(FE_OFN912_n_4727), .o(g64255_sb) );
na02s02 TIMEBOOST_cell_53874 ( .a(TIMEBOOST_net_17154), .b(TIMEBOOST_net_12949), .o(TIMEBOOST_net_10009) );
na03f02 TIMEBOOST_cell_73522 ( .a(TIMEBOOST_net_13360), .b(n_6431), .c(g62588_sb), .o(n_6374) );
na04f04 TIMEBOOST_cell_24715 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_21__Q), .b(g58468_sb), .c(FE_OFN223_n_9844), .d(FE_OFN1441_n_9372), .o(n_9379) );
in01m01 g64256_u0 ( .a(FE_OFN912_n_4727), .o(g64256_sb) );
in01m01 g64257_u0 ( .a(FE_OFN1057_n_4727), .o(g64257_sb) );
na02m10 TIMEBOOST_cell_52667 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q), .o(TIMEBOOST_net_16551) );
na02f02 TIMEBOOST_cell_71747 ( .a(TIMEBOOST_net_23081), .b(FE_OCP_RBN1962_FE_OFN1591_n_13741), .o(n_14268) );
na02f02 TIMEBOOST_cell_51694 ( .a(TIMEBOOST_net_16064), .b(n_12115), .o(n_12898) );
in01m01 g64258_u0 ( .a(FE_OFN1032_n_4732), .o(g64258_sb) );
na04f04 TIMEBOOST_cell_24826 ( .a(g55851_sb), .b(n_1628), .c(n_9177), .d(n_1384), .o(n_9180) );
na02f10 TIMEBOOST_cell_68204 ( .a(n_8831), .b(g58788_sb), .o(TIMEBOOST_net_21310) );
na04f02 TIMEBOOST_cell_24827 ( .a(n_10991), .b(n_10216), .c(n_10221), .d(n_12589), .o(n_12851) );
in01m08 g64259_u0 ( .a(FE_OFN1057_n_4727), .o(g64259_sb) );
na02f02 TIMEBOOST_cell_71393 ( .a(TIMEBOOST_net_22904), .b(g59112_sb), .o(n_8705) );
in01f01 g64260_u0 ( .a(FE_OFN1055_n_4727), .o(g64260_sb) );
na02s01 TIMEBOOST_cell_39740 ( .a(g57897_sb), .b(FE_OFN201_n_9230), .o(TIMEBOOST_net_11482) );
na03m02 TIMEBOOST_cell_72654 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(FE_OFN929_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q), .o(TIMEBOOST_net_23235) );
in01s01 g64261_u0 ( .a(FE_OFN1057_n_4727), .o(g64261_sb) );
na02m02 TIMEBOOST_cell_68827 ( .a(TIMEBOOST_net_21621), .b(n_4488), .o(TIMEBOOST_net_13239) );
na02s01 g64261_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(FE_OFN1057_n_4727), .o(g64261_db) );
na03f02 TIMEBOOST_cell_73636 ( .a(TIMEBOOST_net_13243), .b(FE_OFN1270_n_4095), .c(g62671_sb), .o(n_6196) );
in01m02 g64262_u0 ( .a(FE_OFN1058_n_4727), .o(g64262_sb) );
na03f02 TIMEBOOST_cell_72828 ( .a(g64171_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q), .c(TIMEBOOST_net_12613), .o(TIMEBOOST_net_15726) );
na02m03 TIMEBOOST_cell_48026 ( .a(TIMEBOOST_net_14230), .b(FE_OFN1013_n_4734), .o(TIMEBOOST_net_12541) );
in01m01 g64263_u0 ( .a(FE_OFN1055_n_4727), .o(g64263_sb) );
na02s01 TIMEBOOST_cell_45459 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q), .o(TIMEBOOST_net_13624) );
na02f02 TIMEBOOST_cell_72245 ( .a(TIMEBOOST_net_23330), .b(g63034_sb), .o(n_5179) );
in01m01 g64264_u0 ( .a(FE_OFN912_n_4727), .o(g64264_sb) );
in01m01 g64265_u0 ( .a(FE_OFN1055_n_4727), .o(g64265_sb) );
na03f02 TIMEBOOST_cell_67008 ( .a(FE_OFN1589_n_13736), .b(TIMEBOOST_net_16520), .c(FE_OCP_RBN1997_n_13971), .o(g53174_p) );
in01m01 g64266_u0 ( .a(FE_OFN1037_n_4732), .o(g64266_sb) );
in01m02 g64267_u0 ( .a(FE_OFN1036_n_4732), .o(g64267_sb) );
na03m02 TIMEBOOST_cell_72769 ( .a(n_4476), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q), .c(TIMEBOOST_net_12545), .o(TIMEBOOST_net_20615) );
in01m01 g64268_u0 ( .a(FE_OFN928_n_4730), .o(g64268_sb) );
in01s01 g64269_u0 ( .a(FE_OFN928_n_4730), .o(g64269_sb) );
in01m02 g64270_u0 ( .a(FE_OFN928_n_4730), .o(g64270_sb) );
na02f10 TIMEBOOST_cell_43949 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_779), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q), .o(TIMEBOOST_net_12869) );
na03f02 TIMEBOOST_cell_34840 ( .a(TIMEBOOST_net_9390), .b(FE_OFN1387_n_8567), .c(g57577_sb), .o(n_11174) );
na03f02 TIMEBOOST_cell_65879 ( .a(FE_OFN720_n_8060), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q), .c(n_1873), .o(TIMEBOOST_net_15054) );
in01m01 g64271_u0 ( .a(FE_OFN928_n_4730), .o(g64271_sb) );
na03f02 TIMEBOOST_cell_72671 ( .a(TIMEBOOST_net_16583), .b(FE_OFN784_n_2678), .c(g65233_sb), .o(n_2654) );
in01m02 g64272_u0 ( .a(FE_OFN1032_n_4732), .o(g64272_sb) );
na04f02 TIMEBOOST_cell_24828 ( .a(n_10672), .b(n_10096), .c(n_10675), .d(n_12577), .o(n_12839) );
na03m02 TIMEBOOST_cell_72692 ( .a(TIMEBOOST_net_23160), .b(g65028_sb), .c(TIMEBOOST_net_21784), .o(TIMEBOOST_net_17097) );
in01m10 g64273_u0 ( .a(FE_OFN928_n_4730), .o(g64273_sb) );
na02f02 TIMEBOOST_cell_70808 ( .a(TIMEBOOST_net_16700), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_22612) );
na02m06 g64273_u2 ( .a(FE_OFN928_n_4730), .b(pci_target_unit_fifos_pciw_addr_data_in_134), .o(g64273_db) );
in01m01 g64274_u0 ( .a(FE_OFN928_n_4730), .o(g64274_sb) );
na02f01 TIMEBOOST_cell_44268 ( .a(TIMEBOOST_net_13028), .b(FE_OFN1095_g64577_p), .o(n_6951) );
in01m02 g64275_u0 ( .a(FE_OFN928_n_4730), .o(g64275_sb) );
na03f02 TIMEBOOST_cell_72389 ( .a(n_378), .b(TIMEBOOST_net_13), .c(n_2494), .o(TIMEBOOST_net_118) );
na03f02 TIMEBOOST_cell_34842 ( .a(TIMEBOOST_net_9336), .b(FE_OFN1411_n_8567), .c(g57104_sb), .o(n_11641) );
na02m02 TIMEBOOST_cell_63770 ( .a(TIMEBOOST_net_12693), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q), .o(TIMEBOOST_net_20871) );
in01s01 g64276_u0 ( .a(FE_OFN928_n_4730), .o(g64276_sb) );
na02f10 TIMEBOOST_cell_43951 ( .a(pci_target_unit_pcit_if_pcir_fifo_data_in_774), .b(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q), .o(TIMEBOOST_net_12870) );
na02m01 g64276_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(FE_OFN928_n_4730), .o(g64276_db) );
in01m02 g64277_u0 ( .a(FE_OFN930_n_4730), .o(g64277_sb) );
na02m02 g64277_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q), .b(g64277_sb), .o(g64277_da) );
na02m04 g64277_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(FE_OFN930_n_4730), .o(g64277_db) );
in01m01 g64278_u0 ( .a(FE_OFN917_n_4725), .o(g64278_sb) );
na02s02 TIMEBOOST_cell_64090 ( .a(FE_OFN264_n_9849), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q), .o(TIMEBOOST_net_21031) );
in01m01 g64279_u0 ( .a(FE_OFN930_n_4730), .o(g64279_sb) );
na02s01 TIMEBOOST_cell_51839 ( .a(wbs_dat_i_17_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q), .o(TIMEBOOST_net_16137) );
na02s01 TIMEBOOST_cell_51840 ( .a(TIMEBOOST_net_16137), .b(g61943_sb), .o(TIMEBOOST_net_12832) );
in01m01 g64280_u0 ( .a(FE_OFN928_n_4730), .o(g64280_sb) );
na02f02 TIMEBOOST_cell_70807 ( .a(TIMEBOOST_net_22611), .b(g62042_sb), .o(n_7771) );
na02m01 g64280_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(FE_OFN928_n_4730), .o(g64280_db) );
na02s01 TIMEBOOST_cell_51841 ( .a(wbs_dat_i_23_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q), .o(TIMEBOOST_net_16138) );
in01m02 g64281_u0 ( .a(FE_OFN930_n_4730), .o(g64281_sb) );
na02s01 TIMEBOOST_cell_51842 ( .a(TIMEBOOST_net_16138), .b(g61943_sb), .o(TIMEBOOST_net_12833) );
na03f02 TIMEBOOST_cell_34844 ( .a(TIMEBOOST_net_9412), .b(FE_OFN1388_n_8567), .c(g57454_sb), .o(n_11280) );
na02f10 TIMEBOOST_cell_43953 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_771), .o(TIMEBOOST_net_12871) );
in01m01 g64282_u0 ( .a(FE_OFN928_n_4730), .o(g64282_sb) );
na03f02 TIMEBOOST_cell_66701 ( .a(TIMEBOOST_net_17119), .b(FE_OFN1314_n_6624), .c(g62523_sb), .o(n_6530) );
in01s01 g64283_u0 ( .a(FE_OFN1037_n_4732), .o(g64283_sb) );
na02m01 TIMEBOOST_cell_64130 ( .a(n_8272), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q), .o(TIMEBOOST_net_21051) );
na02m01 g64283_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(FE_OFN1037_n_4732), .o(g64283_db) );
na03f02 TIMEBOOST_cell_73464 ( .a(TIMEBOOST_net_17543), .b(FE_OFN1213_n_4151), .c(g62629_sb), .o(n_6297) );
in01m01 g64284_u0 ( .a(FE_OFN928_n_4730), .o(g64284_sb) );
na02m02 TIMEBOOST_cell_68956 ( .a(g64961_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q), .o(TIMEBOOST_net_21686) );
na02m02 TIMEBOOST_cell_68111 ( .a(TIMEBOOST_net_21263), .b(g54207_sb), .o(TIMEBOOST_net_14036) );
in01f01 g64285_u0 ( .a(FE_OFN930_n_4730), .o(g64285_sb) );
in01f02 g64286_u0 ( .a(FE_OFN927_n_4730), .o(g64286_sb) );
na02s01 TIMEBOOST_cell_51563 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q), .o(TIMEBOOST_net_15999) );
in01m01 g64287_u0 ( .a(FE_OFN928_n_4730), .o(g64287_sb) );
na02m01 TIMEBOOST_cell_54016 ( .a(TIMEBOOST_net_17225), .b(FE_OFN928_n_4730), .o(TIMEBOOST_net_14479) );
na03m02 TIMEBOOST_cell_72808 ( .a(n_4479), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q), .c(TIMEBOOST_net_12537), .o(TIMEBOOST_net_17517) );
in01m02 g64288_u0 ( .a(FE_OFN1031_n_4732), .o(g64288_sb) );
na03f02 TIMEBOOST_cell_34874 ( .a(TIMEBOOST_net_9396), .b(FE_OFN1421_n_8567), .c(g57069_sb), .o(n_11672) );
na02f02 g64288_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(FE_OFN1031_n_4732), .o(g64288_db) );
na02m02 TIMEBOOST_cell_53063 ( .a(n_6136), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(TIMEBOOST_net_16749) );
in01m01 g64289_u0 ( .a(FE_OFN927_n_4730), .o(g64289_sb) );
na02f02 TIMEBOOST_cell_71518 ( .a(n_12313), .b(TIMEBOOST_net_13535), .o(TIMEBOOST_net_22967) );
in01m02 g64290_u0 ( .a(FE_OFN927_n_4730), .o(g64290_sb) );
in01s01 TIMEBOOST_cell_73933 ( .a(TIMEBOOST_net_23497), .o(TIMEBOOST_net_23498) );
na03f02 TIMEBOOST_cell_66362 ( .a(g62945_sb), .b(FE_OFN1234_n_6391), .c(TIMEBOOST_net_17497), .o(n_5991) );
in01m01 g64291_u0 ( .a(FE_OFN929_n_4730), .o(g64291_sb) );
na02m02 TIMEBOOST_cell_72118 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q), .b(pci_target_unit_fifos_pciw_cbe_in_152), .o(TIMEBOOST_net_23267) );
in01m02 g64292_u0 ( .a(FE_OFN927_n_4730), .o(g64292_sb) );
in01m01 g64293_u0 ( .a(FE_OFN929_n_4730), .o(g64293_sb) );
na03f02 TIMEBOOST_cell_73637 ( .a(TIMEBOOST_net_20623), .b(FE_OFN1268_n_4095), .c(g62681_sb), .o(n_6177) );
in01m04 TIMEBOOST_cell_35479 ( .a(TIMEBOOST_net_10069), .o(TIMEBOOST_net_10070) );
na02s01 TIMEBOOST_cell_53875 ( .a(g58450_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q), .o(TIMEBOOST_net_17155) );
in01m02 g64295_u0 ( .a(FE_OFN927_n_4730), .o(g64295_sb) );
na02f02 TIMEBOOST_cell_49717 ( .a(n_3932), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q), .o(TIMEBOOST_net_15076) );
na02m01 TIMEBOOST_cell_68534 ( .a(n_3739), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q), .o(TIMEBOOST_net_21475) );
in01m01 g64296_u0 ( .a(FE_OFN917_n_4725), .o(g64296_sb) );
na03f04 TIMEBOOST_cell_71448 ( .a(n_3290), .b(pciu_bar0_in_372), .c(FE_RN_570_0), .o(TIMEBOOST_net_22932) );
na02m02 TIMEBOOST_cell_62462 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_132), .o(TIMEBOOST_net_20178) );
no02f03 TIMEBOOST_cell_42847 ( .a(TIMEBOOST_net_102), .b(n_2430), .o(TIMEBOOST_net_12318) );
in01m08 g64297_u0 ( .a(FE_OFN1034_n_4732), .o(g64297_sb) );
na03f02 TIMEBOOST_cell_64469 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q), .b(FE_OFN575_n_9902), .c(TIMEBOOST_net_20195), .o(TIMEBOOST_net_14938) );
na02m02 TIMEBOOST_cell_49212 ( .a(g65820_db), .b(TIMEBOOST_net_14823), .o(n_1896) );
na03m08 TIMEBOOST_cell_64300 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q), .b(n_504), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_409), .o(TIMEBOOST_net_16955) );
in01m04 g64298_u0 ( .a(FE_OFN929_n_4730), .o(g64298_sb) );
na02f01 TIMEBOOST_cell_68608 ( .a(TIMEBOOST_net_170), .b(n_2341), .o(TIMEBOOST_net_21512) );
oa12m01 g64299_u0 ( .a(n_3807), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_1__192), .c(n_4730), .o(n_4729) );
in01m02 g64300_u0 ( .a(FE_OFN1031_n_4732), .o(g64300_sb) );
na02s08 TIMEBOOST_cell_62808 ( .a(pci_target_unit_fifos_pcir_data_in_185), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_20351) );
na02m10 TIMEBOOST_cell_45233 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q), .o(TIMEBOOST_net_13511) );
in01m02 g64301_u0 ( .a(FE_OFN929_n_4730), .o(g64301_sb) );
na03f02 TIMEBOOST_cell_73413 ( .a(TIMEBOOST_net_17559), .b(FE_OFN1248_n_4093), .c(g62490_sb), .o(n_6605) );
na03f02 TIMEBOOST_cell_34846 ( .a(TIMEBOOST_net_9427), .b(FE_OFN1388_n_8567), .c(g57113_sb), .o(n_11633) );
na02f01 TIMEBOOST_cell_68846 ( .a(TIMEBOOST_net_10278), .b(g65325_sb), .o(TIMEBOOST_net_21631) );
in01m01 g64302_u0 ( .a(FE_OFN929_n_4730), .o(g64302_sb) );
na02f01 g64302_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_125), .b(FE_OFN929_n_4730), .o(g64302_db) );
na02m01 TIMEBOOST_cell_71841 ( .a(TIMEBOOST_net_23128), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_397), .o(TIMEBOOST_net_16792) );
na02s01 TIMEBOOST_cell_49990 ( .a(TIMEBOOST_net_15212), .b(g57904_db), .o(TIMEBOOST_net_10013) );
na02s02 TIMEBOOST_cell_48028 ( .a(TIMEBOOST_net_14231), .b(FE_OFN523_n_9428), .o(TIMEBOOST_net_10774) );
in01m01 g64304_u0 ( .a(FE_OFN928_n_4730), .o(g64304_sb) );
na04f02 TIMEBOOST_cell_67804 ( .a(g58789_sb), .b(n_8831), .c(wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q), .d(wbu_addr_in_251), .o(n_9118) );
na02s01 TIMEBOOST_cell_68614 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q), .o(TIMEBOOST_net_21515) );
in01s01 g64306_u0 ( .a(FE_OFN928_n_4730), .o(g64306_sb) );
in01s01 TIMEBOOST_cell_63610 ( .a(TIMEBOOST_net_20790), .o(TIMEBOOST_net_20737) );
na03s02 TIMEBOOST_cell_72861 ( .a(g58004_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q), .c(TIMEBOOST_net_12911), .o(TIMEBOOST_net_14640) );
in01m01 g64307_u0 ( .a(FE_OFN1033_n_4732), .o(g64307_sb) );
in01s01 TIMEBOOST_cell_45982 ( .a(TIMEBOOST_net_13942), .o(TIMEBOOST_net_13943) );
in01s01 TIMEBOOST_cell_45983 ( .a(conf_wb_err_bc_in_847), .o(TIMEBOOST_net_13944) );
in01m01 g64308_u0 ( .a(FE_OFN1037_n_4732), .o(g64308_sb) );
in01s01 TIMEBOOST_cell_63549 ( .a(TIMEBOOST_net_20728), .o(TIMEBOOST_net_20729) );
in01s01 TIMEBOOST_cell_73934 ( .a(wbm_dat_i_18_), .o(TIMEBOOST_net_23499) );
in01f01 g64309_u0 ( .a(FE_OFN1032_n_4732), .o(g64309_sb) );
na04f04 TIMEBOOST_cell_24830 ( .a(wbu_addr_in_262), .b(g52597_sb), .c(g52597_db), .d(TIMEBOOST_net_772), .o(n_11874) );
na02m02 TIMEBOOST_cell_54628 ( .a(TIMEBOOST_net_17531), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_15370) );
na04f02 TIMEBOOST_cell_24831 ( .a(n_10131), .b(n_10708), .c(n_10711), .d(n_12581), .o(n_12843) );
in01m02 g64310_u0 ( .a(FE_OFN1032_n_4732), .o(g64310_sb) );
na04f04 TIMEBOOST_cell_24832 ( .a(n_10002), .b(n_10007), .c(n_16840), .d(n_16841), .o(n_12140) );
na04f02 TIMEBOOST_cell_73111 ( .a(n_1981), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q), .c(FE_OFN716_n_8176), .d(g61794_sb), .o(n_8210) );
na04f04 TIMEBOOST_cell_24833 ( .a(n_9993), .b(n_16844), .c(n_16845), .d(n_10577), .o(n_12137) );
in01m01 g64311_u0 ( .a(FE_OFN1032_n_4732), .o(g64311_sb) );
na03f02 TIMEBOOST_cell_72868 ( .a(TIMEBOOST_net_21729), .b(g65433_sb), .c(TIMEBOOST_net_22116), .o(TIMEBOOST_net_17136) );
na02f02 TIMEBOOST_cell_40853 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_12038), .o(n_12735) );
in01m02 g64312_u0 ( .a(FE_OFN1037_n_4732), .o(g64312_sb) );
na02m02 g64312_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(FE_OFN1037_n_4732), .o(g64312_db) );
na02f02 TIMEBOOST_cell_40855 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_12039), .o(n_12686) );
in01m01 g64313_u0 ( .a(FE_OFN1037_n_4732), .o(g64313_sb) );
na02s01 TIMEBOOST_cell_49232 ( .a(TIMEBOOST_net_14833), .b(g52466_da), .o(TIMEBOOST_net_11893) );
na04f04 TIMEBOOST_cell_67702 ( .a(TIMEBOOST_net_16862), .b(FE_OFN2200_n_10256), .c(g52598_sb), .d(TIMEBOOST_net_708), .o(n_11872) );
in01m01 g64314_u0 ( .a(FE_OFN1034_n_4732), .o(g64314_sb) );
na02m01 TIMEBOOST_cell_69802 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q), .o(TIMEBOOST_net_22109) );
na02f02 TIMEBOOST_cell_40859 ( .a(FE_OFN1577_n_12028), .b(TIMEBOOST_net_12041), .o(n_12631) );
in01f01 g64315_u0 ( .a(FE_OFN959_n_2299), .o(g64315_sb) );
na03m02 TIMEBOOST_cell_72647 ( .a(TIMEBOOST_net_21489), .b(g64839_sb), .c(TIMEBOOST_net_21675), .o(TIMEBOOST_net_17377) );
na02m02 TIMEBOOST_cell_69276 ( .a(n_4444), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q), .o(TIMEBOOST_net_21846) );
in01m02 g64316_u0 ( .a(FE_OFN1033_n_4732), .o(g64316_sb) );
na03m02 TIMEBOOST_cell_68011 ( .a(TIMEBOOST_net_14941), .b(FE_OFN272_n_9828), .c(TIMEBOOST_net_15079), .o(TIMEBOOST_net_9515) );
in01f01 g64317_u0 ( .a(FE_OFN930_n_4730), .o(g64317_sb) );
na04m04 TIMEBOOST_cell_67509 ( .a(n_1870), .b(FE_OFN704_n_8069), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q), .d(g61915_sb), .o(n_7991) );
na03f02 TIMEBOOST_cell_66707 ( .a(TIMEBOOST_net_17051), .b(n_6319), .c(g62979_sb), .o(n_5924) );
na04f04 TIMEBOOST_cell_73112 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q), .b(FE_OFN706_n_8119), .c(n_1937), .d(g61787_sb), .o(n_8229) );
in01m10 g64318_u0 ( .a(FE_OFN1037_n_4732), .o(g64318_sb) );
na03f02 TIMEBOOST_cell_24834 ( .a(n_14895), .b(n_13488), .c(n_14833), .o(n_14897) );
na03f02 TIMEBOOST_cell_24835 ( .a(n_14895), .b(n_13487), .c(n_14832), .o(n_14894) );
in01m01 g64319_u0 ( .a(FE_OFN1034_n_4732), .o(g64319_sb) );
na02m04 TIMEBOOST_cell_69794 ( .a(g65040_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q), .o(TIMEBOOST_net_22105) );
na04f04 TIMEBOOST_cell_65980 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q), .b(FE_OCPN1909_n_16497), .c(pci_target_unit_pcit_if_pcir_fifo_data_in), .d(g54330_sb), .o(n_12986) );
in01m02 g64320_u0 ( .a(FE_OFN1031_n_4732), .o(g64320_sb) );
na02s01 TIMEBOOST_cell_63260 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q), .b(FE_OFN516_n_9697), .o(TIMEBOOST_net_20577) );
na02f02 TIMEBOOST_cell_52850 ( .a(TIMEBOOST_net_16642), .b(g61908_sb), .o(n_8005) );
in01f01 g64321_u0 ( .a(FE_OFN1033_n_4732), .o(g64321_sb) );
na02m02 TIMEBOOST_cell_44246 ( .a(TIMEBOOST_net_13017), .b(g63618_sb), .o(n_7141) );
na02m10 TIMEBOOST_cell_53023 ( .a(configuration_pci_err_data_520), .b(wbm_dat_o_19_), .o(TIMEBOOST_net_16729) );
in01m01 g64322_u0 ( .a(FE_OFN1034_n_4732), .o(g64322_sb) );
no02f06 TIMEBOOST_cell_68065 ( .a(TIMEBOOST_net_21240), .b(n_1291), .o(TIMEBOOST_net_46) );
na03s01 TIMEBOOST_cell_67845 ( .a(n_2507), .b(g66398_sb), .c(g66421_db), .o(n_2508) );
na02m02 TIMEBOOST_cell_64050 ( .a(TIMEBOOST_net_7590), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q), .o(TIMEBOOST_net_21011) );
in01m01 g64323_u0 ( .a(FE_OFN1034_n_4732), .o(g64323_sb) );
na02f02 TIMEBOOST_cell_50386 ( .a(TIMEBOOST_net_15410), .b(g63167_sb), .o(n_5804) );
na02m04 TIMEBOOST_cell_69588 ( .a(g64984_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q), .o(TIMEBOOST_net_22002) );
in01f01 g64324_u0 ( .a(FE_OFN1034_n_4732), .o(g64324_sb) );
na02s01 TIMEBOOST_cell_29097 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q), .b(FE_OFN2054_n_8831), .o(TIMEBOOST_net_8653) );
na03m02 TIMEBOOST_cell_72782 ( .a(n_4470), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q), .c(TIMEBOOST_net_10631), .o(TIMEBOOST_net_17389) );
in01m02 g64325_u0 ( .a(FE_OFN1031_n_4732), .o(g64325_sb) );
na02f01 TIMEBOOST_cell_29099 ( .a(n_8511), .b(g63590_sb), .o(TIMEBOOST_net_8654) );
in01m01 g64326_u0 ( .a(FE_OFN1035_n_4732), .o(g64326_sb) );
na03f01 TIMEBOOST_cell_72432 ( .a(TIMEBOOST_net_10174), .b(FE_OFN945_n_2248), .c(g65857_sb), .o(n_1581) );
na03s01 TIMEBOOST_cell_41626 ( .a(g57993_sb), .b(FE_OFN227_n_9841), .c(g57993_db), .o(n_9802) );
in01m02 g64327_u0 ( .a(FE_OFN916_n_4725), .o(g64327_sb) );
na03m04 TIMEBOOST_cell_72838 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q), .b(g65434_sb), .c(TIMEBOOST_net_23288), .o(TIMEBOOST_net_17031) );
na03m04 TIMEBOOST_cell_72616 ( .a(FE_OFN1013_n_4734), .b(TIMEBOOST_net_20255), .c(g64130_sb), .o(n_4032) );
in01s01 TIMEBOOST_cell_73938 ( .a(wbm_dat_i_1_), .o(TIMEBOOST_net_23503) );
in01s01 g64328_u0 ( .a(FE_OFN917_n_4725), .o(g64328_sb) );
na03m01 TIMEBOOST_cell_22747 ( .a(FE_OFN258_n_9862), .b(g58199_sb), .c(g58199_db), .o(n_9586) );
na02f01 g64328_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_133), .b(FE_OFN917_n_4725), .o(g64328_db) );
na03s02 TIMEBOOST_cell_22746 ( .a(FE_OFN260_n_9860), .b(g58200_sb), .c(g58200_db), .o(n_9585) );
in01m02 g64329_u0 ( .a(FE_OFN917_n_4725), .o(g64329_sb) );
na02f01 TIMEBOOST_cell_48002 ( .a(TIMEBOOST_net_14218), .b(FE_OFN636_n_4669), .o(TIMEBOOST_net_10618) );
in01s01 TIMEBOOST_cell_67785 ( .a(TIMEBOOST_net_21212), .o(wbs_adr_i_27_) );
na03s01 TIMEBOOST_cell_22748 ( .a(FE_OFN260_n_9860), .b(g58140_sb), .c(g58140_db), .o(n_9655) );
in01m01 g64330_u0 ( .a(FE_OFN917_n_4725), .o(g64330_sb) );
na02m01 TIMEBOOST_cell_71910 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q), .b(FE_OFN685_n_4417), .o(TIMEBOOST_net_23163) );
na02m01 g64330_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_136), .b(FE_OFN917_n_4725), .o(g64330_db) );
na02m20 TIMEBOOST_cell_53099 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_14__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_397), .o(TIMEBOOST_net_16767) );
in01m02 g64331_u0 ( .a(FE_OFN917_n_4725), .o(g64331_sb) );
na03f02 TIMEBOOST_cell_66922 ( .a(FE_OFN1553_n_12104), .b(TIMEBOOST_net_16493), .c(FE_OCP_RBN1980_n_10273), .o(n_16597) );
na02m06 TIMEBOOST_cell_62532 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_151), .o(TIMEBOOST_net_20213) );
na03m02 TIMEBOOST_cell_72928 ( .a(FE_OFN1678_n_4655), .b(n_4482), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_23295) );
in01m02 g64332_u0 ( .a(FE_OFN1057_n_4727), .o(g64332_sb) );
na02m02 TIMEBOOST_cell_29483 ( .a(configuration_wb_err_addr_533), .b(n_2960), .o(TIMEBOOST_net_8846) );
na02f01 TIMEBOOST_cell_69611 ( .a(TIMEBOOST_net_22013), .b(FE_OFN1034_n_4732), .o(TIMEBOOST_net_20414) );
in01m01 g64333_u0 ( .a(FE_OFN917_n_4725), .o(g64333_sb) );
na03f02 TIMEBOOST_cell_73343 ( .a(n_17048), .b(n_4880), .c(n_17034), .o(TIMEBOOST_net_430) );
na02s01 TIMEBOOST_cell_45543 ( .a(n_351), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q), .o(TIMEBOOST_net_13666) );
in01m01 g64334_u0 ( .a(FE_OFN917_n_4725), .o(g64334_sb) );
na03f02 TIMEBOOST_cell_73690 ( .a(TIMEBOOST_net_22950), .b(g52439_db), .c(TIMEBOOST_net_22959), .o(n_14813) );
na02f02 TIMEBOOST_cell_49156 ( .a(TIMEBOOST_net_14795), .b(g61869_sb), .o(n_8097) );
in01f01 g64335_u0 ( .a(FE_OFN917_n_4725), .o(g64335_sb) );
na03s02 TIMEBOOST_cell_22759 ( .a(FE_OFN270_n_9836), .b(g58088_sb), .c(g58088_db), .o(n_9708) );
in01f02 g64336_u0 ( .a(FE_OFN916_n_4725), .o(g64336_sb) );
na02m10 TIMEBOOST_cell_45545 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q), .o(TIMEBOOST_net_13667) );
na02m04 TIMEBOOST_cell_70235 ( .a(TIMEBOOST_net_22325), .b(FE_OFN719_n_8060), .o(TIMEBOOST_net_15037) );
na03f02 TIMEBOOST_cell_73414 ( .a(TIMEBOOST_net_17386), .b(FE_OFN1196_n_4090), .c(g62573_sb), .o(n_6407) );
in01m06 g64337_u0 ( .a(FE_OFN912_n_4727), .o(g64337_sb) );
na04f02 TIMEBOOST_cell_73415 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q), .b(n_4358), .c(FE_OFN1243_n_4092), .d(g62509_sb), .o(n_6561) );
na02m04 g64337_u2 ( .a(FE_OFN912_n_4727), .b(pci_target_unit_fifos_pciw_addr_data_in_151), .o(g64337_db) );
na02m01 TIMEBOOST_cell_69818 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q), .o(TIMEBOOST_net_22117) );
oa12m01 g64338_u0 ( .a(n_3797), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_3__270), .c(n_4725), .o(n_4726) );
in01m02 g64339_u0 ( .a(FE_OFN1057_n_4727), .o(g64339_sb) );
na04f04 TIMEBOOST_cell_67544 ( .a(g61881_sb), .b(FE_OFN706_n_8119), .c(n_1864), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q), .o(n_8068) );
na03f08 TIMEBOOST_cell_64313 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q), .b(n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_414), .o(TIMEBOOST_net_14864) );
na02s01 TIMEBOOST_cell_70268 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q), .o(TIMEBOOST_net_22342) );
in01m02 g64340_u0 ( .a(FE_OFN918_n_4725), .o(g64340_sb) );
na02m02 TIMEBOOST_cell_70217 ( .a(TIMEBOOST_net_22316), .b(g61912_sb), .o(n_7997) );
na03m02 TIMEBOOST_cell_72475 ( .a(TIMEBOOST_net_16566), .b(FE_OFN905_n_4736), .c(g64126_sb), .o(TIMEBOOST_net_13112) );
in01f01 g64341_u0 ( .a(FE_OFN1056_n_4727), .o(g64341_sb) );
na02m06 TIMEBOOST_cell_68570 ( .a(FE_OFN625_n_4409), .b(n_156), .o(TIMEBOOST_net_21493) );
in01m02 g64342_u0 ( .a(FE_OFN1056_n_4727), .o(g64342_sb) );
na04f04 TIMEBOOST_cell_73441 ( .a(n_3768), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q), .c(FE_OFN1216_n_4151), .d(g62359_sb), .o(n_6880) );
na03f02 TIMEBOOST_cell_73523 ( .a(TIMEBOOST_net_13359), .b(n_6645), .c(g62400_sb), .o(n_6799) );
na02s02 TIMEBOOST_cell_48876 ( .a(TIMEBOOST_net_14655), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_10857) );
in01f02 g64343_u0 ( .a(FE_OFN918_n_4725), .o(g64343_sb) );
na03f02 TIMEBOOST_cell_68380 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q), .b(FE_OFN906_n_4736), .c(pci_target_unit_fifos_pciw_addr_data_in_148), .o(TIMEBOOST_net_21398) );
na04m02 TIMEBOOST_cell_67413 ( .a(TIMEBOOST_net_14517), .b(FE_OFN1676_n_4655), .c(g65365_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q), .o(TIMEBOOST_net_16776) );
na02m02 TIMEBOOST_cell_68405 ( .a(TIMEBOOST_net_21410), .b(TIMEBOOST_net_16189), .o(TIMEBOOST_net_13094) );
in01m02 g64344_u0 ( .a(FE_OFN917_n_4725), .o(g64344_sb) );
na03s01 TIMEBOOST_cell_22767 ( .a(FE_OFN270_n_9836), .b(g58056_sb), .c(g58056_db), .o(n_9733) );
na02f01 TIMEBOOST_cell_70610 ( .a(TIMEBOOST_net_13039), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_22513) );
in01m10 g64345_u0 ( .a(FE_OFN918_n_4725), .o(g64345_sb) );
in01m01 g64346_u0 ( .a(FE_OFN930_n_4730), .o(g64346_sb) );
na03f02 TIMEBOOST_cell_34848 ( .a(TIMEBOOST_net_9429), .b(FE_OFN1421_n_8567), .c(g57351_sb), .o(n_11398) );
na04f06 TIMEBOOST_cell_73177 ( .a(TIMEBOOST_net_17282), .b(FE_OFN1150_n_13249), .c(n_2116), .d(g54140_sb), .o(n_13667) );
in01m01 g64347_u0 ( .a(FE_OFN1055_n_4727), .o(g64347_sb) );
na02s02 TIMEBOOST_cell_70869 ( .a(TIMEBOOST_net_22642), .b(FE_OFN569_n_9528), .o(TIMEBOOST_net_16762) );
na02s01 TIMEBOOST_cell_45461 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q), .o(TIMEBOOST_net_13625) );
in01m02 g64348_u0 ( .a(FE_OFN917_n_4725), .o(g64348_sb) );
na03s02 TIMEBOOST_cell_22771 ( .a(FE_OFN260_n_9860), .b(g58041_sb), .c(g58041_db), .o(n_9747) );
na02m01 TIMEBOOST_cell_54025 ( .a(FE_OFN686_n_4417), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q), .o(TIMEBOOST_net_17230) );
na03f02 TIMEBOOST_cell_34943 ( .a(TIMEBOOST_net_8563), .b(FE_OFN1398_n_8567), .c(g58574_sb), .o(n_9194) );
in01m01 g64349_u0 ( .a(FE_OFN1031_n_4732), .o(g64349_sb) );
na02s01 TIMEBOOST_cell_62992 ( .a(configuration_wb_err_cs_bit31_24), .b(conf_wb_err_bc_in), .o(TIMEBOOST_net_20443) );
na02f01 g64349_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(FE_OFN1031_n_4732), .o(g64349_db) );
na02m06 g64866_u2 ( .a(FE_OFN612_n_4501), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q), .o(g64866_db) );
in01m01 g64350_u0 ( .a(FE_OFN930_n_4730), .o(g64350_sb) );
in01s01 TIMEBOOST_cell_63609 ( .a(TIMEBOOST_net_20789), .o(TIMEBOOST_net_20788) );
na02s01 TIMEBOOST_cell_44023 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q), .b(FE_OFN585_n_9692), .o(TIMEBOOST_net_12906) );
in01m01 g64351_u0 ( .a(FE_OFN917_n_4725), .o(g64351_sb) );
na02f40 TIMEBOOST_cell_45003 ( .a(n_7398), .b(n_16914), .o(TIMEBOOST_net_13396) );
na02s01 TIMEBOOST_cell_48880 ( .a(TIMEBOOST_net_14657), .b(FE_OFN247_n_9112), .o(TIMEBOOST_net_9439) );
na03f02 TIMEBOOST_cell_66597 ( .a(TIMEBOOST_net_17008), .b(FE_OFN1208_n_6356), .c(g62578_sb), .o(n_6398) );
in01m01 g64352_u0 ( .a(FE_OFN918_n_4725), .o(g64352_sb) );
na02m01 g64352_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(FE_OFN918_n_4725), .o(g64352_db) );
na02m02 TIMEBOOST_cell_44911 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q), .b(g58289_sb), .o(TIMEBOOST_net_13350) );
in01m02 g64353_u0 ( .a(FE_OFN916_n_4725), .o(g64353_sb) );
na03s01 TIMEBOOST_cell_22774 ( .a(g58027_db), .b(g58027_sb), .c(FE_OFN270_n_9836), .o(n_9761) );
na02f04 TIMEBOOST_cell_71449 ( .a(TIMEBOOST_net_22932), .b(FE_RN_571_0), .o(FE_RN_573_0) );
in01f01 g64354_u0 ( .a(FE_OFN918_n_4725), .o(g64354_sb) );
na03s01 TIMEBOOST_cell_22777 ( .a(g58010_db), .b(g58010_sb), .c(FE_OFN260_n_9860), .o(n_9783) );
na02f02 g64354_u2 ( .a(FE_OFN918_n_4725), .b(pci_target_unit_fifos_pciw_addr_data_in_125), .o(g64354_db) );
na03m02 TIMEBOOST_cell_73010 ( .a(TIMEBOOST_net_21867), .b(FE_OFN1809_n_4454), .c(TIMEBOOST_net_22105), .o(TIMEBOOST_net_17516) );
in01m02 g64355_u0 ( .a(FE_OFN916_n_4725), .o(g64355_sb) );
na03f02 TIMEBOOST_cell_67642 ( .a(TIMEBOOST_net_15565), .b(FE_OFN1274_n_4096), .c(g62362_sb), .o(n_7392) );
na03s02 TIMEBOOST_cell_72431 ( .a(FE_OFN602_n_9687), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q), .c(TIMEBOOST_net_22341), .o(TIMEBOOST_net_20424) );
in01m02 g64356_u0 ( .a(FE_OFN916_n_4725), .o(g64356_sb) );
na04f02 TIMEBOOST_cell_67927 ( .a(n_3296), .b(n_2622), .c(n_3374), .d(n_3399), .o(n_5549) );
na02m02 TIMEBOOST_cell_62502 ( .a(n_3783), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q), .o(TIMEBOOST_net_20198) );
in01m01 g64357_u0 ( .a(FE_OFN918_n_4725), .o(g64357_sb) );
na02m01 TIMEBOOST_cell_64110 ( .a(n_13541), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q), .o(TIMEBOOST_net_21041) );
na02f02 TIMEBOOST_cell_70852 ( .a(TIMEBOOST_net_16696), .b(FE_OFN1302_n_5763), .o(TIMEBOOST_net_22634) );
na02s02 TIMEBOOST_cell_52730 ( .a(TIMEBOOST_net_16582), .b(g58102_db), .o(n_9696) );
in01m01 g64358_u0 ( .a(FE_OFN918_n_4725), .o(g64358_sb) );
na02s01 TIMEBOOST_cell_42809 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q), .o(TIMEBOOST_net_12299) );
na02m01 g64358_u2 ( .a(pci_target_unit_fifos_pciw_cbe_in), .b(FE_OFN918_n_4725), .o(g64358_db) );
na03f02 TIMEBOOST_cell_67079 ( .a(FE_OFN1596_n_13741), .b(n_13873), .c(TIMEBOOST_net_13799), .o(n_14264) );
in01m01 g64359_u0 ( .a(FE_OFN918_n_4725), .o(g64359_sb) );
na02m04 TIMEBOOST_cell_72304 ( .a(FE_OFN272_n_9828), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q), .o(TIMEBOOST_net_23360) );
in01m02 g64360_u0 ( .a(FE_OFN916_n_4725), .o(g64360_sb) );
na04m06 TIMEBOOST_cell_72740 ( .a(n_4470), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q), .c(FE_OFN640_n_4669), .d(TIMEBOOST_net_21883), .o(TIMEBOOST_net_17549) );
in01m02 g64361_u0 ( .a(FE_OFN918_n_4725), .o(g64361_sb) );
na02s01 TIMEBOOST_cell_52326 ( .a(TIMEBOOST_net_16380), .b(g58059_sb), .o(TIMEBOOST_net_9494) );
in01m02 g64362_u0 ( .a(FE_OFN918_n_4725), .o(g64362_sb) );
na04f02 TIMEBOOST_cell_36820 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q), .b(FE_OFN1379_n_8567), .c(n_9454), .d(FE_OFN1426_n_8567), .o(n_11224) );
na03s02 TIMEBOOST_cell_71944 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q), .b(FE_OFN685_n_4417), .c(n_4493), .o(TIMEBOOST_net_23180) );
na04f02 TIMEBOOST_cell_36822 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q), .b(FE_OFN1379_n_8567), .c(n_9201), .d(FE_OFN1426_n_8567), .o(n_10800) );
in01m02 g64363_u0 ( .a(FE_OFN916_n_4725), .o(g64363_sb) );
na02m02 TIMEBOOST_cell_68732 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q), .b(g64825_sb), .o(TIMEBOOST_net_21574) );
na03s02 TIMEBOOST_cell_22792 ( .a(g57924_sb), .b(FE_OFN264_n_9849), .c(g57924_db), .o(n_9886) );
oa12m02 g64364_u0 ( .a(n_3808), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_0__153), .c(FE_OFN1059_n_4727), .o(n_4722) );
na03f02 TIMEBOOST_cell_65881 ( .a(TIMEBOOST_net_16361), .b(g64349_db), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q), .o(TIMEBOOST_net_14891) );
na02s01 TIMEBOOST_cell_39742 ( .a(FE_OFN201_n_9230), .b(g57903_sb), .o(TIMEBOOST_net_11483) );
in01f01 g64366_u0 ( .a(FE_OFN1033_n_4732), .o(g64366_sb) );
na04f04 TIMEBOOST_cell_42519 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_786), .c(FE_OFN2134_n_13124), .d(g54351_sb), .o(n_13090) );
na02f01 TIMEBOOST_cell_72242 ( .a(TIMEBOOST_net_13052), .b(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_23329) );
na04m04 TIMEBOOST_cell_67860 ( .a(TIMEBOOST_net_14263), .b(FE_OFN929_n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q), .d(g64301_sb), .o(TIMEBOOST_net_8324) );
in01f01 g64367_u0 ( .a(FE_OFN918_n_4725), .o(g64367_sb) );
na02m01 TIMEBOOST_cell_69096 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q), .b(FE_OFN1663_n_4490), .o(TIMEBOOST_net_21756) );
na04f02 TIMEBOOST_cell_36824 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN1394_n_8567), .c(n_8556), .d(g58592_sb), .o(n_8906) );
no02f02 g64368_u0 ( .a(wbu_addr_in_260), .b(n_2694), .o(g64368_p) );
ao12f02 g64368_u1 ( .a(g64368_p), .b(wbu_addr_in_260), .c(n_2694), .o(n_2695) );
no02m02 g64369_u0 ( .a(n_2419), .b(wbm_adr_o_11_), .o(g64369_p) );
ao12f02 g64369_u1 ( .a(g64369_p), .b(wbm_adr_o_11_), .c(n_2419), .o(n_2693) );
no02f04 g64370_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_9_), .b(n_1633), .o(g64370_p) );
ao12f02 g64370_u1 ( .a(g64370_p), .b(pci_target_unit_del_sync_comp_cycle_count_9_), .c(n_1633), .o(n_2423) );
no02m04 g64371_u0 ( .a(n_1992), .b(n_1631), .o(g64371_p) );
ao12f02 g64371_u1 ( .a(g64371_p), .b(n_1992), .c(n_1631), .o(n_2422) );
in01f01 g64372_u0 ( .a(n_1669), .o(n_1463) );
in01s01 g64373_u0 ( .a(n_1438), .o(n_1190) );
in01s01 g64374_u0 ( .a(n_1476), .o(n_1213) );
no02f04 g64375_u0 ( .a(conf_wb_err_addr_in_952), .b(n_2691), .o(g64375_p) );
ao12f02 g64375_u1 ( .a(g64375_p), .b(conf_wb_err_addr_in_952), .c(n_2691), .o(n_2692) );
no02f04 g64376_u0 ( .a(conf_wb_err_addr_in_949), .b(n_2260), .o(g64376_p) );
ao12f02 g64376_u1 ( .a(g64376_p), .b(conf_wb_err_addr_in_949), .c(n_2260), .o(n_2261) );
no02f04 g64377_u0 ( .a(wbm_adr_o_8_), .b(n_2258), .o(g64377_p) );
ao12f02 g64377_u1 ( .a(g64377_p), .b(wbm_adr_o_8_), .c(n_2258), .o(n_2259) );
no02s01 g64378_u0 ( .a(n_2256), .b(wbu_addr_in_257), .o(g64378_p) );
ao12s01 g64378_u1 ( .a(g64378_p), .b(wbu_addr_in_257), .c(n_2256), .o(n_2257) );
no02f08 g64379_u0 ( .a(n_1396), .b(n_1395), .o(g64379_p) );
ao12f08 g64379_u1 ( .a(g64379_p), .b(n_1396), .c(n_1395), .o(n_2255) );
no02f08 g64380_u0 ( .a(n_1393), .b(n_1404), .o(g64380_p) );
ao12f06 g64380_u1 ( .a(g64380_p), .b(n_1393), .c(n_1404), .o(n_2254) );
no02f08 g64382_u0 ( .a(n_1400), .b(n_1398), .o(g64382_p) );
ao12f08 g64382_u1 ( .a(g64382_p), .b(n_1400), .c(n_1398), .o(n_2252) );
no02f08 g64383_u0 ( .a(n_1449), .b(n_1405), .o(g64383_p) );
ao12f08 g64383_u1 ( .a(g64383_p), .b(n_1449), .c(n_1405), .o(n_2251) );
no02f10 g64384_u0 ( .a(n_1402), .b(n_1401), .o(g64384_p) );
ao12f08 g64384_u1 ( .a(g64384_p), .b(n_1402), .c(n_1401), .o(n_2250) );
no02f06 g64385_u0 ( .a(n_1394), .b(n_1439), .o(g64385_p) );
ao12f06 g64385_u1 ( .a(g64385_p), .b(n_1394), .c(n_1439), .o(n_2249) );
na02f06 g64450_u0 ( .a(n_2219), .b(pci_gnt_i), .o(n_3126) );
na02f02 g64451_u0 ( .a(n_3115), .b(configuration_icr_bit2_0), .o(n_2898) );
na02f06 g64452_u0 ( .a(n_3290), .b(pciu_bar0_in_364), .o(n_3292) );
na02f01 g64454_u0 ( .a(n_4718), .b(n_3314), .o(g64454_p) );
in01f02 g64454_u1 ( .a(g64454_p), .o(n_3289) );
na03f02 TIMEBOOST_cell_73670 ( .a(TIMEBOOST_net_8331), .b(FE_OFN2106_g64577_p), .c(g63099_sb), .o(n_5056) );
na02m01 g64456_u0 ( .a(n_4512), .b(n_4669), .o(n_4514) );
na02m04 TIMEBOOST_cell_69551 ( .a(TIMEBOOST_net_21983), .b(TIMEBOOST_net_12689), .o(TIMEBOOST_net_17494) );
na02m01 TIMEBOOST_cell_47559 ( .a(g58789_sb), .b(n_8831), .o(TIMEBOOST_net_13997) );
no02f03 g64459_u0 ( .a(n_2726), .b(n_3023), .o(n_3812) );
na02m01 g64460_u0 ( .a(n_4512), .b(n_4677), .o(n_4513) );
no02m06 g64461_u0 ( .a(n_2248), .b(n_1621), .o(g64461_p) );
in01m04 g64461_u1 ( .a(g64461_p), .o(n_7835) );
na02m01 g64462_u0 ( .a(n_4512), .b(FE_OFN1678_n_4655), .o(n_4511) );
na02f01 g64463_u0 ( .a(n_4512), .b(FE_OFN1640_n_4671), .o(n_4510) );
no02f20 g64464_u0 ( .a(n_15324), .b(n_2308), .o(n_2897) );
no02f02 g64465_u0 ( .a(n_3016), .b(n_2449), .o(g64465_p) );
in01f02 g64465_u1 ( .a(g64465_p), .o(n_3390) );
no02m04 g64466_u0 ( .a(n_1623), .b(n_4725), .o(g64466_p) );
in01m02 g64466_u1 ( .a(g64466_p), .o(n_2247) );
na02s01 TIMEBOOST_cell_42798 ( .a(TIMEBOOST_net_12293), .b(FE_OFN936_n_2292), .o(TIMEBOOST_net_10232) );
na02f40 g64577_u0 ( .a(n_2399), .b(pci_target_unit_fifos_pciw_wenable_in), .o(g64577_p) );
na02f08 g64578_u0 ( .a(n_1482), .b(n_2691), .o(g64578_p) );
in01f06 g64578_u1 ( .a(g64578_p), .o(n_3130) );
na03m02 TIMEBOOST_cell_67158 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q), .b(n_3792), .c(FE_OFN1640_n_4671), .o(TIMEBOOST_net_14441) );
na02m01 g64580_u0 ( .a(n_4512), .b(FE_OFN651_n_4508), .o(n_4509) );
na02f10 g64581_u0 ( .a(n_1388), .b(n_2260), .o(g64581_p) );
in01f08 g64581_u1 ( .a(g64581_p), .o(n_2722) );
na02f04 g64582_u0 ( .a(n_1437), .b(pci_target_unit_wishbone_master_rty_counter_3_), .o(g64582_p) );
in01f04 g64582_u1 ( .a(g64582_p), .o(n_1273) );
na02f10 g64583_u0 ( .a(n_3023), .b(FE_OFN2121_n_2687), .o(n_6986) );
in01f01 g64584_u0 ( .a(n_3313), .o(n_2888) );
na02f40 g64585_u0 ( .a(n_4718), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(g64585_p) );
in01f10 g64585_u1 ( .a(g64585_p), .o(n_3313) );
na03m02 TIMEBOOST_cell_46696 ( .a(TIMEBOOST_net_12805), .b(g58379_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q), .o(TIMEBOOST_net_9466) );
no02f02 g64587_u0 ( .a(FE_OFN2100_n_3281), .b(n_3280), .o(g64587_p) );
in01f02 g64587_u1 ( .a(g64587_p), .o(n_3282) );
in01s01 g64588_u0 ( .a(n_2245), .o(n_2246) );
no02f04 g64589_u0 ( .a(n_3395), .b(FE_OFN999_n_15978), .o(n_2245) );
na02f08 g64590_u0 ( .a(n_3089), .b(n_2308), .o(n_3090) );
no02f02 g64591_u0 ( .a(n_3388), .b(n_3275), .o(n_3389) );
no02m01 g64592_u0 ( .a(n_3388), .b(n_3265), .o(n_3387) );
no02f02 g64593_u0 ( .a(n_3278), .b(n_3277), .o(n_3279) );
na02f06 g64595_u0 ( .a(n_4718), .b(n_2685), .o(g64595_p) );
in01f06 g64595_u1 ( .a(g64595_p), .o(n_3119) );
na02f10 g64596_u0 ( .a(n_1282), .b(n_2256), .o(g64596_p) );
in01f08 g64596_u1 ( .a(g64596_p), .o(n_2437) );
na02f10 g64597_u0 ( .a(n_1373), .b(n_2419), .o(g64597_p) );
in01f08 g64597_u1 ( .a(g64597_p), .o(n_2931) );
oa12f01 g64598_u0 ( .a(n_2406), .b(n_990), .c(n_691), .o(n_2418) );
na02f01 g64599_u0 ( .a(n_3810), .b(n_4084), .o(n_3811) );
no02f02 g64601_u0 ( .a(n_3278), .b(n_3275), .o(n_3276) );
no02f80 g64602_u0 ( .a(pci_target_unit_pci_target_sm_state_transfere_reg), .b(n_532), .o(n_2887) );
in01f01 g64603_u0 ( .a(n_4533), .o(n_3809) );
na02m02 g64605_u0 ( .a(FE_OFN1059_n_4727), .b(n_3806), .o(n_3808) );
no02m02 g64606_u0 ( .a(n_3386), .b(n_3395), .o(n_3385) );
no02m01 g64607_u0 ( .a(n_3388), .b(n_3273), .o(n_3384) );
no02f01 g64608_u0 ( .a(n_3278), .b(n_3273), .o(n_3274) );
na02m02 g64609_u0 ( .a(n_4730), .b(n_3806), .o(n_3807) );
no02f08 g64610_u0 ( .a(n_13820), .b(n_2415), .o(g64610_p) );
in01f04 g64610_u1 ( .a(g64610_p), .o(n_2416) );
na02m06 g64611_u0 ( .a(FE_OFN1036_n_4732), .b(n_3806), .o(n_3805) );
na04f04 TIMEBOOST_cell_24209 ( .a(n_9517), .b(g57423_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q), .d(FE_OFN1424_n_8567), .o(n_11314) );
na03s02 TIMEBOOST_cell_72442 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(FE_OFN946_n_2248), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q), .o(TIMEBOOST_net_21406) );
na04f04 TIMEBOOST_cell_73260 ( .a(TIMEBOOST_net_20413), .b(TIMEBOOST_net_11010), .c(FE_OFN1095_g64577_p), .d(g61963_sb), .o(n_6948) );
in01s02 g64630_u3 ( .a(g64630_p), .o(n_1995) );
na02f04 g64631_u0 ( .a(n_3089), .b(n_2742), .o(g64631_p) );
in01f02 g64631_u1 ( .a(g64631_p), .o(n_3271) );
no02m02 g64632_u0 ( .a(n_3798), .b(n_2464), .o(g64632_p) );
in01s02 g64632_u1 ( .a(g64632_p), .o(n_3800) );
na02f08 g64633_u0 ( .a(n_2694), .b(n_1479), .o(g64633_p) );
in01f06 g64633_u1 ( .a(g64633_p), .o(n_3132) );
no02f10 g64639_u0 ( .a(n_3278), .b(n_3030), .o(g64639_p) );
in01f08 g64639_u1 ( .a(g64639_p), .o(n_4630) );
no02f02 g64641_u0 ( .a(n_3798), .b(n_2319), .o(n_3799) );
no02f01 g64642_u0 ( .a(n_4720), .b(n_3280), .o(n_4721) );
na02f10 g64643_u0 ( .a(n_1241), .b(n_2258), .o(g64643_p) );
in01f10 g64643_u1 ( .a(g64643_p), .o(n_2441) );
no02f40 g64644_u0 ( .a(n_842), .b(n_938), .o(n_1434) );
no02f08 g64645_u0 ( .a(n_1987), .b(n_1974), .o(n_2414) );
no02f01 g64646_u0 ( .a(n_4718), .b(n_691), .o(g64646_p) );
in01f02 g64646_u1 ( .a(g64646_p), .o(n_3087) );
na02m02 g64647_u0 ( .a(n_4725), .b(n_3806), .o(n_3797) );
na02s01 g64649_u0 ( .a(n_3267), .b(n_2966), .o(n_3268) );
no02f10 g64650_u0 ( .a(n_3395), .b(n_1514), .o(n_2443) );
no02f01 g64651_u0 ( .a(n_3278), .b(n_3265), .o(n_3266) );
no02f02 g64652_u0 ( .a(n_3388), .b(n_3277), .o(n_3381) );
in01f20 g64667_u0 ( .a(n_15260), .o(n_13249) );
na02f02 g64670_u0 ( .a(n_1961), .b(n_2337), .o(n_4152) );
no02f08 g64671_u0 ( .a(n_3388), .b(n_3030), .o(g64671_p) );
in01f06 g64671_u1 ( .a(g64671_p), .o(n_4783) );
in01m02 g64676_u0 ( .a(n_2727), .o(n_2412) );
ao12f10 g64677_u0 ( .a(n_1588), .b(n_1211), .c(n_545), .o(n_2727) );
na02f04 g64678_u0 ( .a(n_1533), .b(n_3795), .o(g64678_p) );
in01f02 g64678_u1 ( .a(g64678_p), .o(n_3796) );
na02s02 TIMEBOOST_cell_39179 ( .a(TIMEBOOST_net_11201), .b(g58217_db), .o(n_9569) );
na04s02 TIMEBOOST_cell_72906 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q), .b(g65822_sb), .c(g65822_db), .d(TIMEBOOST_net_14826), .o(n_8071) );
ao12s01 g64685_u0 ( .a(pci_target_unit_del_sync_req_comp_pending), .b(pci_target_unit_del_sync_req_rty_exp_reg), .c(pci_target_unit_del_sync_req_rty_exp_clr), .o(n_646) );
no02f02 g64687_u0 ( .a(n_2070), .b(n_3261), .o(g64687_p) );
in01f02 g64687_u1 ( .a(g64687_p), .o(n_3262) );
na03s02 TIMEBOOST_cell_64466 ( .a(TIMEBOOST_net_10238), .b(g65699_sb), .c(TIMEBOOST_net_20846), .o(n_8368) );
ao12s01 g64689_u0 ( .a(n_152), .b(n_2765), .c(output_backup_trdy_out_reg_Q), .o(n_3380) );
na02f01 g64694_u0 ( .a(n_2303), .b(n_4718), .o(g64694_p) );
in01f01 g64694_u1 ( .a(g64694_p), .o(n_3081) );
oa12m01 g64695_u0 ( .a(n_2803), .b(n_15762), .c(n_3022), .o(n_2900) );
na03f10 TIMEBOOST_cell_64292 ( .a(n_1441), .b(n_529), .c(n_2982), .o(TIMEBOOST_net_185) );
na02m02 g64697_u0 ( .a(n_3481), .b(n_4718), .o(g64697_p) );
in01m02 g64697_u1 ( .a(g64697_p), .o(n_4719) );
ao22f02 g64698_u0 ( .a(n_2555), .b(n_14909), .c(n_2358), .d(n_2331), .o(n_3259) );
ao12f04 g64699_u0 ( .a(n_2086), .b(n_3123), .c(n_1554), .o(n_2878) );
na02f02 g64700_u0 ( .a(n_2065), .b(FE_OFN197_n_2683), .o(g64700_p) );
in01f02 g64700_u1 ( .a(g64700_p), .o(n_2684) );
no02f02 g64701_u0 ( .a(n_2072), .b(n_3261), .o(g64701_p) );
in01f02 g64701_u1 ( .a(g64701_p), .o(n_3258) );
no02f04 g64702_u0 ( .a(n_3261), .b(n_2068), .o(g64702_p) );
in01f02 g64702_u1 ( .a(g64702_p), .o(n_3257) );
ao12f02 g64703_u0 ( .a(n_2409), .b(n_8498), .c(pci_target_unit_pcit_if_req_req_pending_in), .o(n_2410) );
no02f01 g64704_u0 ( .a(n_3261), .b(n_8540), .o(g64704_p) );
in01f01 g64704_u1 ( .a(g64704_p), .o(n_3256) );
no02f02 g64705_u0 ( .a(n_2080), .b(n_3261), .o(g64705_p) );
in01f02 g64705_u1 ( .a(g64705_p), .o(n_3255) );
ao12s01 g64706_u0 ( .a(n_1659), .b(wishbone_slave_unit_pci_initiator_if_read_count_2_), .c(n_660), .o(n_1660) );
na02f08 g64707_u0 ( .a(n_3163), .b(n_3378), .o(g64707_p) );
in01f06 g64707_u1 ( .a(g64707_p), .o(n_3379) );
no02f06 g64708_u0 ( .a(n_1832), .b(n_1834), .o(n_8564) );
ao12m01 g64709_u0 ( .a(n_1178), .b(n_1011), .c(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(n_1658) );
in01s01 g64710_u0 ( .a(n_2682), .o(n_2877) );
ao12s01 g64711_u0 ( .a(wishbone_slave_unit_del_sync_req_comp_pending), .b(wishbone_slave_unit_del_sync_req_rty_exp_reg), .c(wishbone_slave_unit_del_sync_req_rty_exp_clr), .o(n_2682) );
no02f01 g64712_u0 ( .a(n_2079), .b(n_3261), .o(g64712_p) );
in01f01 g64712_u1 ( .a(g64712_p), .o(n_3254) );
oa12f01 g64714_u0 ( .a(n_2406), .b(wishbone_slave_unit_pci_initiator_if_read_count_0_), .c(n_691), .o(n_2407) );
oa12f02 g64715_u0 ( .a(n_2406), .b(n_292), .c(n_692), .o(n_2405) );
ao12f02 g64716_u0 ( .a(n_2049), .b(wbu_cache_line_size_in_206), .c(n_691), .o(n_2234) );
na02f02 TIMEBOOST_cell_38247 ( .a(TIMEBOOST_net_10735), .b(g65709_db), .o(n_1946) );
na04f04 TIMEBOOST_cell_24191 ( .a(n_8557), .b(g58591_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q), .d(FE_OFN1403_n_8567), .o(n_8908) );
na03f04 TIMEBOOST_cell_73181 ( .a(TIMEBOOST_net_23279), .b(g64297_sb), .c(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_22455) );
na02s01 TIMEBOOST_cell_18561 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q), .b(FE_OFN2079_n_8069), .o(TIMEBOOST_net_5644) );
na02f04 g64727_u0 ( .a(n_2399), .b(n_1976), .o(g64727_p) );
in01f04 g64727_u1 ( .a(g64727_p), .o(n_3335) );
oa22f08 g64728_u0 ( .a(n_1809), .b(n_16168), .c(n_16160), .d(n_3250), .o(n_5751) );
ao12f04 g64729_u0 ( .a(n_3026), .b(n_16000), .c(n_3078), .o(n_3079) );
na04f02 TIMEBOOST_cell_73416 ( .a(n_4382), .b(FE_OFN1223_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q), .d(g62649_sb), .o(n_6249) );
na04f04 TIMEBOOST_cell_25003 ( .a(n_10614), .b(n_9260), .c(n_10026), .d(n_10023), .o(n_12144) );
na03f02 TIMEBOOST_cell_73824 ( .a(TIMEBOOST_net_13801), .b(n_13903), .c(FE_OFN1596_n_13741), .o(n_14302) );
na03s02 TIMEBOOST_cell_73011 ( .a(TIMEBOOST_net_20824), .b(g65758_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q), .o(TIMEBOOST_net_23364) );
ao22f04 g64735_u0 ( .a(n_2339), .b(n_14910), .c(configuration_wb_err_data_572), .d(FE_OFN1071_n_15729), .o(n_3077) );
no02s01 g64736_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_5_), .b(n_1425), .o(g64736_p) );
ao12s01 g64736_u1 ( .a(g64736_p), .b(pci_target_unit_del_sync_comp_cycle_count_5_), .c(n_1425), .o(n_1701) );
ao22s01 g64738_u0 ( .a(n_547), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_2_), .c(n_401), .d(n_1471), .o(n_1472) );
ao12f01 g64739_u0 ( .a(n_2806), .b(pci_target_unit_wishbone_master_read_count_1_), .c(n_3250), .o(n_3251) );
no02f02 g64740_u0 ( .a(n_1469), .b(pci_target_unit_wishbone_master_rty_counter_5_), .o(g64740_p) );
ao12f02 g64740_u1 ( .a(g64740_p), .b(pci_target_unit_wishbone_master_rty_counter_5_), .c(n_1469), .o(n_2291) );
oa12f02 g64741_u0 ( .a(n_2002), .b(n_2001), .c(pci_target_unit_wishbone_master_rty_counter_6_), .o(n_2396) );
ao22f02 g64742_u0 ( .a(configuration_isr_bit_631), .b(n_3246), .c(n_3248), .d(configuration_sync_command_bit0), .o(n_15436) );
in01s01 g64743_u0 ( .a(n_3377), .o(n_3794) );
na02f01 TIMEBOOST_cell_68167 ( .a(TIMEBOOST_net_21291), .b(wbu_addr_in_276), .o(TIMEBOOST_net_12305) );
ao22f01 g64745_u0 ( .a(configuration_command_bit), .b(n_3248), .c(n_3246), .d(configuration_isr_bit_618), .o(n_3247) );
no02m01 g64746_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_5_), .b(n_1426), .o(g64746_p) );
ao12m01 g64746_u1 ( .a(g64746_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_5_), .c(n_1426), .o(n_1656) );
no02f06 g64747_u0 ( .a(n_1279), .b(n_1081), .o(g64747_p) );
ao12f08 g64747_u1 ( .a(g64747_p), .b(n_1081), .c(n_1279), .o(n_2227) );
in01m01 g64748_u0 ( .a(FE_OFN672_n_4505), .o(g64748_sb) );
na02s02 TIMEBOOST_cell_38563 ( .a(TIMEBOOST_net_10893), .b(g58191_db), .o(n_9593) );
na03m06 TIMEBOOST_cell_72618 ( .a(FE_OFN1013_n_4734), .b(TIMEBOOST_net_20256), .c(g63545_sb), .o(n_4611) );
in01m02 g64749_u0 ( .a(FE_OFN682_n_4460), .o(g64749_sb) );
na04f02 TIMEBOOST_cell_36826 ( .a(n_354), .b(FE_OFN1394_n_8567), .c(n_8549), .d(g58607_sb), .o(n_8900) );
in01m01 g64750_u0 ( .a(FE_OFN671_n_4505), .o(g64750_sb) );
na02s01 TIMEBOOST_cell_49445 ( .a(FE_OFN262_n_9851), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_14940) );
na03f02 TIMEBOOST_cell_73196 ( .a(TIMEBOOST_net_20877), .b(FE_OFN1092_g64577_p), .c(g63573_sb), .o(n_4108) );
in01s01 TIMEBOOST_cell_73921 ( .a(TIMEBOOST_net_23485), .o(TIMEBOOST_net_23486) );
in01m02 g64751_u0 ( .a(FE_OFN614_n_4501), .o(g64751_sb) );
na04f02 TIMEBOOST_cell_68013 ( .a(n_3931), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q), .c(g62777_sb), .d(FE_OFN1140_g64577_p), .o(n_4993) );
na03m02 TIMEBOOST_cell_72805 ( .a(n_4452), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q), .c(TIMEBOOST_net_12596), .o(TIMEBOOST_net_20531) );
na02m10 TIMEBOOST_cell_52447 ( .a(configuration_pci_err_addr_487), .b(wbm_adr_o_17_), .o(TIMEBOOST_net_16441) );
in01s01 g64752_u0 ( .a(FE_OFN678_n_4460), .o(g64752_sb) );
na04f04 TIMEBOOST_cell_36828 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN1415_n_8567), .c(n_9781), .d(g57143_sb), .o(n_11606) );
na02m01 g64752_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q), .b(FE_OFN678_n_4460), .o(g64752_db) );
in01m06 g64753_u0 ( .a(FE_OFN618_n_4490), .o(g64753_sb) );
na02s02 TIMEBOOST_cell_52230 ( .a(TIMEBOOST_net_16332), .b(TIMEBOOST_net_12327), .o(n_9674) );
na03f02 TIMEBOOST_cell_34752 ( .a(TIMEBOOST_net_9404), .b(FE_OFN1400_n_8567), .c(g57357_sb), .o(n_10386) );
na03f02 TIMEBOOST_cell_66919 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_16497), .c(FE_OFN1513_n_14987), .o(n_12661) );
in01m08 g64754_u0 ( .a(FE_OFN672_n_4505), .o(g64754_sb) );
in01m02 g64755_u0 ( .a(FE_OFN671_n_4505), .o(g64755_sb) );
na02s01 TIMEBOOST_cell_38581 ( .a(TIMEBOOST_net_10902), .b(g58144_db), .o(n_9651) );
na02s02 TIMEBOOST_cell_48581 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q), .o(TIMEBOOST_net_14508) );
na02s01 TIMEBOOST_cell_38583 ( .a(TIMEBOOST_net_10903), .b(g58143_db), .o(n_9069) );
in01m01 g64756_u0 ( .a(FE_OFN619_n_4490), .o(g64756_sb) );
na03f02 TIMEBOOST_cell_34754 ( .a(TIMEBOOST_net_9406), .b(FE_OFN1374_n_8567), .c(g57453_sb), .o(n_11281) );
na03s02 TIMEBOOST_cell_41710 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q), .b(g58329_sb), .c(g58329_db), .o(n_9485) );
in01m01 g64757_u0 ( .a(FE_OFN646_n_4497), .o(g64757_sb) );
na02m02 TIMEBOOST_cell_68115 ( .a(TIMEBOOST_net_21265), .b(g61880_sb), .o(TIMEBOOST_net_17292) );
in01m01 g64758_u0 ( .a(FE_OFN667_n_4495), .o(g64758_sb) );
na03s02 TIMEBOOST_cell_42119 ( .a(g58171_sb), .b(FE_OFN260_n_9860), .c(g58171_db), .o(n_9619) );
na02m02 g64758_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q), .b(FE_OFN667_n_4495), .o(g64758_db) );
na03f02 TIMEBOOST_cell_34869 ( .a(TIMEBOOST_net_9344), .b(FE_OFN1414_n_8567), .c(g57391_sb), .o(n_11352) );
in01m04 g64759_u0 ( .a(FE_OFN670_n_4505), .o(g64759_sb) );
na03f04 TIMEBOOST_cell_73578 ( .a(TIMEBOOST_net_7617), .b(FE_OFN1084_n_13221), .c(g54178_da), .o(TIMEBOOST_net_22889) );
na03f02 TIMEBOOST_cell_66487 ( .a(TIMEBOOST_net_17382), .b(FE_OFN1207_n_6356), .c(g62715_sb), .o(n_6140) );
in01m04 g64760_u0 ( .a(FE_OFN1806_n_4501), .o(g64760_sb) );
na02s01 TIMEBOOST_cell_43019 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_139), .o(TIMEBOOST_net_12404) );
na02m02 TIMEBOOST_cell_69469 ( .a(TIMEBOOST_net_21942), .b(TIMEBOOST_net_16261), .o(TIMEBOOST_net_17562) );
na03f02 TIMEBOOST_cell_66662 ( .a(TIMEBOOST_net_17130), .b(FE_OFN1323_n_6436), .c(g62633_sb), .o(n_6286) );
in01m02 g64761_u0 ( .a(FE_OFN669_n_4505), .o(g64761_sb) );
na03s02 TIMEBOOST_cell_73012 ( .a(TIMEBOOST_net_20823), .b(g65742_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q), .o(TIMEBOOST_net_23363) );
na02f02 TIMEBOOST_cell_68609 ( .a(TIMEBOOST_net_21512), .b(n_3019), .o(TIMEBOOST_net_454) );
in01m04 g64762_u0 ( .a(FE_OFN1663_n_4490), .o(g64762_sb) );
na02m02 TIMEBOOST_cell_68611 ( .a(TIMEBOOST_net_21513), .b(TIMEBOOST_net_12354), .o(TIMEBOOST_net_17519) );
na03m02 TIMEBOOST_cell_66464 ( .a(n_3827), .b(g63127_db), .c(FE_OFN1138_g64577_p), .o(n_4999) );
in01m04 g64763_u0 ( .a(FE_OFN1806_n_4501), .o(g64763_sb) );
in01s01 TIMEBOOST_cell_73922 ( .a(wbm_dat_i_12_), .o(TIMEBOOST_net_23487) );
na02f04 TIMEBOOST_cell_68069 ( .a(TIMEBOOST_net_21242), .b(n_928), .o(TIMEBOOST_net_263) );
in01m02 g64764_u0 ( .a(FE_OFN1659_n_4490), .o(g64764_sb) );
na02s01 TIMEBOOST_cell_68293 ( .a(TIMEBOOST_net_21354), .b(TIMEBOOST_net_20161), .o(n_9846) );
na03f02 TIMEBOOST_cell_34756 ( .a(TIMEBOOST_net_9408), .b(FE_OFN1397_n_8567), .c(g57066_sb), .o(n_11676) );
na02f01 TIMEBOOST_cell_44312 ( .a(TIMEBOOST_net_13050), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_11322) );
in01m01 g64765_u0 ( .a(FE_OFN1660_n_4490), .o(g64765_sb) );
na03f02 TIMEBOOST_cell_34758 ( .a(TIMEBOOST_net_9410), .b(FE_OFN1399_n_8567), .c(g57062_sb), .o(n_11677) );
na03f02 TIMEBOOST_cell_73638 ( .a(TIMEBOOST_net_17461), .b(FE_OFN1268_n_4095), .c(g62706_sb), .o(n_6154) );
in01m01 g64766_u0 ( .a(FE_OFN666_n_4495), .o(g64766_sb) );
na03s01 TIMEBOOST_cell_72410 ( .a(wbs_dat_i_31_), .b(g61885_sb), .c(TIMEBOOST_net_9649), .o(TIMEBOOST_net_12834) );
na03m08 TIMEBOOST_cell_72715 ( .a(FE_OFN2108_n_2047), .b(TIMEBOOST_net_20277), .c(g65690_sb), .o(n_1953) );
na03m01 TIMEBOOST_cell_32106 ( .a(g58107_sb), .b(g58107_db), .c(FE_OFN258_n_9862), .o(n_9686) );
in01m01 g64767_u0 ( .a(FE_OFN620_n_4490), .o(g64767_sb) );
na02m02 TIMEBOOST_cell_68295 ( .a(TIMEBOOST_net_21355), .b(n_1079), .o(TIMEBOOST_net_21060) );
na02m04 TIMEBOOST_cell_68750 ( .a(g64895_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q), .o(TIMEBOOST_net_21583) );
in01m04 g64768_u0 ( .a(FE_OFN1660_n_4490), .o(g64768_sb) );
na02f02 TIMEBOOST_cell_71090 ( .a(TIMEBOOST_net_20542), .b(FE_OFN1247_n_4093), .o(TIMEBOOST_net_22753) );
na03f01 TIMEBOOST_cell_72509 ( .a(TIMEBOOST_net_21331), .b(wbu_addr_in_272), .c(g58782_sb), .o(n_9880) );
na02m02 TIMEBOOST_cell_71858 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q), .b(g65962_sb), .o(TIMEBOOST_net_23137) );
in01m02 g64769_u0 ( .a(FE_OFN670_n_4505), .o(g64769_sb) );
na02f02 TIMEBOOST_cell_70349 ( .a(TIMEBOOST_net_22382), .b(g63596_sb), .o(n_7182) );
na03f02 TIMEBOOST_cell_66155 ( .a(TIMEBOOST_net_16744), .b(FE_OFN1184_n_3476), .c(g60653_sb), .o(n_5670) );
na02s02 TIMEBOOST_cell_39746 ( .a(g58307_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q), .o(TIMEBOOST_net_11485) );
in01m01 g64770_u0 ( .a(FE_OFN671_n_4505), .o(g64770_sb) );
na03f02 TIMEBOOST_cell_72874 ( .a(TIMEBOOST_net_21745), .b(g64176_sb), .c(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_22507) );
na03f02 TIMEBOOST_cell_73261 ( .a(TIMEBOOST_net_22313), .b(FE_OFN2212_n_8407), .c(g61733_sb), .o(n_8353) );
in01m01 g64771_u0 ( .a(FE_OFN671_n_4505), .o(g64771_sb) );
no02f02 TIMEBOOST_cell_45411 ( .a(TIMEBOOST_net_7531), .b(FE_RN_374_0), .o(TIMEBOOST_net_13600) );
no02f04 TIMEBOOST_cell_51526 ( .a(TIMEBOOST_net_15980), .b(FE_RN_735_0), .o(n_13787) );
na02s02 TIMEBOOST_cell_38585 ( .a(TIMEBOOST_net_10904), .b(g58092_db), .o(n_9705) );
in01m02 g64772_u0 ( .a(FE_OFN670_n_4505), .o(g64772_sb) );
na02s01 TIMEBOOST_cell_63002 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q), .o(TIMEBOOST_net_20448) );
na03f02 TIMEBOOST_cell_66157 ( .a(TIMEBOOST_net_16434), .b(FE_OFN1185_n_3476), .c(g60645_sb), .o(n_5682) );
na02m02 TIMEBOOST_cell_39748 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q), .b(g58339_sb), .o(TIMEBOOST_net_11486) );
in01m02 g64773_u0 ( .a(FE_OFN670_n_4505), .o(g64773_sb) );
na02s01 TIMEBOOST_cell_38597 ( .a(TIMEBOOST_net_10910), .b(g58014_db), .o(n_9779) );
na02m02 TIMEBOOST_cell_68444 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q), .b(FE_OFN669_n_4505), .o(TIMEBOOST_net_21430) );
na04s02 TIMEBOOST_cell_46767 ( .a(g57957_db), .b(g57957_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q), .d(FE_OFN266_n_9884), .o(TIMEBOOST_net_9462) );
in01m04 g64774_u0 ( .a(FE_OFN670_n_4505), .o(g64774_sb) );
na04f06 TIMEBOOST_cell_68015 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_410), .b(g54191_sb), .c(TIMEBOOST_net_7609), .d(FE_OFN1085_n_13221), .o(n_13426) );
na02m06 g64774_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q), .b(FE_OFN670_n_4505), .o(g64774_db) );
na03f02 TIMEBOOST_cell_73732 ( .a(TIMEBOOST_net_8602), .b(FE_OFN2209_n_11027), .c(n_12362), .o(n_12806) );
in01m01 g64775_u0 ( .a(FE_OFN672_n_4505), .o(g64775_sb) );
na03f02 TIMEBOOST_cell_72528 ( .a(TIMEBOOST_net_21394), .b(g64119_sb), .c(FE_OFN1137_g64577_p), .o(TIMEBOOST_net_22471) );
na02m02 g64775_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q), .b(FE_OFN670_n_4505), .o(g64775_db) );
na03f03 TIMEBOOST_cell_73733 ( .a(TIMEBOOST_net_13629), .b(FE_OFN2209_n_11027), .c(n_12362), .o(n_16408) );
in01m01 g64776_u0 ( .a(FE_OFN671_n_4505), .o(g64776_sb) );
na02f02 TIMEBOOST_cell_50316 ( .a(TIMEBOOST_net_15375), .b(g62364_sb), .o(n_6872) );
na02m02 g64776_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q), .b(FE_OFN671_n_4505), .o(g64776_db) );
na03f02 TIMEBOOST_cell_73417 ( .a(TIMEBOOST_net_20952), .b(FE_OFN1200_n_4090), .c(g62651_sb), .o(n_6243) );
in01m01 g64777_u0 ( .a(FE_OFN671_n_4505), .o(g64777_sb) );
na03m02 TIMEBOOST_cell_73171 ( .a(g64313_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q), .c(TIMEBOOST_net_14747), .o(TIMEBOOST_net_8334) );
na02s01 TIMEBOOST_cell_53535 ( .a(pci_target_unit_fifos_inGreyCount_reg_1__Q), .b(n_852), .o(TIMEBOOST_net_16985) );
in01m01 g64778_u0 ( .a(FE_OFN670_n_4505), .o(g64778_sb) );
na02s01 TIMEBOOST_cell_38601 ( .a(TIMEBOOST_net_10912), .b(g58006_db), .o(n_9788) );
na02m02 TIMEBOOST_cell_68701 ( .a(TIMEBOOST_net_21558), .b(TIMEBOOST_net_14202), .o(TIMEBOOST_net_17450) );
na02s01 TIMEBOOST_cell_38591 ( .a(TIMEBOOST_net_10907), .b(g58074_db), .o(n_9086) );
in01m01 g64779_u0 ( .a(FE_OFN669_n_4505), .o(g64779_sb) );
na02s01 TIMEBOOST_cell_37313 ( .a(TIMEBOOST_net_10268), .b(FE_OFN1003_n_2047), .o(TIMEBOOST_net_8223) );
na02m02 TIMEBOOST_cell_39750 ( .a(g58395_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q), .o(TIMEBOOST_net_11487) );
in01m06 g64780_u0 ( .a(FE_OFN670_n_4505), .o(g64780_sb) );
na02m08 g64780_u2 ( .a(FE_OFN670_n_4505), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q), .o(g64780_db) );
na02s01 TIMEBOOST_cell_49491 ( .a(FE_OFN258_n_9862), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q), .o(TIMEBOOST_net_14963) );
in01m01 g64781_u0 ( .a(FE_OFN672_n_4505), .o(g64781_sb) );
na02f01 TIMEBOOST_cell_68829 ( .a(TIMEBOOST_net_21622), .b(n_4447), .o(TIMEBOOST_net_17380) );
na02m02 g64781_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q), .b(FE_OFN672_n_4505), .o(g64781_db) );
in01m08 g64782_u0 ( .a(FE_OFN672_n_4505), .o(g64782_sb) );
na02s01 TIMEBOOST_cell_45247 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q), .o(TIMEBOOST_net_13518) );
in01m02 g64783_u0 ( .a(FE_OFN669_n_4505), .o(g64783_sb) );
na03f04 TIMEBOOST_cell_70860 ( .a(wbm_adr_o_12_), .b(g62068_sb), .c(g52441_sb), .o(TIMEBOOST_net_22638) );
na03m02 TIMEBOOST_cell_66097 ( .a(pci_target_unit_wishbone_master_bc_register_reg_2__Q), .b(g52592_sb), .c(TIMEBOOST_net_5511), .o(n_14685) );
in01m02 g64784_u0 ( .a(FE_OFN1660_n_4490), .o(g64784_sb) );
na02m02 TIMEBOOST_cell_48791 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q), .b(g58304_sb), .o(TIMEBOOST_net_14613) );
na03f02 TIMEBOOST_cell_34760 ( .a(TIMEBOOST_net_9468), .b(FE_OFN1409_n_8567), .c(g57513_sb), .o(n_11229) );
in01m02 g64785_u0 ( .a(FE_OFN669_n_4505), .o(g64785_sb) );
na02s01 TIMEBOOST_cell_62976 ( .a(conf_wb_err_addr_in_945), .b(configuration_wb_err_addr_536), .o(TIMEBOOST_net_20435) );
na03m06 TIMEBOOST_cell_68802 ( .a(TIMEBOOST_net_17213), .b(FE_OFN918_n_4725), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q), .o(TIMEBOOST_net_21609) );
in01f01 g64786_u0 ( .a(FE_OFN1659_n_4490), .o(g64786_sb) );
na02m01 g64786_u2 ( .a(n_3763), .b(FE_OFN1659_n_4490), .o(g64786_db) );
na03f02 TIMEBOOST_cell_73665 ( .a(TIMEBOOST_net_21063), .b(FE_OFN1135_g64577_p), .c(g62856_sb), .o(n_5255) );
in01m02 g64787_u0 ( .a(FE_OFN671_n_4505), .o(g64787_sb) );
na02m02 TIMEBOOST_cell_53456 ( .a(TIMEBOOST_net_16945), .b(FE_OFN1074_n_4740), .o(TIMEBOOST_net_14880) );
in01m01 g64788_u0 ( .a(FE_OFN667_n_4495), .o(g64788_sb) );
na02f02 TIMEBOOST_cell_69206 ( .a(TIMEBOOST_net_14192), .b(n_6136), .o(TIMEBOOST_net_21811) );
na03f02 TIMEBOOST_cell_66600 ( .a(TIMEBOOST_net_17094), .b(FE_OFN1310_n_6624), .c(g62898_sb), .o(n_6081) );
na02f02 TIMEBOOST_cell_51576 ( .a(TIMEBOOST_net_16005), .b(n_10134), .o(n_12156) );
in01m01 g64789_u0 ( .a(FE_OFN666_n_4495), .o(g64789_sb) );
na03m02 TIMEBOOST_cell_73175 ( .a(g64308_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q), .c(TIMEBOOST_net_14752), .o(TIMEBOOST_net_8332) );
na02m02 TIMEBOOST_cell_53090 ( .a(TIMEBOOST_net_16762), .b(TIMEBOOST_net_13022), .o(TIMEBOOST_net_9563) );
in01m02 g64790_u0 ( .a(FE_OFN669_n_4505), .o(g64790_sb) );
na02f02 TIMEBOOST_cell_70853 ( .a(TIMEBOOST_net_22634), .b(g62034_sb), .o(n_7782) );
na02m08 TIMEBOOST_cell_43029 ( .a(pci_target_unit_fifos_pciw_addr_data_in_149), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q), .o(TIMEBOOST_net_12409) );
in01m01 g64791_u0 ( .a(FE_OFN667_n_4495), .o(g64791_sb) );
na03m02 TIMEBOOST_cell_68942 ( .a(g64934_sb), .b(n_4442), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q), .o(TIMEBOOST_net_21679) );
in01m01 g64792_u0 ( .a(FE_OFN667_n_4495), .o(g64792_sb) );
na03f02 TIMEBOOST_cell_73465 ( .a(TIMEBOOST_net_23332), .b(FE_OFN1223_n_6391), .c(g62634_sb), .o(n_6284) );
na02f02 TIMEBOOST_cell_68071 ( .a(TIMEBOOST_net_21243), .b(n_2237), .o(n_1372) );
in01m01 g64793_u0 ( .a(FE_OFN667_n_4495), .o(g64793_sb) );
na02s02 TIMEBOOST_cell_38527 ( .a(TIMEBOOST_net_10875), .b(g58204_db), .o(n_9583) );
na02s02 TIMEBOOST_cell_38525 ( .a(TIMEBOOST_net_10874), .b(g58000_db), .o(n_9793) );
in01m02 g64794_u0 ( .a(FE_OFN665_n_4495), .o(g64794_sb) );
na02f01 TIMEBOOST_cell_69056 ( .a(FE_OFN651_n_4508), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q), .o(TIMEBOOST_net_21736) );
in01m01 g64795_u0 ( .a(FE_OFN666_n_4495), .o(g64795_sb) );
na02m02 TIMEBOOST_cell_52426 ( .a(TIMEBOOST_net_16430), .b(g58302_sb), .o(n_9028) );
na02m01 g64795_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q), .b(FE_OFN666_n_4495), .o(g64795_db) );
na02s01 TIMEBOOST_cell_38529 ( .a(TIMEBOOST_net_10876), .b(g58162_db), .o(n_9626) );
in01m02 g64796_u0 ( .a(FE_OFN618_n_4490), .o(g64796_sb) );
na03s02 TIMEBOOST_cell_46608 ( .a(TIMEBOOST_net_12831), .b(g63603_sb), .c(g63603_db), .o(n_7207) );
na03f02 TIMEBOOST_cell_73734 ( .a(TIMEBOOST_net_13628), .b(FE_OFN2209_n_11027), .c(n_12362), .o(n_16601) );
in01m02 g64797_u0 ( .a(FE_OFN671_n_4505), .o(g64797_sb) );
na02s01 TIMEBOOST_cell_39729 ( .a(TIMEBOOST_net_11476), .b(g57901_db), .o(n_9224) );
na02f02 TIMEBOOST_cell_49822 ( .a(TIMEBOOST_net_15128), .b(g63074_sb), .o(n_5102) );
in01m02 g64798_u0 ( .a(FE_OFN664_n_4495), .o(g64798_sb) );
na02m02 TIMEBOOST_cell_47905 ( .a(pci_target_unit_fifos_pciw_cbe_in_152), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q), .o(TIMEBOOST_net_14170) );
na04f04 TIMEBOOST_cell_73262 ( .a(n_1571), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q), .c(FE_OFN2212_n_8407), .d(g61941_sb), .o(n_7941) );
in01m02 g64799_u0 ( .a(FE_OFN664_n_4495), .o(g64799_sb) );
na02s01 TIMEBOOST_cell_52728 ( .a(TIMEBOOST_net_16581), .b(FE_OFN237_n_9118), .o(TIMEBOOST_net_9526) );
no04f06 TIMEBOOST_cell_68036 ( .a(TIMEBOOST_net_463), .b(FE_RN_573_0), .c(TIMEBOOST_net_8835), .d(FE_RN_562_0), .o(FE_RN_577_0) );
in01m01 g64800_u0 ( .a(FE_OFN1663_n_4490), .o(g64800_sb) );
na02m04 TIMEBOOST_cell_69388 ( .a(FE_OFN647_n_4497), .b(n_4429), .o(TIMEBOOST_net_21902) );
na03f02 TIMEBOOST_cell_34762 ( .a(TIMEBOOST_net_9361), .b(FE_OFN1370_n_8567), .c(g57086_sb), .o(n_10491) );
na02m03 TIMEBOOST_cell_72149 ( .a(TIMEBOOST_net_23282), .b(g64247_sb), .o(n_3925) );
in01m01 g64801_u0 ( .a(FE_OFN664_n_4495), .o(g64801_sb) );
no03f02 TIMEBOOST_cell_47341 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(TIMEBOOST_net_13635), .c(FE_RN_729_0), .o(n_12636) );
na02m01 g64801_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q), .b(FE_OFN664_n_4495), .o(g64801_db) );
in01m02 g64802_u0 ( .a(FE_OFN664_n_4495), .o(g64802_sb) );
na02s01 TIMEBOOST_cell_45807 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q), .o(TIMEBOOST_net_13798) );
in01m02 g64803_u0 ( .a(FE_OFN671_n_4505), .o(g64803_sb) );
na02m02 g64803_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q), .b(FE_OFN671_n_4505), .o(g64803_db) );
na03m02 TIMEBOOST_cell_69656 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q), .b(TIMEBOOST_net_7039), .c(g65817_db), .o(TIMEBOOST_net_22036) );
in01m04 g64804_u0 ( .a(FE_OFN669_n_4505), .o(g64804_sb) );
na02m02 TIMEBOOST_cell_18075 ( .a(n_272), .b(FE_OCP_RBN1917_wbs_cti_i_1_), .o(TIMEBOOST_net_5401) );
in01s01 TIMEBOOST_cell_73849 ( .a(TIMEBOOST_net_23413), .o(TIMEBOOST_net_23414) );
in01m01 g64805_u0 ( .a(FE_OFN649_n_4497), .o(g64805_sb) );
na03m02 TIMEBOOST_cell_70362 ( .a(FE_OFN2021_n_4778), .b(TIMEBOOST_net_16653), .c(TIMEBOOST_net_638), .o(TIMEBOOST_net_22389) );
na02s02 g65920_u2 ( .a(FE_OFN948_n_2248), .b(TIMEBOOST_net_20729), .o(g65920_db) );
in01m04 g64806_u0 ( .a(FE_OFN670_n_4505), .o(g64806_sb) );
na02s01 TIMEBOOST_cell_63254 ( .a(g58433_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q), .o(TIMEBOOST_net_20574) );
na02f01 TIMEBOOST_cell_43411 ( .a(n_3764), .b(g64786_sb), .o(TIMEBOOST_net_12600) );
in01m04 g64807_u0 ( .a(FE_OFN614_n_4501), .o(g64807_sb) );
na02f04 TIMEBOOST_cell_70196 ( .a(TIMEBOOST_net_14903), .b(g54305_sb), .o(TIMEBOOST_net_22306) );
na02m10 TIMEBOOST_cell_52449 ( .a(configuration_pci_err_addr_483), .b(wbm_adr_o_13_), .o(TIMEBOOST_net_16442) );
in01m02 g64808_u0 ( .a(FE_OFN664_n_4495), .o(g64808_sb) );
na02s01 TIMEBOOST_cell_42985 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q), .o(TIMEBOOST_net_12387) );
na02m01 TIMEBOOST_cell_64108 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q), .b(n_13544), .o(TIMEBOOST_net_21040) );
in01m02 g64809_u0 ( .a(FE_OFN672_n_4505), .o(g64809_sb) );
na02s01 TIMEBOOST_cell_42877 ( .a(pci_target_unit_fifos_pcir_control_in_192), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q), .o(TIMEBOOST_net_12333) );
na02s02 TIMEBOOST_cell_39760 ( .a(FE_OFN245_n_9114), .b(g57941_sb), .o(TIMEBOOST_net_11492) );
in01s01 g64810_u0 ( .a(n_4460), .o(g64810_sb) );
na02s02 TIMEBOOST_cell_71416 ( .a(g58001_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_22916) );
na02m01 g64810_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q), .b(n_4460), .o(g64810_db) );
na03s02 TIMEBOOST_cell_278 ( .a(n_1709), .b(g61746_sb), .c(g61922_db), .o(n_7977) );
in01m04 g64811_u0 ( .a(FE_OFN681_n_4460), .o(g64811_sb) );
na03f04 TIMEBOOST_cell_70308 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_410), .b(g54145_sb), .c(n_2105), .o(TIMEBOOST_net_22362) );
na02m02 TIMEBOOST_cell_50512 ( .a(TIMEBOOST_net_15473), .b(g62538_sb), .o(n_6493) );
na03s02 TIMEBOOST_cell_41701 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q), .b(g58404_sb), .c(g58404_db), .o(n_9003) );
in01m01 g64812_u0 ( .a(FE_OFN681_n_4460), .o(g64812_sb) );
na03m02 TIMEBOOST_cell_73140 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(g64116_sb), .c(g64116_db), .o(n_4044) );
na02s01 TIMEBOOST_cell_43037 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q), .o(TIMEBOOST_net_12413) );
in01s01 TIMEBOOST_cell_73965 ( .a(TIMEBOOST_net_23529), .o(TIMEBOOST_net_23530) );
in01m01 g64813_u0 ( .a(n_4460), .o(g64813_sb) );
na02s01 TIMEBOOST_cell_49492 ( .a(TIMEBOOST_net_14963), .b(FE_OFN572_n_9502), .o(TIMEBOOST_net_11198) );
no02f02 TIMEBOOST_cell_45412 ( .a(TIMEBOOST_net_13600), .b(n_7709), .o(n_13566) );
na02m02 TIMEBOOST_cell_69112 ( .a(n_4312), .b(FE_OFN618_n_4490), .o(TIMEBOOST_net_21764) );
in01m01 g64814_u0 ( .a(n_4460), .o(g64814_sb) );
na02s01 TIMEBOOST_cell_38803 ( .a(TIMEBOOST_net_11013), .b(g65858_sb), .o(n_2482) );
na02m01 g64814_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q), .b(n_4460), .o(g64814_db) );
na02m01 TIMEBOOST_cell_42814 ( .a(TIMEBOOST_net_12301), .b(g65835_sb), .o(TIMEBOOST_net_8781) );
in01m01 g64815_u0 ( .a(n_4460), .o(g64815_sb) );
na02m01 g64815_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q), .b(n_4460), .o(g64815_db) );
na02m08 TIMEBOOST_cell_69408 ( .a(pci_target_unit_fifos_pciw_addr_data_in), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q), .o(TIMEBOOST_net_21912) );
in01m02 g64816_u0 ( .a(FE_OFN682_n_4460), .o(g64816_sb) );
na02f02 TIMEBOOST_cell_71319 ( .a(TIMEBOOST_net_22867), .b(TIMEBOOST_net_21049), .o(TIMEBOOST_net_9524) );
na02m02 g64816_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q), .b(n_4460), .o(g64816_db) );
na03f02 TIMEBOOST_cell_73418 ( .a(TIMEBOOST_net_20519), .b(FE_OFN1212_n_4151), .c(g62913_sb), .o(n_6053) );
in01m04 g64817_u0 ( .a(FE_OFN681_n_4460), .o(g64817_sb) );
na02m02 TIMEBOOST_cell_71524 ( .a(TIMEBOOST_net_13538), .b(FE_OCPN1825_n_12030), .o(TIMEBOOST_net_22970) );
na02s01 TIMEBOOST_cell_69158 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q), .b(g65952_sb), .o(TIMEBOOST_net_21787) );
na04f04 TIMEBOOST_cell_36830 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q), .b(FE_OFN1404_n_8567), .c(n_9068), .d(g57290_sb), .o(n_10411) );
in01m01 g64818_u0 ( .a(FE_OFN682_n_4460), .o(g64818_sb) );
na02s01 TIMEBOOST_cell_43077 ( .a(FE_OFN243_n_9116), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q), .o(TIMEBOOST_net_12433) );
in01f01 g64819_u0 ( .a(FE_OFN623_n_4409), .o(g64819_sb) );
na02f01 TIMEBOOST_cell_69172 ( .a(g64286_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q), .o(TIMEBOOST_net_21794) );
na02f01 g64819_u2 ( .a(n_3738), .b(FE_OFN623_n_4409), .o(g64819_db) );
na02m01 TIMEBOOST_cell_53061 ( .a(configuration_pci_err_addr_501), .b(wbm_adr_o_31_), .o(TIMEBOOST_net_16748) );
in01m04 g64820_u0 ( .a(FE_OFN682_n_4460), .o(g64820_sb) );
na04m02 TIMEBOOST_cell_67251 ( .a(n_3749), .b(g64907_sb), .c(g64907_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q), .o(TIMEBOOST_net_17099) );
na02s01 TIMEBOOST_cell_43069 ( .a(FE_OFN243_n_9116), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q), .o(TIMEBOOST_net_12429) );
na02s02 TIMEBOOST_cell_63055 ( .a(TIMEBOOST_net_20474), .b(g58214_sb), .o(n_9563) );
in01m01 g64821_u0 ( .a(n_4460), .o(g64821_sb) );
na04f04 TIMEBOOST_cell_73263 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q), .b(FE_OFN2212_n_8407), .c(n_1598), .d(g61822_sb), .o(n_8144) );
na02s01 TIMEBOOST_cell_30979 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_3__Q), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9594) );
na02f02 TIMEBOOST_cell_18331 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_5529) );
in01m04 g64822_u0 ( .a(FE_OFN682_n_4460), .o(g64822_sb) );
na02m06 g64822_u2 ( .a(FE_OFN682_n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q), .o(g64822_db) );
na04s02 TIMEBOOST_cell_72884 ( .a(g61749_sb), .b(g61749_db), .c(g65763_db), .d(g65763_da), .o(n_8319) );
in01m01 g64823_u0 ( .a(FE_OFN682_n_4460), .o(g64823_sb) );
na02m10 TIMEBOOST_cell_45709 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_13749) );
na02m02 TIMEBOOST_cell_68117 ( .a(TIMEBOOST_net_21266), .b(g54219_sb), .o(TIMEBOOST_net_12277) );
na02f02 TIMEBOOST_cell_53309 ( .a(n_17044), .b(n_10069), .o(TIMEBOOST_net_16872) );
in01m01 g64824_u0 ( .a(FE_OFN679_n_4460), .o(g64824_sb) );
na03f02 TIMEBOOST_cell_72712 ( .a(g65074_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q), .c(TIMEBOOST_net_10603), .o(TIMEBOOST_net_17571) );
na02s02 TIMEBOOST_cell_43085 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q), .o(TIMEBOOST_net_12437) );
na02m02 TIMEBOOST_cell_68683 ( .a(TIMEBOOST_net_21549), .b(g64330_db), .o(n_3846) );
in01m01 g64825_u0 ( .a(FE_OFN679_n_4460), .o(g64825_sb) );
in01m02 g64826_u0 ( .a(FE_OFN629_n_4454), .o(g64826_sb) );
in01s01 TIMEBOOST_cell_72350 ( .a(pci_target_unit_fifos_pcir_data_in_161), .o(TIMEBOOST_net_23383) );
na02s01 TIMEBOOST_cell_38499 ( .a(TIMEBOOST_net_10861), .b(g57970_db), .o(n_9831) );
in01m01 g64827_u0 ( .a(FE_OFN1810_n_4454), .o(g64827_sb) );
na03m04 TIMEBOOST_cell_72652 ( .a(TIMEBOOST_net_21494), .b(g65034_sb), .c(TIMEBOOST_net_21676), .o(TIMEBOOST_net_17048) );
na02f01 TIMEBOOST_cell_71650 ( .a(FE_OFN1761_n_10780), .b(TIMEBOOST_net_13520), .o(TIMEBOOST_net_23033) );
in01m02 g64828_u0 ( .a(FE_OFN631_n_4454), .o(g64828_sb) );
in01m01 g64829_u0 ( .a(FE_OFN634_n_4454), .o(g64829_sb) );
in01s01 TIMEBOOST_cell_63576 ( .a(TIMEBOOST_net_20756), .o(wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_Q) );
na04f02 TIMEBOOST_cell_35119 ( .a(wbs_dat_o_22_), .b(g52517_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_121), .d(FE_OFN1472_g52675_p), .o(n_13798) );
in01m04 g64830_u0 ( .a(FE_OFN631_n_4454), .o(g64830_sb) );
na02m01 TIMEBOOST_cell_42730 ( .a(TIMEBOOST_net_12259), .b(wbu_addr_in_253), .o(TIMEBOOST_net_10150) );
in01m01 g64831_u0 ( .a(FE_OFN1810_n_4454), .o(g64831_sb) );
na03f02 TIMEBOOST_cell_34906 ( .a(TIMEBOOST_net_9485), .b(FE_OFN1380_n_8567), .c(g57156_sb), .o(n_10462) );
in01m02 g64832_u0 ( .a(FE_OFN1810_n_4454), .o(g64832_sb) );
na03f02 TIMEBOOST_cell_34908 ( .a(TIMEBOOST_net_9486), .b(FE_OFN1383_n_8567), .c(g57326_sb), .o(n_11424) );
na03m02 TIMEBOOST_cell_65431 ( .a(TIMEBOOST_net_16245), .b(g64837_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q), .o(TIMEBOOST_net_17552) );
na02m04 TIMEBOOST_cell_69424 ( .a(FE_OFN646_n_4497), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q), .o(TIMEBOOST_net_21920) );
in01m02 g64833_u0 ( .a(FE_OFN633_n_4454), .o(g64833_sb) );
na02m02 g64833_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q), .b(FE_OFN633_n_4454), .o(g64833_db) );
na03m02 TIMEBOOST_cell_68874 ( .a(g64932_sb), .b(n_4493), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q), .o(TIMEBOOST_net_21645) );
in01m01 g64834_u0 ( .a(FE_OFN1809_n_4454), .o(g64834_sb) );
na02m02 TIMEBOOST_cell_51943 ( .a(FE_OFN905_n_4736), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q), .o(TIMEBOOST_net_16189) );
na02m02 TIMEBOOST_cell_68169 ( .a(TIMEBOOST_net_21292), .b(TIMEBOOST_net_12277), .o(TIMEBOOST_net_16806) );
in01s01 TIMEBOOST_cell_63593 ( .a(TIMEBOOST_net_20773), .o(TIMEBOOST_net_20772) );
in01m01 g64835_u0 ( .a(FE_OFN1809_n_4454), .o(g64835_sb) );
na02s04 TIMEBOOST_cell_68128 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_89), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_21272) );
na02f01 g64835_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q), .b(FE_OFN1809_n_4454), .o(g64835_db) );
na02s01 TIMEBOOST_cell_18007 ( .a(n_1816), .b(n_709), .o(TIMEBOOST_net_5367) );
in01m02 g64836_u0 ( .a(FE_OFN629_n_4454), .o(g64836_sb) );
na02s01 TIMEBOOST_cell_45809 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_13799) );
na02s02 TIMEBOOST_cell_38503 ( .a(TIMEBOOST_net_10863), .b(g58221_sb), .o(n_9565) );
in01m01 g64837_u0 ( .a(FE_OFN631_n_4454), .o(g64837_sb) );
na02m01 TIMEBOOST_cell_52363 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(FE_OFN1032_n_4732), .o(TIMEBOOST_net_16399) );
in01m01 g64838_u0 ( .a(FE_OFN631_n_4454), .o(g64838_sb) );
na02s02 TIMEBOOST_cell_38541 ( .a(TIMEBOOST_net_10882), .b(n_8892), .o(n_9435) );
na02m04 TIMEBOOST_cell_72012 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q), .b(g65871_sb), .o(TIMEBOOST_net_23214) );
in01m01 g64839_u0 ( .a(FE_OFN634_n_4454), .o(g64839_sb) );
na03f02 TIMEBOOST_cell_69482 ( .a(TIMEBOOST_net_21175), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q), .c(g65965_sb), .o(TIMEBOOST_net_21949) );
na02s01 TIMEBOOST_cell_38501 ( .a(TIMEBOOST_net_10862), .b(g58228_db), .o(n_9561) );
in01m02 g64840_u0 ( .a(FE_OFN628_n_4454), .o(g64840_sb) );
na02s01 TIMEBOOST_cell_39764 ( .a(FE_OFN245_n_9114), .b(g57973_sb), .o(TIMEBOOST_net_11494) );
in01s01 TIMEBOOST_cell_73898 ( .a(n_8144), .o(TIMEBOOST_net_23463) );
in01s02 TIMEBOOST_cell_45935 ( .a(TIMEBOOST_net_13896), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_86) );
in01m02 g64841_u0 ( .a(FE_OFN630_n_4454), .o(g64841_sb) );
na02m01 TIMEBOOST_cell_68442 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q), .b(FE_OFN669_n_4505), .o(TIMEBOOST_net_21429) );
na03s02 TIMEBOOST_cell_72909 ( .a(n_1569), .b(g61931_sb), .c(g61931_db), .o(n_7961) );
na02m02 TIMEBOOST_cell_37688 ( .a(FE_OFN1624_n_4438), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_10456) );
in01m01 g64842_u0 ( .a(FE_OFN689_n_4438), .o(g64842_sb) );
in01m01 g64843_u0 ( .a(FE_OFN1625_n_4438), .o(g64843_sb) );
na04f04 TIMEBOOST_cell_36856 ( .a(n_2925), .b(n_2858), .c(n_3068), .d(n_2870), .o(n_4172) );
na02m01 g64843_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q), .b(FE_OFN1625_n_4438), .o(g64843_db) );
na04f02 TIMEBOOST_cell_36858 ( .a(g52619_sb), .b(n_10256), .c(TIMEBOOST_net_9585), .d(TIMEBOOST_net_767), .o(n_11851) );
in01m02 g64844_u0 ( .a(FE_OFN1624_n_4438), .o(g64844_sb) );
na03f02 TIMEBOOST_cell_73524 ( .a(TIMEBOOST_net_17062), .b(n_6645), .c(g62435_sb), .o(n_6726) );
in01s01 TIMEBOOST_cell_63608 ( .a(TIMEBOOST_net_20788), .o(TIMEBOOST_net_20725) );
in01m02 g64845_u0 ( .a(FE_OFN1625_n_4438), .o(g64845_sb) );
na02s01 TIMEBOOST_cell_43129 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q), .o(TIMEBOOST_net_12459) );
in01m01 g64846_u0 ( .a(FE_OFN1624_n_4438), .o(g64846_sb) );
na02s01 TIMEBOOST_cell_43035 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_130), .o(TIMEBOOST_net_12412) );
in01s01 TIMEBOOST_cell_67723 ( .a(pci_target_unit_fifos_pcir_data_in_172), .o(TIMEBOOST_net_21150) );
in01m01 g64847_u0 ( .a(FE_OFN1625_n_4438), .o(g64847_sb) );
na02s02 TIMEBOOST_cell_43111 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q), .b(pci_target_unit_fifos_pcir_data_in_160), .o(TIMEBOOST_net_12450) );
na02s08 TIMEBOOST_cell_72090 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q), .b(pci_target_unit_fifos_pciw_control_in_156), .o(TIMEBOOST_net_23253) );
in01m01 g64848_u0 ( .a(FE_OFN1625_n_4438), .o(g64848_sb) );
na02m10 TIMEBOOST_cell_52659 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q), .o(TIMEBOOST_net_16547) );
na02s02 TIMEBOOST_cell_43073 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_12431) );
na02s01 TIMEBOOST_cell_31017 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_1__Q), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_9613) );
in01m02 g64849_u0 ( .a(FE_OFN1626_n_4438), .o(g64849_sb) );
na02m02 g64849_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q), .b(FE_OFN1626_n_4438), .o(g64849_db) );
na02m01 TIMEBOOST_cell_62953 ( .a(TIMEBOOST_net_20423), .b(g57923_db), .o(n_9887) );
in01m02 g64850_u0 ( .a(FE_OFN1628_n_4438), .o(g64850_sb) );
na03f02 TIMEBOOST_cell_73419 ( .a(TIMEBOOST_net_20971), .b(FE_OFN1208_n_6356), .c(g62682_sb), .o(n_6175) );
na04f06 TIMEBOOST_cell_68016 ( .a(TIMEBOOST_net_16779), .b(g54183_sb), .c(wishbone_slave_unit_del_sync_addr_out_reg_20__Q), .d(FE_OFN1084_n_13221), .o(n_13430) );
na02m04 TIMEBOOST_cell_68864 ( .a(n_4444), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q), .o(TIMEBOOST_net_21640) );
in01m01 g64851_u0 ( .a(FE_OFN1624_n_4438), .o(g64851_sb) );
na02f01 TIMEBOOST_cell_44410 ( .a(TIMEBOOST_net_13099), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_11443) );
na02s01 TIMEBOOST_cell_43109 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q), .b(FE_OFN535_n_9823), .o(TIMEBOOST_net_12449) );
in01m01 g64852_u0 ( .a(FE_OFN1625_n_4438), .o(g64852_sb) );
na02s04 TIMEBOOST_cell_71150 ( .a(FE_OFN241_n_9830), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q), .o(TIMEBOOST_net_22783) );
na02s02 TIMEBOOST_cell_64029 ( .a(TIMEBOOST_net_21000), .b(FE_OFN241_n_9830), .o(n_9729) );
in01m04 g64853_u0 ( .a(FE_OFN1626_n_4438), .o(g64853_sb) );
na02s01 TIMEBOOST_cell_43107 ( .a(pci_target_unit_fifos_pcir_data_in), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q), .o(TIMEBOOST_net_12448) );
na04m04 TIMEBOOST_cell_67232 ( .a(g64783_sb), .b(n_3764), .c(g64783_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q), .o(TIMEBOOST_net_17492) );
in01m01 g64854_u0 ( .a(FE_OFN1626_n_4438), .o(g64854_sb) );
in01s01 TIMEBOOST_cell_67725 ( .a(pci_target_unit_fifos_pcir_data_in_178), .o(TIMEBOOST_net_21152) );
na03f02 TIMEBOOST_cell_70706 ( .a(n_4611), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q), .c(FE_OFN1118_g64577_p), .o(TIMEBOOST_net_22561) );
na04f02 TIMEBOOST_cell_73466 ( .a(n_4402), .b(FE_OFN1223_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q), .d(g62605_sb), .o(n_6342) );
in01m06 g64855_u0 ( .a(FE_OFN1626_n_4438), .o(g64855_sb) );
na04f02 TIMEBOOST_cell_72477 ( .a(TIMEBOOST_net_21352), .b(g64114_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q), .d(FE_OFN717_n_8176), .o(TIMEBOOST_net_22580) );
na03f02 TIMEBOOST_cell_73756 ( .a(n_13901), .b(TIMEBOOST_net_13696), .c(FE_OFN1593_n_13741), .o(g53263_p) );
in01m01 g64856_u0 ( .a(FE_OFN689_n_4438), .o(g64856_sb) );
na04s04 TIMEBOOST_cell_46496 ( .a(TIMEBOOST_net_12722), .b(FE_OFN1802_n_9690), .c(g58242_sb), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q), .o(TIMEBOOST_net_9424) );
na02m08 TIMEBOOST_cell_45463 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q), .o(TIMEBOOST_net_13626) );
in01m02 g64857_u0 ( .a(FE_OFN1623_n_4438), .o(g64857_sb) );
na03m04 TIMEBOOST_cell_72929 ( .a(g65277_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q), .c(TIMEBOOST_net_12641), .o(TIMEBOOST_net_17159) );
in01m01 g64858_u0 ( .a(FE_OFN615_n_4501), .o(g64858_sb) );
na03f02 TIMEBOOST_cell_34764 ( .a(TIMEBOOST_net_9348), .b(FE_OFN1397_n_8567), .c(g57241_sb), .o(n_11517) );
na02s02 TIMEBOOST_cell_44141 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_12965) );
in01m01 g64859_u0 ( .a(FE_OFN612_n_4501), .o(g64859_sb) );
na03f02 TIMEBOOST_cell_66789 ( .a(TIMEBOOST_net_17012), .b(FE_OFN1272_n_4096), .c(g63002_sb), .o(n_5878) );
na03f02 TIMEBOOST_cell_34766 ( .a(TIMEBOOST_net_9357), .b(FE_OFN1368_n_8567), .c(g57321_sb), .o(n_11429) );
na03f02 TIMEBOOST_cell_73639 ( .a(TIMEBOOST_net_17547), .b(FE_OFN1253_n_4143), .c(g62413_sb), .o(n_6772) );
in01m04 g64860_u0 ( .a(FE_OFN647_n_4497), .o(g64860_sb) );
na02s01 TIMEBOOST_cell_49291 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q), .b(FE_OFN519_n_9697), .o(TIMEBOOST_net_14863) );
na02m10 TIMEBOOST_cell_45609 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q), .o(TIMEBOOST_net_13699) );
in01m01 g64861_u0 ( .a(FE_OFN1663_n_4490), .o(g64861_sb) );
na02f02 TIMEBOOST_cell_40040 ( .a(wbm_adr_o_13_), .b(g59387_sb), .o(TIMEBOOST_net_11632) );
in01m02 g64862_u0 ( .a(FE_OFN615_n_4501), .o(g64862_sb) );
na03f02 TIMEBOOST_cell_73420 ( .a(TIMEBOOST_net_20585), .b(FE_OFN1207_n_6356), .c(g62597_sb), .o(n_6358) );
na03s02 TIMEBOOST_cell_46610 ( .a(TIMEBOOST_net_12838), .b(g63607_sb), .c(g63607_db), .o(n_7151) );
in01m04 g64863_u0 ( .a(FE_OFN615_n_4501), .o(g64863_sb) );
na03f02 TIMEBOOST_cell_34768 ( .a(TIMEBOOST_net_9350), .b(FE_OFN1383_n_8567), .c(g57426_sb), .o(n_11309) );
in01f01 g64864_u0 ( .a(FE_OFN1807_n_4501), .o(g64864_sb) );
na02m10 TIMEBOOST_cell_41066 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q), .o(TIMEBOOST_net_12145) );
na02m01 g64864_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q), .b(FE_OFN1807_n_4501), .o(g64864_db) );
na02s01 TIMEBOOST_cell_71156 ( .a(TIMEBOOST_net_12799), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q), .o(TIMEBOOST_net_22786) );
in01m04 g64865_u0 ( .a(FE_OFN615_n_4501), .o(g64865_sb) );
na03f02 TIMEBOOST_cell_34770 ( .a(TIMEBOOST_net_9351), .b(FE_OFN1409_n_8567), .c(g57147_sb), .o(n_11603) );
na02m02 TIMEBOOST_cell_63369 ( .a(TIMEBOOST_net_20631), .b(TIMEBOOST_net_12970), .o(TIMEBOOST_net_9405) );
in01m04 g64866_u0 ( .a(FE_OFN612_n_4501), .o(g64866_sb) );
na02m02 TIMEBOOST_cell_70237 ( .a(TIMEBOOST_net_22326), .b(FE_OFN720_n_8060), .o(TIMEBOOST_net_15035) );
na03m02 TIMEBOOST_cell_70110 ( .a(n_4476), .b(g64972_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q), .o(TIMEBOOST_net_22263) );
na03m02 TIMEBOOST_cell_69748 ( .a(n_4473), .b(FE_OFN1642_n_4671), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q), .o(TIMEBOOST_net_22082) );
in01m04 g64867_u0 ( .a(FE_OFN1807_n_4501), .o(g64867_sb) );
na02m02 TIMEBOOST_cell_69544 ( .a(g64921_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q), .o(TIMEBOOST_net_21980) );
na02s01 TIMEBOOST_cell_45413 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q), .o(TIMEBOOST_net_13601) );
in01m04 g64868_u0 ( .a(FE_OFN615_n_4501), .o(g64868_sb) );
na03f02 TIMEBOOST_cell_34772 ( .a(TIMEBOOST_net_9352), .b(FE_OFN1390_n_8567), .c(g57382_sb), .o(n_11363) );
na02s01 TIMEBOOST_cell_63124 ( .a(FE_OFN203_n_9228), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q), .o(TIMEBOOST_net_20509) );
in01m01 g64869_u0 ( .a(FE_OFN1806_n_4501), .o(g64869_sb) );
na03m02 TIMEBOOST_cell_72503 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q), .b(FE_OFN671_n_4505), .c(TIMEBOOST_net_21669), .o(TIMEBOOST_net_17428) );
na03f02 TIMEBOOST_cell_73640 ( .a(TIMEBOOST_net_17438), .b(FE_OFN1284_n_4097), .c(g62384_sb), .o(n_6833) );
in01m01 g64870_u0 ( .a(FE_OFN1807_n_4501), .o(g64870_sb) );
na03m02 TIMEBOOST_cell_70364 ( .a(FE_OFN2021_n_4778), .b(TIMEBOOST_net_16651), .c(TIMEBOOST_net_631), .o(TIMEBOOST_net_22390) );
na02m01 TIMEBOOST_cell_69266 ( .a(n_4444), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q), .o(TIMEBOOST_net_21841) );
na03s01 TIMEBOOST_cell_72569 ( .a(pci_target_unit_del_sync_addr_in_222), .b(g66403_sb), .c(g66409_db), .o(n_2528) );
in01m01 g64871_u0 ( .a(FE_OFN612_n_4501), .o(g64871_sb) );
na02f02 TIMEBOOST_cell_30944 ( .a(TIMEBOOST_net_9576), .b(n_2852), .o(n_4649) );
in01m01 g64872_u0 ( .a(FE_OFN615_n_4501), .o(g64872_sb) );
na02m01 TIMEBOOST_cell_52813 ( .a(n_1117), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .o(TIMEBOOST_net_16624) );
na02f04 TIMEBOOST_cell_62811 ( .a(TIMEBOOST_net_20352), .b(n_2722), .o(n_2723) );
na03f02 TIMEBOOST_cell_73735 ( .a(FE_OFN2209_n_11027), .b(TIMEBOOST_net_8606), .c(n_12362), .o(n_16592) );
in01m01 g64873_u0 ( .a(FE_OFN1807_n_4501), .o(g64873_sb) );
na02f01 TIMEBOOST_cell_62807 ( .a(TIMEBOOST_net_20350), .b(FE_OFN1059_n_4727), .o(TIMEBOOST_net_14703) );
na03s01 TIMEBOOST_cell_64737 ( .a(pci_target_unit_del_sync_addr_in_214), .b(g66406_sb), .c(g66416_db), .o(n_2517) );
in01m01 g64874_u0 ( .a(FE_OFN614_n_4501), .o(g64874_sb) );
na02m02 g64874_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q), .b(FE_OFN614_n_4501), .o(g64874_db) );
in01m01 g64875_u0 ( .a(FE_OFN664_n_4495), .o(g64875_sb) );
na02s01 TIMEBOOST_cell_47509 ( .a(parchk_pci_ad_reg_in_1225), .b(g67085_db), .o(TIMEBOOST_net_13972) );
na04f04 TIMEBOOST_cell_68017 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_406), .b(g54187_sb), .c(TIMEBOOST_net_7606), .d(FE_OFN1085_n_13221), .o(n_13428) );
na02m06 TIMEBOOST_cell_47541 ( .a(FE_OFN2115_wishbone_slave_unit_pci_initiator_if_data_source), .b(wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_13988) );
in01m01 g64876_u0 ( .a(FE_OFN612_n_4501), .o(g64876_sb) );
na02s01 TIMEBOOST_cell_30981 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_2__Q), .b(FE_OFN237_n_9118), .o(TIMEBOOST_net_9595) );
na03f02 TIMEBOOST_cell_73757 ( .a(TIMEBOOST_net_16058), .b(FE_OFN1774_n_13800), .c(FE_OFN1770_n_14054), .o(g53167_p) );
na02f02 TIMEBOOST_cell_70249 ( .a(TIMEBOOST_net_22332), .b(g61836_sb), .o(n_6975) );
in01m04 g64877_u0 ( .a(FE_OFN612_n_4501), .o(g64877_sb) );
na02s02 TIMEBOOST_cell_49274 ( .a(TIMEBOOST_net_14854), .b(TIMEBOOST_net_10857), .o(TIMEBOOST_net_9425) );
na02m01 TIMEBOOST_cell_69528 ( .a(n_4498), .b(n_95), .o(TIMEBOOST_net_21972) );
in01m01 g64878_u0 ( .a(FE_OFN665_n_4495), .o(g64878_sb) );
na02s02 TIMEBOOST_cell_48210 ( .a(TIMEBOOST_net_14322), .b(g57959_sb), .o(TIMEBOOST_net_10442) );
na03m06 TIMEBOOST_cell_64797 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q), .b(FE_OFN579_n_9531), .c(g58403_sb), .o(TIMEBOOST_net_14977) );
na02s01 TIMEBOOST_cell_48859 ( .a(FE_OFN239_n_9832), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q), .o(TIMEBOOST_net_14647) );
in01m04 g64879_u0 ( .a(FE_OFN686_n_4417), .o(g64879_sb) );
na02s01 TIMEBOOST_cell_52944 ( .a(TIMEBOOST_net_16689), .b(TIMEBOOST_net_12429), .o(TIMEBOOST_net_9516) );
no02f02 TIMEBOOST_cell_45131 ( .a(n_4144), .b(n_7552), .o(TIMEBOOST_net_13460) );
in01m04 g64880_u0 ( .a(FE_OFN686_n_4417), .o(g64880_sb) );
na02s01 TIMEBOOST_cell_31019 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_5__Q), .b(n_9114), .o(TIMEBOOST_net_9614) );
no02f02 TIMEBOOST_cell_45132 ( .a(TIMEBOOST_net_13460), .b(n_7214), .o(g59721_p) );
na02s02 TIMEBOOST_cell_48212 ( .a(TIMEBOOST_net_14323), .b(g58414_sb), .o(TIMEBOOST_net_9324) );
in01m02 g64881_u0 ( .a(FE_OFN685_n_4417), .o(g64881_sb) );
na02m02 TIMEBOOST_cell_69678 ( .a(g65354_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q), .o(TIMEBOOST_net_22047) );
in01m01 g64882_u0 ( .a(FE_OFN685_n_4417), .o(g64882_sb) );
na04f02 TIMEBOOST_cell_73447 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q), .b(n_4917), .c(FE_OFN1243_n_4092), .d(g62689_sb), .o(n_7366) );
na02m02 TIMEBOOST_cell_72247 ( .a(TIMEBOOST_net_23331), .b(g58288_sb), .o(TIMEBOOST_net_9557) );
in01m01 g64883_u0 ( .a(FE_OFN686_n_4417), .o(g64883_sb) );
na04f04 TIMEBOOST_cell_67511 ( .a(TIMEBOOST_net_16399), .b(TIMEBOOST_net_8767), .c(g63101_db), .d(g63101_sb), .o(n_5052) );
na02s01 TIMEBOOST_cell_31021 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_23__Q), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_9615) );
in01m01 g64884_u0 ( .a(FE_OFN686_n_4417), .o(g64884_sb) );
na02f10 TIMEBOOST_cell_68068 ( .a(n_193), .b(n_245), .o(TIMEBOOST_net_21242) );
na02s02 TIMEBOOST_cell_53070 ( .a(TIMEBOOST_net_16752), .b(FE_OFN584_n_9692), .o(TIMEBOOST_net_10872) );
in01m01 g64885_u0 ( .a(FE_OFN686_n_4417), .o(g64885_sb) );
na02s02 TIMEBOOST_cell_70493 ( .a(TIMEBOOST_net_22454), .b(g58029_sb), .o(n_9099) );
na02f02 TIMEBOOST_cell_45136 ( .a(TIMEBOOST_net_13462), .b(g63023_sb), .o(n_5200) );
na03f02 TIMEBOOST_cell_34737 ( .a(TIMEBOOST_net_9397), .b(FE_OFN1388_n_8567), .c(g57149_sb), .o(n_11601) );
in01m01 g64886_u0 ( .a(FE_OFN686_n_4417), .o(g64886_sb) );
na03f02 TIMEBOOST_cell_70392 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q), .b(FE_OFN720_n_8060), .c(n_1613), .o(TIMEBOOST_net_22404) );
na02m01 TIMEBOOST_cell_68302 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q), .b(n_4460), .o(TIMEBOOST_net_21359) );
in01m01 g64887_u0 ( .a(FE_OFN687_n_4417), .o(g64887_sb) );
na03f02 TIMEBOOST_cell_66234 ( .a(TIMEBOOST_net_20964), .b(FE_OFN1258_n_4143), .c(g62908_sb), .o(n_6061) );
na03m06 TIMEBOOST_cell_68288 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q), .b(FE_OFN937_n_2292), .c(pci_target_unit_fifos_pcir_control_in_192), .o(TIMEBOOST_net_21352) );
in01m02 g64888_u0 ( .a(FE_OFN685_n_4417), .o(g64888_sb) );
in01s01 TIMEBOOST_cell_67787 ( .a(TIMEBOOST_net_21214), .o(wbs_adr_i_23_) );
na02m02 g64888_u2 ( .a(FE_OFN685_n_4417), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q), .o(g64888_db) );
na03f02 TIMEBOOST_cell_72857 ( .a(g65406_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q), .c(TIMEBOOST_net_20843), .o(TIMEBOOST_net_17370) );
in01m01 g64889_u0 ( .a(FE_OFN685_n_4417), .o(g64889_sb) );
no02f02 TIMEBOOST_cell_51522 ( .a(TIMEBOOST_net_15978), .b(n_7091), .o(n_13568) );
in01m04 g64890_u0 ( .a(FE_OFN686_n_4417), .o(g64890_sb) );
na02s01 TIMEBOOST_cell_44025 ( .a(FE_OFN554_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q), .o(TIMEBOOST_net_12907) );
na02s01 TIMEBOOST_cell_47635 ( .a(g54219_sb), .b(TIMEBOOST_net_6805), .o(TIMEBOOST_net_14035) );
in01m02 g64891_u0 ( .a(FE_OFN687_n_4417), .o(g64891_sb) );
na03m02 TIMEBOOST_cell_70458 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q), .c(g58378_sb), .o(TIMEBOOST_net_22437) );
in01m02 g64892_u0 ( .a(FE_OFN687_n_4417), .o(g64892_sb) );
na03f02 TIMEBOOST_cell_34876 ( .a(TIMEBOOST_net_9467), .b(FE_OFN1407_n_8567), .c(g57517_sb), .o(n_11223) );
in01m01 g64893_u0 ( .a(FE_OFN686_n_4417), .o(g64893_sb) );
na02f10 TIMEBOOST_cell_43963 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_775), .o(TIMEBOOST_net_12876) );
na02m06 TIMEBOOST_cell_72336 ( .a(TIMEBOOST_net_15866), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_), .o(TIMEBOOST_net_23376) );
in01m02 g64894_u0 ( .a(FE_OFN687_n_4417), .o(g64894_sb) );
na03f02 TIMEBOOST_cell_73736 ( .a(FE_OFN1572_n_11027), .b(TIMEBOOST_net_8604), .c(n_12362), .o(n_16603) );
in01m02 g64895_u0 ( .a(FE_OFN687_n_4417), .o(g64895_sb) );
na03f02 TIMEBOOST_cell_73737 ( .a(FE_OFN1740_n_11019), .b(TIMEBOOST_net_8600), .c(FE_OFN1734_n_16317), .o(n_16589) );
in01s01 g64896_u0 ( .a(n_4417), .o(g64896_sb) );
na03s02 TIMEBOOST_cell_281 ( .a(n_1574), .b(g61894_sb), .c(g61928_db), .o(n_7967) );
na02s01 g64896_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q), .b(n_4417), .o(g64896_db) );
in01m02 g64897_u0 ( .a(FE_OFN684_n_4417), .o(g64897_sb) );
na02m02 TIMEBOOST_cell_68171 ( .a(TIMEBOOST_net_21293), .b(TIMEBOOST_net_16140), .o(TIMEBOOST_net_16793) );
na03f02 TIMEBOOST_cell_66596 ( .a(TIMEBOOST_net_17104), .b(FE_OFN1323_n_6436), .c(g62560_sb), .o(n_6440) );
na02m02 TIMEBOOST_cell_52714 ( .a(TIMEBOOST_net_16574), .b(FE_OFN917_n_4725), .o(TIMEBOOST_net_14301) );
in01m01 g64898_u0 ( .a(FE_OFN684_n_4417), .o(g64898_sb) );
na03m02 TIMEBOOST_cell_72479 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q), .b(FE_OFN1785_n_1699), .c(TIMEBOOST_net_21407), .o(n_4520) );
na02m01 TIMEBOOST_cell_52185 ( .a(configuration_wb_err_addr_562), .b(conf_wb_err_addr_in_971), .o(TIMEBOOST_net_16310) );
in01m01 g64899_u0 ( .a(FE_OFN624_n_4409), .o(g64899_sb) );
na02s01 TIMEBOOST_cell_39768 ( .a(g58034_sb), .b(FE_OFN245_n_9114), .o(TIMEBOOST_net_11496) );
na03f02 TIMEBOOST_cell_66810 ( .a(TIMEBOOST_net_16843), .b(FE_OFN1345_n_8567), .c(g57565_sb), .o(n_11187) );
na02s02 TIMEBOOST_cell_48642 ( .a(TIMEBOOST_net_14538), .b(TIMEBOOST_net_12734), .o(TIMEBOOST_net_9570) );
in01m01 g64900_u0 ( .a(FE_OFN624_n_4409), .o(g64900_sb) );
na02m02 TIMEBOOST_cell_68301 ( .a(TIMEBOOST_net_21358), .b(n_3749), .o(TIMEBOOST_net_16152) );
in01s06 TIMEBOOST_cell_67727 ( .a(TIMEBOOST_net_21154), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_90) );
in01m04 g64901_u0 ( .a(FE_OFN625_n_4409), .o(g64901_sb) );
na02f02 TIMEBOOST_cell_68411 ( .a(TIMEBOOST_net_21413), .b(n_1784), .o(TIMEBOOST_net_20880) );
na02m06 g64901_u2 ( .a(FE_OFN625_n_4409), .b(n_4410), .o(g64901_db) );
na03f02 TIMEBOOST_cell_34923 ( .a(TIMEBOOST_net_9472), .b(FE_OFN1404_n_8567), .c(g57070_sb), .o(n_11671) );
in01m01 g64902_u0 ( .a(FE_OFN625_n_4409), .o(g64902_sb) );
na02m02 TIMEBOOST_cell_68462 ( .a(FE_OFN672_n_4505), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q), .o(TIMEBOOST_net_21439) );
na02m01 TIMEBOOST_cell_42919 ( .a(FE_OFN622_n_4409), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q), .o(TIMEBOOST_net_12354) );
na02m02 TIMEBOOST_cell_69238 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q), .b(FE_OFN1676_n_4655), .o(TIMEBOOST_net_21827) );
in01m04 g64903_u0 ( .a(FE_OFN623_n_4409), .o(g64903_sb) );
na02s01 TIMEBOOST_cell_39770 ( .a(g58133_sb), .b(FE_OFN245_n_9114), .o(TIMEBOOST_net_11497) );
na02m04 g64903_u2 ( .a(n_3691), .b(FE_OFN623_n_4409), .o(g64903_db) );
in01f04 TIMEBOOST_cell_47507 ( .a(TIMEBOOST_net_13970), .o(n_13415) );
in01m01 g64904_u0 ( .a(FE_OFN623_n_4409), .o(g64904_sb) );
na03f04 TIMEBOOST_cell_47150 ( .a(TIMEBOOST_net_7603), .b(n_13625), .c(n_7695), .o(n_14485) );
na03f02 TIMEBOOST_cell_72807 ( .a(n_4493), .b(FE_OFN638_n_4669), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q), .o(TIMEBOOST_net_22019) );
na02s01 TIMEBOOST_cell_39797 ( .a(TIMEBOOST_net_11510), .b(g58439_db), .o(n_9200) );
in01m08 g64905_u0 ( .a(FE_OFN624_n_4409), .o(g64905_sb) );
na03f02 TIMEBOOST_cell_65665 ( .a(TIMEBOOST_net_16354), .b(g64217_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q), .o(TIMEBOOST_net_17322) );
in01m01 g64906_u0 ( .a(FE_OFN624_n_4409), .o(g64906_sb) );
na02f02 TIMEBOOST_cell_71743 ( .a(TIMEBOOST_net_23079), .b(FE_OCP_RBN1962_FE_OFN1591_n_13741), .o(n_16243) );
na02s02 TIMEBOOST_cell_39772 ( .a(g58095_sb), .b(FE_OFN245_n_9114), .o(TIMEBOOST_net_11498) );
in01m01 g64907_u0 ( .a(FE_OFN624_n_4409), .o(g64907_sb) );
in01s01 TIMEBOOST_cell_67729 ( .a(pci_target_unit_fifos_pcir_data_in_187), .o(TIMEBOOST_net_21156) );
na02m01 g64907_u2 ( .a(FE_OFN624_n_4409), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q), .o(g64907_db) );
in01m04 g64908_u0 ( .a(FE_OFN625_n_4409), .o(g64908_sb) );
na03m02 TIMEBOOST_cell_73197 ( .a(g65335_db), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q), .c(TIMEBOOST_net_12898), .o(TIMEBOOST_net_13238) );
in01m01 g64909_u0 ( .a(FE_OFN625_n_4409), .o(g64909_sb) );
na03f02 TIMEBOOST_cell_73467 ( .a(TIMEBOOST_net_17391), .b(FE_OFN1289_n_4098), .c(g62886_sb), .o(n_6105) );
na02m02 g64909_u2 ( .a(n_4403), .b(FE_OFN625_n_4409), .o(g64909_db) );
in01m06 g64910_u0 ( .a(FE_OFN625_n_4409), .o(g64910_sb) );
na02s01 TIMEBOOST_cell_25399 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_93), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6804) );
na03m02 TIMEBOOST_cell_72467 ( .a(TIMEBOOST_net_14078), .b(g65863_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_23230) );
in01m02 g64911_u0 ( .a(FE_OFN622_n_4409), .o(g64911_sb) );
na03m02 TIMEBOOST_cell_72481 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q), .b(FE_OFN1786_n_1699), .c(TIMEBOOST_net_21384), .o(n_1594) );
in01m02 g64912_u0 ( .a(FE_OFN623_n_4409), .o(g64912_sb) );
na02f02 TIMEBOOST_cell_45428 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13608), .o(TIMEBOOST_net_12039) );
na02f02 TIMEBOOST_cell_38781 ( .a(TIMEBOOST_net_11002), .b(g52625_sb), .o(n_14681) );
in01m01 g64913_u0 ( .a(FE_OFN625_n_4409), .o(g64913_sb) );
na03f02 TIMEBOOST_cell_68019 ( .a(TIMEBOOST_net_17421), .b(FE_OFN1260_n_4143), .c(g62377_sb), .o(n_6849) );
na02s01 TIMEBOOST_cell_38523 ( .a(TIMEBOOST_net_10873), .b(g58198_db), .o(n_9588) );
in01m01 g64914_u0 ( .a(FE_OFN622_n_4409), .o(g64914_sb) );
na03f02 TIMEBOOST_cell_66507 ( .a(TIMEBOOST_net_17105), .b(FE_OFN1322_n_6436), .c(g62351_sb), .o(n_6898) );
na03f02 TIMEBOOST_cell_35103 ( .a(TIMEBOOST_net_10024), .b(FE_OFN2155_n_16439), .c(g58827_sb), .o(n_8613) );
in01m02 g64915_u0 ( .a(FE_OFN624_n_4409), .o(g64915_sb) );
na04m06 TIMEBOOST_cell_72837 ( .a(n_3774), .b(g64774_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q), .d(g64774_db), .o(TIMEBOOST_net_17069) );
in01m08 g64916_u0 ( .a(FE_OFN622_n_4409), .o(g64916_sb) );
na02m01 TIMEBOOST_cell_53435 ( .a(TIMEBOOST_net_10731), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q), .o(TIMEBOOST_net_16935) );
na02f02 TIMEBOOST_cell_70251 ( .a(TIMEBOOST_net_22333), .b(g63039_sb), .o(n_7125) );
in01m02 g64917_u0 ( .a(FE_OFN1663_n_4490), .o(g64917_sb) );
na02f02 g59382_u2 ( .a(n_2987), .b(FE_OFN1699_n_5751), .o(g59382_db) );
in01m01 g64918_u0 ( .a(FE_OFN662_n_4392), .o(g64918_sb) );
na03f02 TIMEBOOST_cell_73666 ( .a(TIMEBOOST_net_17578), .b(FE_OFN1285_n_4097), .c(g62668_sb), .o(n_6201) );
in01m04 g64919_u0 ( .a(FE_OFN1810_n_4454), .o(g64919_sb) );
in01s01 TIMEBOOST_cell_73923 ( .a(TIMEBOOST_net_23487), .o(TIMEBOOST_net_23488) );
na03f02 TIMEBOOST_cell_66921 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_16498), .c(FE_OFN1513_n_14987), .o(n_12685) );
in01m01 g64920_u0 ( .a(FE_OFN618_n_4490), .o(g64920_sb) );
in01m01 g64921_u0 ( .a(FE_OFN660_n_4392), .o(g64921_sb) );
na02f08 TIMEBOOST_cell_69471 ( .a(TIMEBOOST_net_21943), .b(n_13341), .o(TIMEBOOST_net_20457) );
na02m02 TIMEBOOST_cell_68173 ( .a(TIMEBOOST_net_21294), .b(TIMEBOOST_net_12276), .o(TIMEBOOST_net_16810) );
in01m04 g64922_u0 ( .a(FE_OFN660_n_4392), .o(g64922_sb) );
na02s01 TIMEBOOST_cell_53876 ( .a(TIMEBOOST_net_17155), .b(TIMEBOOST_net_12978), .o(TIMEBOOST_net_9391) );
na03m06 TIMEBOOST_cell_65099 ( .a(n_3774), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q), .c(FE_OFN649_n_4497), .o(TIMEBOOST_net_12689) );
na02m01 TIMEBOOST_cell_47756 ( .a(TIMEBOOST_net_14095), .b(FE_OFN959_n_2299), .o(TIMEBOOST_net_10319) );
in01m01 g64923_u0 ( .a(FE_OFN661_n_4392), .o(g64923_sb) );
na03f02 TIMEBOOST_cell_73468 ( .a(TIMEBOOST_net_17464), .b(FE_OFN1288_n_4098), .c(g62482_sb), .o(n_6623) );
in01m02 g64924_u0 ( .a(FE_OFN660_n_4392), .o(g64924_sb) );
na02m02 TIMEBOOST_cell_72048 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q), .b(g65838_sb), .o(TIMEBOOST_net_23232) );
na04m01 TIMEBOOST_cell_67132 ( .a(TIMEBOOST_net_6769), .b(g54171_sb), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_386), .d(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q), .o(TIMEBOOST_net_16808) );
in01s01 TIMEBOOST_cell_73860 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_), .o(TIMEBOOST_net_23425) );
in01m01 g64925_u0 ( .a(FE_OFN619_n_4490), .o(g64925_sb) );
na03s01 TIMEBOOST_cell_64712 ( .a(pci_target_unit_del_sync_addr_in_229), .b(g66406_sb), .c(g66406_db), .o(n_2533) );
na03f02 TIMEBOOST_cell_34774 ( .a(TIMEBOOST_net_9327), .b(FE_OFN1377_n_8567), .c(g57166_sb), .o(n_10459) );
in01m04 g64926_u0 ( .a(FE_OFN662_n_4392), .o(g64926_sb) );
na03f02 TIMEBOOST_cell_66493 ( .a(TIMEBOOST_net_17138), .b(FE_OFN1316_n_6624), .c(g63159_sb), .o(n_5819) );
na02m08 g64926_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q), .b(FE_OFN662_n_4392), .o(g64926_db) );
in01s01 TIMEBOOST_cell_72356 ( .a(pci_target_unit_fifos_pcir_data_in_175), .o(TIMEBOOST_net_23389) );
in01m01 g64927_u0 ( .a(FE_OFN662_n_4392), .o(g64927_sb) );
na03m02 TIMEBOOST_cell_72796 ( .a(TIMEBOOST_net_23167), .b(g64857_sb), .c(TIMEBOOST_net_21833), .o(TIMEBOOST_net_16781) );
in01m01 g64928_u0 ( .a(FE_OFN661_n_4392), .o(g64928_sb) );
na03f02 TIMEBOOST_cell_66702 ( .a(TIMEBOOST_net_17493), .b(FE_OFN2063_n_6391), .c(g62457_sb), .o(n_6682) );
na03m02 TIMEBOOST_cell_70170 ( .a(FE_OFN1075_n_4740), .b(pci_target_unit_fifos_pciw_addr_data_in_128), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q), .o(TIMEBOOST_net_22293) );
in01m01 g64929_u0 ( .a(FE_OFN661_n_4392), .o(g64929_sb) );
na02m01 g64929_u2 ( .a(FE_OFN661_n_4392), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q), .o(g64929_db) );
na04f04 TIMEBOOST_cell_67929 ( .a(n_2198), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q), .c(FE_OFN720_n_8060), .d(g61699_sb), .o(n_8430) );
in01m02 g64930_u0 ( .a(FE_OFN660_n_4392), .o(g64930_sb) );
na03s01 TIMEBOOST_cell_32487 ( .a(g58015_sb), .b(FE_OFN217_n_9889), .c(g58015_db), .o(n_9777) );
na03m02 TIMEBOOST_cell_72483 ( .a(TIMEBOOST_net_14052), .b(g65958_db), .c(TIMEBOOST_net_22040), .o(TIMEBOOST_net_14768) );
in01m01 g64931_u0 ( .a(FE_OFN659_n_4392), .o(g64931_sb) );
na02m03 TIMEBOOST_cell_69280 ( .a(n_4498), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_21848) );
na02s02 TIMEBOOST_cell_43773 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_12781) );
in01m01 g64932_u0 ( .a(FE_OFN660_n_4392), .o(g64932_sb) );
na03m02 TIMEBOOST_cell_64673 ( .a(g64884_sb), .b(FE_OFN686_n_4417), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q), .o(TIMEBOOST_net_9700) );
na02m01 g64932_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q), .b(FE_OFN660_n_4392), .o(g64932_db) );
na02f01 TIMEBOOST_cell_51848 ( .a(TIMEBOOST_net_16141), .b(n_15755), .o(TIMEBOOST_net_169) );
in01m02 g64933_u0 ( .a(FE_OFN664_n_4495), .o(g64933_sb) );
na02m02 g64933_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q), .b(FE_OFN664_n_4495), .o(g64933_db) );
in01m01 g64934_u0 ( .a(FE_OFN660_n_4392), .o(g64934_sb) );
in01m01 g64935_u0 ( .a(FE_OFN661_n_4392), .o(g64935_sb) );
na02s01 TIMEBOOST_cell_68615 ( .a(TIMEBOOST_net_21515), .b(FE_OFN1016_n_2053), .o(TIMEBOOST_net_20373) );
na03f01 TIMEBOOST_cell_68118 ( .a(TIMEBOOST_net_14000), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q), .o(TIMEBOOST_net_21267) );
na02m01 TIMEBOOST_cell_69282 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q), .o(TIMEBOOST_net_21849) );
in01m06 g64936_u0 ( .a(FE_OFN661_n_4392), .o(g64936_sb) );
na03s02 TIMEBOOST_cell_32488 ( .a(g58213_sb), .b(FE_OFN227_n_9841), .c(g58213_db), .o(n_9572) );
na03f02 TIMEBOOST_cell_66399 ( .a(TIMEBOOST_net_17023), .b(FE_OFN1242_n_4092), .c(g62591_sb), .o(n_6371) );
na02m08 TIMEBOOST_cell_53025 ( .a(configuration_pci_err_addr_486), .b(wbm_adr_o_16_), .o(TIMEBOOST_net_16730) );
in01m06 g64937_u0 ( .a(FE_OFN659_n_4392), .o(g64937_sb) );
na02m02 TIMEBOOST_cell_69283 ( .a(TIMEBOOST_net_21849), .b(TIMEBOOST_net_9700), .o(TIMEBOOST_net_17104) );
na02m02 TIMEBOOST_cell_31377 ( .a(pci_target_unit_fifos_pciw_addr_data_in_138), .b(FE_OFN917_n_4725), .o(TIMEBOOST_net_9793) );
in01m04 g64938_u0 ( .a(FE_OFN659_n_4392), .o(g64938_sb) );
na03f02 TIMEBOOST_cell_73421 ( .a(TIMEBOOST_net_20533), .b(FE_OFN1250_n_4093), .c(g62683_sb), .o(n_6173) );
na02f01 TIMEBOOST_cell_70556 ( .a(TIMEBOOST_net_13051), .b(FE_OFN1112_g64577_p), .o(TIMEBOOST_net_22486) );
in01m01 g64939_u0 ( .a(FE_OFN659_n_4392), .o(g64939_sb) );
na04f04 TIMEBOOST_cell_72643 ( .a(TIMEBOOST_net_21408), .b(g59239_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q), .d(FE_OFN1083_n_13221), .o(TIMEBOOST_net_22869) );
na02f01 g64939_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q), .b(FE_OFN659_n_4392), .o(g64939_db) );
na02s03 TIMEBOOST_cell_54017 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q), .o(TIMEBOOST_net_17226) );
in01m04 g64940_u0 ( .a(FE_OFN659_n_4392), .o(g64940_sb) );
na03m06 TIMEBOOST_cell_72194 ( .a(FE_OFN1077_n_4740), .b(TIMEBOOST_net_16659), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q), .o(TIMEBOOST_net_23305) );
na03m04 TIMEBOOST_cell_72485 ( .a(n_3761), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q), .c(TIMEBOOST_net_12472), .o(TIMEBOOST_net_20580) );
na02m10 TIMEBOOST_cell_45611 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q), .o(TIMEBOOST_net_13700) );
in01m01 g64941_u0 ( .a(FE_OFN649_n_4497), .o(g64941_sb) );
na04f04 TIMEBOOST_cell_66925 ( .a(TIMEBOOST_net_503), .b(n_13711), .c(n_14384), .d(n_14087), .o(n_14532) );
in01m06 g64942_u0 ( .a(FE_OFN646_n_4497), .o(g64942_sb) );
in01s01 TIMEBOOST_cell_63542 ( .a(TIMEBOOST_net_20722), .o(wbs_adr_i_6_) );
na02m02 TIMEBOOST_cell_69090 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q), .b(FE_OFN1643_n_4671), .o(TIMEBOOST_net_21753) );
in01m01 g64943_u0 ( .a(FE_OFN648_n_4497), .o(g64943_sb) );
na03m01 TIMEBOOST_cell_68438 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q), .c(FE_OFN1003_n_2047), .o(TIMEBOOST_net_21427) );
na03f02 TIMEBOOST_cell_65619 ( .a(TIMEBOOST_net_20385), .b(g65681_sb), .c(g65681_db), .o(TIMEBOOST_net_13081) );
na03f02 TIMEBOOST_cell_46671 ( .a(TIMEBOOST_net_12868), .b(g64231_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q), .o(TIMEBOOST_net_13099) );
in01m01 g64944_u0 ( .a(FE_OFN649_n_4497), .o(g64944_sb) );
in01s01 TIMEBOOST_cell_73911 ( .a(TIMEBOOST_net_23475), .o(TIMEBOOST_net_23476) );
na02f02 TIMEBOOST_cell_70675 ( .a(TIMEBOOST_net_22545), .b(g63152_sb), .o(n_4959) );
in01m01 g64945_u0 ( .a(FE_OFN649_n_4497), .o(g64945_sb) );
na02f02 TIMEBOOST_cell_50952 ( .a(TIMEBOOST_net_15693), .b(g62596_sb), .o(n_6361) );
na02m01 g64945_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q), .b(FE_OFN649_n_4497), .o(g64945_db) );
na03f02 TIMEBOOST_cell_73344 ( .a(n_3238), .b(n_2768), .c(n_3237), .o(TIMEBOOST_net_22930) );
in01m08 g64946_u0 ( .a(FE_OFN649_n_4497), .o(g64946_sb) );
na02m10 TIMEBOOST_cell_45613 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q), .o(TIMEBOOST_net_13701) );
na04f04 TIMEBOOST_cell_73678 ( .a(n_3960), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q), .c(FE_OFN1137_g64577_p), .d(g62857_sb), .o(n_5253) );
in01m04 g64947_u0 ( .a(FE_OFN649_n_4497), .o(g64947_sb) );
na02m02 TIMEBOOST_cell_72076 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q), .b(g64252_sb), .o(TIMEBOOST_net_23246) );
na02m06 g64947_u2 ( .a(FE_OFN649_n_4497), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q), .o(g64947_db) );
in01m02 g64948_u0 ( .a(FE_OFN649_n_4497), .o(g64948_sb) );
na02s01 TIMEBOOST_cell_62526 ( .a(pci_target_unit_fifos_pcir_data_in_186), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q), .o(TIMEBOOST_net_20210) );
na02f02 TIMEBOOST_cell_71137 ( .a(TIMEBOOST_net_22776), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_14782) );
in01m01 g64949_u0 ( .a(FE_OFN647_n_4497), .o(g64949_sb) );
na03f04 TIMEBOOST_cell_72849 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q), .b(g65418_sb), .c(TIMEBOOST_net_22019), .o(TIMEBOOST_net_17016) );
na02m01 TIMEBOOST_cell_48662 ( .a(TIMEBOOST_net_14548), .b(TIMEBOOST_net_5420), .o(n_2652) );
in01m01 g64950_u0 ( .a(FE_OFN647_n_4497), .o(g64950_sb) );
na02m01 g52483_u1 ( .a(wbs_adr_i_7_), .b(g52470_sb), .o(g52483_da) );
na02m02 g64950_u2 ( .a(n_3665), .b(FE_OFN647_n_4497), .o(g64950_db) );
na02f01 TIMEBOOST_cell_47576 ( .a(TIMEBOOST_net_14005), .b(n_2237), .o(TIMEBOOST_net_124) );
in01m01 g64951_u0 ( .a(FE_OFN649_n_4497), .o(g64951_sb) );
na02s02 TIMEBOOST_cell_63219 ( .a(TIMEBOOST_net_20556), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_12807) );
na02m03 TIMEBOOST_cell_69613 ( .a(TIMEBOOST_net_22014), .b(FE_OFN1032_n_4732), .o(TIMEBOOST_net_20415) );
in01m01 g64952_u0 ( .a(FE_OFN646_n_4497), .o(g64952_sb) );
na02s02 TIMEBOOST_cell_38194 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(g65798_sb), .o(TIMEBOOST_net_10709) );
na02m01 g64952_u2 ( .a(n_74), .b(FE_OFN646_n_4497), .o(g64952_db) );
na03f02 TIMEBOOST_cell_47315 ( .a(FE_OFN1552_n_12104), .b(FE_OCP_RBN1978_n_10273), .c(TIMEBOOST_net_13599), .o(n_12637) );
in01m01 g64953_u0 ( .a(n_4460), .o(g64953_sb) );
na02s01 TIMEBOOST_cell_53633 ( .a(FE_OFN1666_n_9477), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q), .o(TIMEBOOST_net_17034) );
na03f02 TIMEBOOST_cell_66946 ( .a(FE_OFN1572_n_11027), .b(TIMEBOOST_net_13611), .c(FE_OFN1752_n_12086), .o(n_12697) );
in01m01 g64954_u0 ( .a(FE_OFN649_n_4497), .o(g64954_sb) );
na02s01 TIMEBOOST_cell_42810 ( .a(TIMEBOOST_net_12299), .b(FE_OFN937_n_2292), .o(TIMEBOOST_net_10238) );
in01s01 TIMEBOOST_cell_73935 ( .a(TIMEBOOST_net_23499), .o(TIMEBOOST_net_23500) );
na04f02 TIMEBOOST_cell_73422 ( .a(n_4357), .b(FE_OFN1223_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q), .d(g62507_sb), .o(n_6566) );
in01m01 g64955_u0 ( .a(FE_OFN648_n_4497), .o(g64955_sb) );
na02m10 TIMEBOOST_cell_71848 ( .a(TIMEBOOST_net_13891), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q), .o(TIMEBOOST_net_23132) );
in01m04 g64956_u0 ( .a(FE_OFN648_n_4497), .o(g64956_sb) );
na02m10 TIMEBOOST_cell_45615 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q), .o(TIMEBOOST_net_13702) );
na02m02 TIMEBOOST_cell_70111 ( .a(TIMEBOOST_net_22263), .b(TIMEBOOST_net_12746), .o(TIMEBOOST_net_17365) );
in01m01 g64957_u0 ( .a(FE_OFN646_n_4497), .o(g64957_sb) );
in01s01 TIMEBOOST_cell_73831 ( .a(TIMEBOOST_net_23395), .o(TIMEBOOST_net_23396) );
in01m01 g64958_u0 ( .a(FE_OFN646_n_4497), .o(g64958_sb) );
na03m02 TIMEBOOST_cell_73013 ( .a(TIMEBOOST_net_21625), .b(g64875_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q), .o(TIMEBOOST_net_13241) );
na03f08 TIMEBOOST_cell_35094 ( .a(g75181_db), .b(n_16271), .c(FE_OCP_RBN2233_n_16273), .o(n_16554) );
na03m02 TIMEBOOST_cell_65210 ( .a(TIMEBOOST_net_10684), .b(g64284_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q), .o(TIMEBOOST_net_20915) );
in01m01 g64959_u0 ( .a(FE_OFN612_n_4501), .o(g64959_sb) );
na03f02 TIMEBOOST_cell_66215 ( .a(TIMEBOOST_net_17446), .b(FE_OFN1243_n_4092), .c(g62548_sb), .o(n_6470) );
na03f02 TIMEBOOST_cell_34776 ( .a(TIMEBOOST_net_9365), .b(FE_OFN1399_n_8567), .c(g57237_sb), .o(n_11519) );
na02s01 TIMEBOOST_cell_68911 ( .a(TIMEBOOST_net_21663), .b(TIMEBOOST_net_12905), .o(TIMEBOOST_net_17035) );
in01m01 g64960_u0 ( .a(FE_OFN612_n_4501), .o(g64960_sb) );
na03f02 TIMEBOOST_cell_73797 ( .a(TIMEBOOST_net_13750), .b(FE_OFN1601_n_13995), .c(FE_OFN1605_n_13997), .o(n_14514) );
in01m01 g64961_u0 ( .a(FE_OFN614_n_4501), .o(g64961_sb) );
na02s02 TIMEBOOST_cell_44142 ( .a(TIMEBOOST_net_12965), .b(FE_OFN1801_n_9690), .o(TIMEBOOST_net_11174) );
in01s01 TIMEBOOST_cell_63604 ( .a(TIMEBOOST_net_20784), .o(TIMEBOOST_net_20731) );
na02m02 TIMEBOOST_cell_49697 ( .a(n_3510), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q), .o(TIMEBOOST_net_15066) );
in01m02 g64962_u0 ( .a(FE_OFN615_n_4501), .o(g64962_sb) );
na03m02 TIMEBOOST_cell_72813 ( .a(TIMEBOOST_net_21587), .b(g64924_sb), .c(TIMEBOOST_net_23240), .o(TIMEBOOST_net_9955) );
na02m02 g64962_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q), .b(FE_OFN615_n_4501), .o(g64962_db) );
in01s01 TIMEBOOST_cell_73899 ( .a(TIMEBOOST_net_23463), .o(TIMEBOOST_net_23464) );
in01m01 g64963_u0 ( .a(FE_OFN618_n_4490), .o(g64963_sb) );
na02s02 TIMEBOOST_cell_52367 ( .a(g58234_sb), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_16401) );
na02s01 TIMEBOOST_cell_70086 ( .a(n_8498), .b(n_1823), .o(TIMEBOOST_net_22251) );
na02s02 TIMEBOOST_cell_52368 ( .a(TIMEBOOST_net_16401), .b(g58249_db), .o(n_9544) );
na02f02 TIMEBOOST_cell_71058 ( .a(TIMEBOOST_net_17379), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_22737) );
na03f02 TIMEBOOST_cell_34778 ( .a(TIMEBOOST_net_9367), .b(FE_OFN1401_n_8567), .c(g57092_sb), .o(n_11650) );
in01m08 g64965_u0 ( .a(FE_OFN1807_n_4501), .o(g64965_sb) );
na03f02 TIMEBOOST_cell_34878 ( .a(TIMEBOOST_net_9324), .b(FE_OFN1377_n_8567), .c(g57557_sb), .o(n_10300) );
na03f02 TIMEBOOST_cell_34879 ( .a(TIMEBOOST_net_9431), .b(FE_OFN1420_n_8567), .c(g57244_sb), .o(n_11513) );
in01m01 g64966_u0 ( .a(FE_OFN665_n_4495), .o(g64966_sb) );
na02m01 g64966_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q), .b(FE_OFN665_n_4495), .o(g64966_db) );
in01m02 g64967_u0 ( .a(FE_OFN619_n_4490), .o(g64967_sb) );
na03f02 TIMEBOOST_cell_66542 ( .a(g53932_sb), .b(FE_OFN1326_n_13547), .c(TIMEBOOST_net_16806), .o(n_13513) );
na03f02 TIMEBOOST_cell_34780 ( .a(TIMEBOOST_net_9517), .b(FE_OFN1400_n_8567), .c(g57509_sb), .o(n_11230) );
na02f02 TIMEBOOST_cell_50720 ( .a(TIMEBOOST_net_15577), .b(n_13919), .o(n_14308) );
in01m01 g64968_u0 ( .a(FE_OFN618_n_4490), .o(g64968_sb) );
na04m04 TIMEBOOST_cell_67416 ( .a(TIMEBOOST_net_14511), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q), .c(g65395_sb), .d(FE_OFN1678_n_4655), .o(TIMEBOOST_net_17051) );
na02s01 TIMEBOOST_cell_48492 ( .a(TIMEBOOST_net_14463), .b(g58431_sb), .o(TIMEBOOST_net_12574) );
in01m04 g64969_u0 ( .a(FE_OFN615_n_4501), .o(g64969_sb) );
na03f02 TIMEBOOST_cell_34782 ( .a(TIMEBOOST_net_9379), .b(FE_OFN1377_n_8567), .c(g57433_sb), .o(n_10823) );
na02s02 TIMEBOOST_cell_69286 ( .a(TIMEBOOST_net_17227), .b(FE_OFN956_n_1699), .o(TIMEBOOST_net_21851) );
in01m02 g64970_u0 ( .a(FE_OFN667_n_4495), .o(g64970_sb) );
na03f02 TIMEBOOST_cell_73182 ( .a(TIMEBOOST_net_14591), .b(FE_OFN717_n_8176), .c(g61874_sb), .o(n_8084) );
na03f02 TIMEBOOST_cell_66604 ( .a(TIMEBOOST_net_17059), .b(n_6287), .c(g62969_sb), .o(n_5944) );
in01m01 g64971_u0 ( .a(FE_OFN615_n_4501), .o(g64971_sb) );
na03f02 TIMEBOOST_cell_34784 ( .a(TIMEBOOST_net_9529), .b(FE_OFN1390_n_8567), .c(g57301_sb), .o(n_11449) );
in01m02 g64972_u0 ( .a(FE_OFN1807_n_4501), .o(g64972_sb) );
na02s02 TIMEBOOST_cell_29141 ( .a(g58223_sb), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_8675) );
na02m01 TIMEBOOST_cell_68560 ( .a(n_50), .b(FE_OFN625_n_4409), .o(TIMEBOOST_net_21488) );
na02s01 TIMEBOOST_cell_29142 ( .a(TIMEBOOST_net_8675), .b(g58223_db), .o(n_9050) );
in01m01 g64973_u0 ( .a(FE_OFN1807_n_4501), .o(g64973_sb) );
na03f02 TIMEBOOST_cell_34910 ( .a(TIMEBOOST_net_9487), .b(FE_OFN1399_n_8567), .c(g57273_sb), .o(n_11482) );
na02m01 g64973_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q), .b(FE_OFN1807_n_4501), .o(g64973_db) );
na02s02 TIMEBOOST_cell_48214 ( .a(TIMEBOOST_net_14324), .b(g57896_sb), .o(TIMEBOOST_net_9465) );
in01m06 g64974_u0 ( .a(FE_OFN647_n_4497), .o(g64974_sb) );
na03f02 TIMEBOOST_cell_73738 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q), .b(FE_OFN1742_n_11019), .c(TIMEBOOST_net_16029), .o(n_12716) );
na02f01 TIMEBOOST_cell_52061 ( .a(TIMEBOOST_net_12410), .b(FE_OFN1013_n_4734), .o(TIMEBOOST_net_16248) );
na02m01 TIMEBOOST_cell_43628 ( .a(TIMEBOOST_net_12708), .b(FE_OFN1051_n_16657), .o(TIMEBOOST_net_10959) );
in01m01 g64975_u0 ( .a(FE_OFN622_n_4409), .o(g64975_sb) );
na02s01 TIMEBOOST_cell_31329 ( .a(g58243_sb), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_9769) );
na03f20 TIMEBOOST_cell_72391 ( .a(wishbone_slave_unit_pcim_if_wbw_cbe_in), .b(TIMEBOOST_net_12253), .c(n_294), .o(n_13548) );
na03f02 TIMEBOOST_cell_34779 ( .a(TIMEBOOST_net_9368), .b(FE_OFN1400_n_8567), .c(g57171_sb), .o(n_11585) );
in01m01 g64976_u0 ( .a(FE_OFN615_n_4501), .o(g64976_sb) );
na03f02 TIMEBOOST_cell_34786 ( .a(TIMEBOOST_net_9538), .b(FE_OFN1422_n_8567), .c(g57403_sb), .o(n_11338) );
na03f02 TIMEBOOST_cell_65918 ( .a(g62105_sb), .b(FE_OFN1174_n_5592), .c(TIMEBOOST_net_16406), .o(n_5595) );
in01f01 g64977_u0 ( .a(FE_OFN1623_n_4438), .o(g64977_sb) );
na02m04 TIMEBOOST_cell_69680 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q), .b(FE_OFN1676_n_4655), .o(TIMEBOOST_net_22048) );
na02m01 g64977_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q), .b(FE_OFN1623_n_4438), .o(g64977_db) );
na02m02 TIMEBOOST_cell_53989 ( .a(n_3764), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q), .o(TIMEBOOST_net_17212) );
in01m01 g64978_u0 ( .a(FE_OFN665_n_4495), .o(g64978_sb) );
na02s01 TIMEBOOST_cell_51866 ( .a(TIMEBOOST_net_16150), .b(FE_OFN595_n_9694), .o(TIMEBOOST_net_10348) );
na02s01 TIMEBOOST_cell_68318 ( .a(g64896_sb), .b(n_3780), .o(TIMEBOOST_net_21367) );
in01m02 g64979_u0 ( .a(FE_OFN619_n_4490), .o(g64979_sb) );
na03s02 TIMEBOOST_cell_46615 ( .a(TIMEBOOST_net_12837), .b(g63619_sb), .c(g63619_db), .o(n_7200) );
na03f02 TIMEBOOST_cell_34788 ( .a(TIMEBOOST_net_9540), .b(FE_OFN1411_n_8567), .c(g57318_sb), .o(n_11433) );
na03f02 TIMEBOOST_cell_73423 ( .a(TIMEBOOST_net_21022), .b(FE_OFN1268_n_4095), .c(g62410_sb), .o(n_6778) );
in01m01 g64980_u0 ( .a(FE_OFN685_n_4417), .o(g64980_sb) );
na02m02 TIMEBOOST_cell_68682 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q), .b(g64330_sb), .o(TIMEBOOST_net_21549) );
na02m01 TIMEBOOST_cell_69126 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q), .b(FE_OFN1644_n_4671), .o(TIMEBOOST_net_21771) );
na02s01 TIMEBOOST_cell_31330 ( .a(TIMEBOOST_net_9769), .b(g58243_db), .o(n_9045) );
na03s02 TIMEBOOST_cell_46510 ( .a(FE_OFN1657_n_9502), .b(n_8892), .c(g58333_da), .o(n_9484) );
in01m01 g64982_u0 ( .a(FE_OFN1624_n_4438), .o(g64982_sb) );
na02f01 TIMEBOOST_cell_70252 ( .a(TIMEBOOST_net_9946), .b(FE_OFN1100_g64577_p), .o(TIMEBOOST_net_22334) );
na03f02 TIMEBOOST_cell_34759 ( .a(TIMEBOOST_net_9480), .b(FE_OFN1400_n_8567), .c(g57100_sb), .o(n_11647) );
in01m01 g64983_u0 ( .a(FE_OFN647_n_4497), .o(g64983_sb) );
na02m01 g64983_u2 ( .a(FE_OFN647_n_4497), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q), .o(g64983_db) );
na02m04 TIMEBOOST_cell_69193 ( .a(TIMEBOOST_net_21804), .b(g64298_sb), .o(n_3876) );
in01m02 g64984_u0 ( .a(FE_OFN649_n_4497), .o(g64984_sb) );
in01m04 g64985_u0 ( .a(FE_OFN1628_n_4438), .o(g64985_sb) );
na02f02 TIMEBOOST_cell_70733 ( .a(TIMEBOOST_net_22574), .b(g54151_sb), .o(n_13659) );
na02m01 TIMEBOOST_cell_68174 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_413), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q), .o(TIMEBOOST_net_21295) );
na02s01 TIMEBOOST_cell_68140 ( .a(g61885_sb), .b(wbs_dat_i_20_), .o(TIMEBOOST_net_21278) );
in01m01 g64986_u0 ( .a(FE_OFN667_n_4495), .o(g64986_sb) );
na02m01 g64986_u2 ( .a(FE_OFN667_n_4495), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q), .o(g64986_db) );
in01m01 g64987_u0 ( .a(FE_OFN689_n_4438), .o(g64987_sb) );
na03f02 TIMEBOOST_cell_66770 ( .a(TIMEBOOST_net_13369), .b(n_6554), .c(g62493_sb), .o(n_6598) );
na03s02 TIMEBOOST_cell_69654 ( .a(TIMEBOOST_net_10327), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q), .c(TIMEBOOST_net_14277), .o(TIMEBOOST_net_22035) );
in01m01 g64988_u0 ( .a(FE_OFN646_n_4497), .o(g64988_sb) );
na03m02 TIMEBOOST_cell_69180 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_139), .c(FE_OFN930_n_4730), .o(TIMEBOOST_net_21798) );
na02m02 TIMEBOOST_cell_69676 ( .a(n_4493), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q), .o(TIMEBOOST_net_22046) );
na03f02 TIMEBOOST_cell_73758 ( .a(TIMEBOOST_net_16056), .b(FE_OFN1774_n_13800), .c(FE_OFN1771_n_14054), .o(g53314_p) );
in01m04 g64989_u0 ( .a(FE_OFN684_n_4417), .o(g64989_sb) );
na03f02 TIMEBOOST_cell_34761 ( .a(TIMEBOOST_net_9332), .b(FE_OFN1413_n_8567), .c(g57362_sb), .o(n_10385) );
in01m02 g64990_u0 ( .a(FE_OFN1625_n_4438), .o(g64990_sb) );
na02s01 TIMEBOOST_cell_48723 ( .a(FE_OFN560_n_9895), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q), .o(TIMEBOOST_net_14579) );
na03f02 TIMEBOOST_cell_73739 ( .a(TIMEBOOST_net_13573), .b(FE_OFN1739_n_11019), .c(FE_OFN1734_n_16317), .o(n_12501) );
in01m04 g64991_u0 ( .a(FE_OFN1628_n_4438), .o(g64991_sb) );
in01m02 g64992_u0 ( .a(FE_OFN659_n_4392), .o(g64992_sb) );
na03f02 TIMEBOOST_cell_62916 ( .a(g61921_sb), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q), .c(FE_OFN716_n_8176), .o(TIMEBOOST_net_20405) );
in01m06 g64993_u0 ( .a(FE_OFN1624_n_4438), .o(g64993_sb) );
no03f06 TIMEBOOST_cell_64398 ( .a(FE_RN_328_0), .b(FE_RN_332_0), .c(FE_RN_330_0), .o(FE_RN_333_0) );
na03m02 TIMEBOOST_cell_72487 ( .a(n_40), .b(n_3764), .c(FE_OFN646_n_4497), .o(TIMEBOOST_net_10728) );
in01m04 g64994_u0 ( .a(FE_OFN661_n_4392), .o(g64994_sb) );
in01s04 TIMEBOOST_cell_67096 ( .a(TIMEBOOST_net_21130), .o(FE_OFN528_n_9899) );
in01s01 TIMEBOOST_cell_73949 ( .a(TIMEBOOST_net_23513), .o(TIMEBOOST_net_23514) );
na03f02 TIMEBOOST_cell_66495 ( .a(TIMEBOOST_net_17021), .b(FE_OFN1224_n_6391), .c(g62551_sb), .o(n_6463) );
in01m01 g64995_u0 ( .a(FE_OFN664_n_4495), .o(g64995_sb) );
na02m04 TIMEBOOST_cell_72338 ( .a(TIMEBOOST_net_15865), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_), .o(TIMEBOOST_net_23377) );
na02f01 g64995_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q), .b(FE_OFN664_n_4495), .o(g64995_db) );
na02f02 TIMEBOOST_cell_71922 ( .a(TIMEBOOST_net_16885), .b(FE_OFN916_n_4725), .o(TIMEBOOST_net_23169) );
in01m02 g64996_u0 ( .a(FE_OFN1624_n_4438), .o(g64996_sb) );
na03f02 TIMEBOOST_cell_34775 ( .a(TIMEBOOST_net_9376), .b(FE_OFN1403_n_8567), .c(g57438_sb), .o(n_10355) );
in01s01 TIMEBOOST_cell_63603 ( .a(TIMEBOOST_net_20783), .o(TIMEBOOST_net_20782) );
na04m06 TIMEBOOST_cell_67314 ( .a(n_4465), .b(g65095_sb), .c(TIMEBOOST_net_20814), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q), .o(TIMEBOOST_net_20596) );
in01m08 g64997_u0 ( .a(FE_OFN689_n_4438), .o(g64997_sb) );
na04f04 TIMEBOOST_cell_73424 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q), .b(n_4908), .c(FE_OFN365_n_4093), .d(g62676_sb), .o(n_7368) );
na04s02 TIMEBOOST_cell_73641 ( .a(FE_OFN518_n_9697), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q), .c(g58150_sb), .d(FE_OFN221_n_9846), .o(n_9642) );
na04f06 TIMEBOOST_cell_73329 ( .a(n_4031), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q), .c(FE_OFN1136_g64577_p), .d(g62768_sb), .o(n_5458) );
in01m01 g64998_u0 ( .a(FE_OFN1624_n_4438), .o(g64998_sb) );
na03f02 TIMEBOOST_cell_66916 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_16491), .c(FE_OFN1513_n_14987), .o(n_12733) );
na02m01 g64998_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q), .b(FE_OFN1624_n_4438), .o(g64998_db) );
na03f02 TIMEBOOST_cell_73642 ( .a(TIMEBOOST_net_17499), .b(FE_OFN1230_n_6391), .c(g63177_sb), .o(n_5794) );
in01m04 g64999_u0 ( .a(FE_OFN667_n_4495), .o(g64999_sb) );
na02f02 TIMEBOOST_cell_70495 ( .a(TIMEBOOST_net_22455), .b(g63090_sb), .o(n_5074) );
na02s01 TIMEBOOST_cell_43187 ( .a(FE_OFN219_n_9853), .b(g58176_sb), .o(TIMEBOOST_net_12488) );
ao22f02 g64_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q), .b(FE_OFN1529_n_10853), .c(FE_OFN1453_n_10588), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q), .o(n_15528) );
in01m02 g65000_u0 ( .a(FE_OFN1628_n_4438), .o(g65000_sb) );
na02s02 TIMEBOOST_cell_37594 ( .a(g58076_sb), .b(FE_OFN217_n_9889), .o(TIMEBOOST_net_10409) );
na02f01 TIMEBOOST_cell_63051 ( .a(TIMEBOOST_net_20472), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_15131) );
na02s02 TIMEBOOST_cell_37595 ( .a(TIMEBOOST_net_10409), .b(g58076_db), .o(n_9718) );
in01m02 g65001_u0 ( .a(FE_OFN662_n_4392), .o(g65001_sb) );
na03m04 TIMEBOOST_cell_72364 ( .a(pci_target_unit_fifos_pciw_control_in_155), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q), .c(FE_OFN1059_n_4727), .o(TIMEBOOST_net_23245) );
in01m01 g65002_u0 ( .a(FE_OFN647_n_4497), .o(g65002_sb) );
na02m02 g65002_u2 ( .a(n_139), .b(FE_OFN647_n_4497), .o(g65002_db) );
na02m10 TIMEBOOST_cell_52989 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q), .b(wishbone_slave_unit_pcim_sm_data_in_640), .o(TIMEBOOST_net_16712) );
in01m02 g65003_u0 ( .a(FE_OFN685_n_4417), .o(g65003_sb) );
na02m04 g65003_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN685_n_4417), .o(g65003_db) );
in01m01 g65004_u0 ( .a(FE_OFN666_n_4495), .o(g65004_sb) );
na02s01 TIMEBOOST_cell_48031 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q), .o(TIMEBOOST_net_14233) );
na02m02 g65004_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q), .b(FE_OFN666_n_4495), .o(g65004_db) );
na02f01 TIMEBOOST_cell_30959 ( .a(n_3006), .b(wbu_addr_in_259), .o(TIMEBOOST_net_9584) );
in01m01 g65005_u0 ( .a(FE_OFN661_n_4392), .o(g65005_sb) );
na03f02 TIMEBOOST_cell_34795 ( .a(TIMEBOOST_net_9546), .b(FE_OFN1397_n_8567), .c(g57226_sb), .o(n_10434) );
na03f02 TIMEBOOST_cell_66401 ( .a(TIMEBOOST_net_21023), .b(n_8590), .c(g59122_sb), .o(n_8585) );
na03m06 TIMEBOOST_cell_72619 ( .a(FE_OFN1013_n_4734), .b(TIMEBOOST_net_20250), .c(g64175_sb), .o(n_3991) );
in01m01 g65006_u0 ( .a(FE_OFN661_n_4392), .o(g65006_sb) );
na02m02 TIMEBOOST_cell_53536 ( .a(TIMEBOOST_net_16985), .b(n_5546), .o(TIMEBOOST_net_15228) );
in01m01 g65007_u0 ( .a(FE_OFN1625_n_4438), .o(g65007_sb) );
na04m02 TIMEBOOST_cell_67343 ( .a(TIMEBOOST_net_20243), .b(FE_OFN651_n_4508), .c(g65427_sb), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q), .o(TIMEBOOST_net_17142) );
in01m02 g65008_u0 ( .a(FE_OFN1625_n_4438), .o(g65008_sb) );
na02f01 TIMEBOOST_cell_72256 ( .a(TIMEBOOST_net_16743), .b(FE_OFN1182_n_3476), .o(TIMEBOOST_net_23336) );
na03f02 TIMEBOOST_cell_73705 ( .a(TIMEBOOST_net_16481), .b(n_12313), .c(FE_OFN1566_n_12502), .o(n_12600) );
na02s01 g66399_u2 ( .a(parchk_pci_ad_reg_in_1231), .b(n_2520), .o(g66399_db) );
in01m01 g65009_u0 ( .a(FE_OFN648_n_4497), .o(g65009_sb) );
na04f06 TIMEBOOST_cell_64461 ( .a(n_1208), .b(n_1189), .c(n_1169), .d(n_1037), .o(n_2233) );
na03f01 TIMEBOOST_cell_65106 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q), .b(n_3785), .c(FE_OFN681_n_4460), .o(TIMEBOOST_net_10603) );
in01m02 g65010_u0 ( .a(FE_OFN622_n_4409), .o(g65010_sb) );
na02s01 TIMEBOOST_cell_47908 ( .a(TIMEBOOST_net_14171), .b(FE_OFN950_n_2055), .o(TIMEBOOST_net_12483) );
na03f02 TIMEBOOST_cell_73759 ( .a(FE_OFN1774_n_13800), .b(TIMEBOOST_net_13702), .c(FE_OFN1770_n_14054), .o(g53210_p) );
in01m01 g65011_u0 ( .a(FE_OFN1625_n_4438), .o(g65011_sb) );
in01s01 TIMEBOOST_cell_73912 ( .a(n_2524), .o(TIMEBOOST_net_23477) );
in01m01 g65012_u0 ( .a(FE_OFN661_n_4392), .o(g65012_sb) );
na02f01 TIMEBOOST_cell_68970 ( .a(TIMEBOOST_net_16898), .b(FE_OFN1010_n_4734), .o(TIMEBOOST_net_21693) );
na03f02 TIMEBOOST_cell_72930 ( .a(g65287_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q), .c(TIMEBOOST_net_14513), .o(TIMEBOOST_net_17135) );
in01m06 g65013_u0 ( .a(FE_OFN625_n_4409), .o(g65013_sb) );
na02m02 TIMEBOOST_cell_52785 ( .a(TIMEBOOST_net_12680), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q), .o(TIMEBOOST_net_16610) );
in01m01 g65014_u0 ( .a(FE_OFN647_n_4497), .o(g65014_sb) );
na02m06 TIMEBOOST_cell_62524 ( .a(TIMEBOOST_net_12377), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_20209) );
in01m02 g65015_u0 ( .a(FE_OFN1628_n_4438), .o(g65015_sb) );
na03f02 TIMEBOOST_cell_46674 ( .a(n_4527), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q), .c(g62749_sb), .o(TIMEBOOST_net_13155) );
na02s01 TIMEBOOST_cell_71303 ( .a(TIMEBOOST_net_22859), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_20604) );
in01s01 TIMEBOOST_cell_63597 ( .a(TIMEBOOST_net_20777), .o(TIMEBOOST_net_20776) );
in01m01 g65016_u0 ( .a(FE_OFN622_n_4409), .o(g65016_sb) );
na02f01 TIMEBOOST_cell_70930 ( .a(TIMEBOOST_net_20972), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_22673) );
na03f02 TIMEBOOST_cell_72992 ( .a(TIMEBOOST_net_21917), .b(g65043_sb), .c(TIMEBOOST_net_22108), .o(TIMEBOOST_net_17580) );
na02s02 TIMEBOOST_cell_39778 ( .a(g58003_sb), .b(FE_OFN245_n_9114), .o(TIMEBOOST_net_11501) );
in01m02 g65017_u0 ( .a(FE_OFN646_n_4497), .o(g65017_sb) );
in01s01 TIMEBOOST_cell_73900 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(TIMEBOOST_net_23465) );
in01m01 g65018_u0 ( .a(FE_OFN1625_n_4438), .o(g65018_sb) );
na02m02 TIMEBOOST_cell_69242 ( .a(n_4479), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q), .o(TIMEBOOST_net_21829) );
in01s01 TIMEBOOST_cell_72351 ( .a(TIMEBOOST_net_23383), .o(TIMEBOOST_net_23384) );
na02m01 TIMEBOOST_cell_69012 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q), .b(FE_OFN652_n_4508), .o(TIMEBOOST_net_21714) );
in01m01 g65019_u0 ( .a(FE_OFN687_n_4417), .o(g65019_sb) );
na02f01 g65019_u1 ( .a(n_4645), .b(g65019_sb), .o(g65019_da) );
na02m01 g65019_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q), .b(FE_OFN687_n_4417), .o(g65019_db) );
na02s01 TIMEBOOST_cell_38599 ( .a(TIMEBOOST_net_10911), .b(g58013_db), .o(n_9102) );
in01m01 g65020_u0 ( .a(FE_OFN670_n_4505), .o(g65020_sb) );
na02m01 TIMEBOOST_cell_71990 ( .a(n_3777), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q), .o(TIMEBOOST_net_23203) );
na03s02 TIMEBOOST_cell_73183 ( .a(TIMEBOOST_net_10062), .b(g62070_sb), .c(TIMEBOOST_net_5642), .o(n_7828) );
na02m01 TIMEBOOST_cell_69250 ( .a(n_3783), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q), .o(TIMEBOOST_net_21833) );
in01m01 g65021_u0 ( .a(FE_OFN630_n_4454), .o(g65021_sb) );
na03f02 TIMEBOOST_cell_34821 ( .a(TIMEBOOST_net_9382), .b(FE_OFN1409_n_8567), .c(g57545_sb), .o(n_11198) );
in01m02 g65022_u0 ( .a(FE_OFN687_n_4417), .o(g65022_sb) );
na02s02 TIMEBOOST_cell_48935 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q), .b(FE_OFN956_n_1699), .o(TIMEBOOST_net_14685) );
na02f02 TIMEBOOST_cell_70609 ( .a(TIMEBOOST_net_22512), .b(g63134_sb), .o(n_4982) );
na03f02 TIMEBOOST_cell_66159 ( .a(TIMEBOOST_net_16748), .b(FE_OFN1181_n_3476), .c(g60628_sb), .o(n_5709) );
in01m01 g65023_u0 ( .a(FE_OFN667_n_4495), .o(g65023_sb) );
na02m02 TIMEBOOST_cell_42989 ( .a(pci_target_unit_fifos_pciw_addr_data_in_140), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q), .o(TIMEBOOST_net_12389) );
na02m02 g52473_u1 ( .a(g52457_sb), .b(wbs_adr_i_27_), .o(g52473_da) );
in01m01 g65024_u0 ( .a(FE_OFN630_n_4454), .o(g65024_sb) );
na03m04 TIMEBOOST_cell_72971 ( .a(g64956_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q), .c(TIMEBOOST_net_10727), .o(TIMEBOOST_net_17501) );
na02m02 TIMEBOOST_cell_70115 ( .a(TIMEBOOST_net_22265), .b(TIMEBOOST_net_12820), .o(TIMEBOOST_net_17012) );
in01m01 g65025_u0 ( .a(FE_OFN624_n_4409), .o(g65025_sb) );
na04m02 TIMEBOOST_cell_67264 ( .a(n_3749), .b(g64794_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q), .d(FE_OFN665_n_4495), .o(n_3760) );
na03f02 TIMEBOOST_cell_66902 ( .a(FE_OFN1749_n_12004), .b(TIMEBOOST_net_13559), .c(n_12010), .o(n_12737) );
na03f02 TIMEBOOST_cell_67089 ( .a(FE_OFN1596_n_13741), .b(n_13903), .c(TIMEBOOST_net_13791), .o(n_14410) );
in01m02 g65026_u0 ( .a(FE_OFN634_n_4454), .o(g65026_sb) );
in01m01 g65027_u0 ( .a(FE_OFN630_n_4454), .o(g65027_sb) );
na04f04 TIMEBOOST_cell_24192 ( .a(n_9684), .b(g57248_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q), .d(FE_OFN1385_n_8567), .o(n_11509) );
in01m01 g65028_u0 ( .a(FE_OFN665_n_4495), .o(g65028_sb) );
na02f01 g65856_u2 ( .a(FE_OFN948_n_2248), .b(TIMEBOOST_net_20727), .o(g65856_db) );
in01m01 g65029_u0 ( .a(FE_OFN685_n_4417), .o(g65029_sb) );
na02m02 TIMEBOOST_cell_69498 ( .a(n_4645), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q), .o(TIMEBOOST_net_21957) );
na03m02 TIMEBOOST_cell_69082 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q), .b(FE_OFN1012_n_4734), .c(pci_target_unit_fifos_pciw_addr_data_in_126), .o(TIMEBOOST_net_21749) );
na04f04 TIMEBOOST_cell_47201 ( .a(FE_OFN2102_n_2834), .b(n_3505), .c(n_4826), .d(n_6978), .o(n_7338) );
in01m06 g65030_u0 ( .a(FE_OFN634_n_4454), .o(g65030_sb) );
na03f02 TIMEBOOST_cell_68021 ( .a(TIMEBOOST_net_17027), .b(FE_OFN1260_n_4143), .c(g62521_sb), .o(n_6534) );
na02f02 TIMEBOOST_cell_70809 ( .a(TIMEBOOST_net_22612), .b(g62047_sb), .o(n_7764) );
in01m01 g65031_u0 ( .a(FE_OFN685_n_4417), .o(g65031_sb) );
na02f02 TIMEBOOST_cell_63189 ( .a(TIMEBOOST_net_20541), .b(FE_OFN1275_n_4096), .o(TIMEBOOST_net_15352) );
na02m06 TIMEBOOST_cell_52753 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q), .o(TIMEBOOST_net_16594) );
in01m01 g65032_u0 ( .a(FE_OFN660_n_4392), .o(g65032_sb) );
na02m01 TIMEBOOST_cell_68617 ( .a(TIMEBOOST_net_21516), .b(FE_OFN927_n_4730), .o(TIMEBOOST_net_14667) );
na02f02 TIMEBOOST_cell_70611 ( .a(TIMEBOOST_net_22513), .b(g63032_sb), .o(n_5183) );
na02f02 TIMEBOOST_cell_69657 ( .a(TIMEBOOST_net_22036), .b(FE_OFN714_n_8140), .o(TIMEBOOST_net_14795) );
in01m01 g65033_u0 ( .a(FE_OFN629_n_4454), .o(g65033_sb) );
na02s04 TIMEBOOST_cell_62460 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q), .o(TIMEBOOST_net_20177) );
na02m01 g65033_u2 ( .a(FE_OFN629_n_4454), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q), .o(g65033_db) );
na03s01 TIMEBOOST_cell_72408 ( .a(pci_target_unit_fifos_pcir_data_in), .b(n_2299), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q), .o(TIMEBOOST_net_14055) );
in01m04 g65034_u0 ( .a(FE_OFN633_n_4454), .o(g65034_sb) );
na02s01 TIMEBOOST_cell_47624 ( .a(TIMEBOOST_net_14029), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_398), .o(n_13180) );
na03f02 TIMEBOOST_cell_66749 ( .a(TIMEBOOST_net_17136), .b(FE_OFN1313_n_6624), .c(g62956_sb), .o(n_5969) );
in01m01 g65035_u0 ( .a(FE_OFN1810_n_4454), .o(g65035_sb) );
na02s01 TIMEBOOST_cell_43016 ( .a(TIMEBOOST_net_12402), .b(FE_OFN229_n_9120), .o(TIMEBOOST_net_9371) );
na03f02 TIMEBOOST_cell_73706 ( .a(TIMEBOOST_net_13526), .b(n_12313), .c(FE_OFN1562_n_12502), .o(n_12655) );
na03f02 TIMEBOOST_cell_73469 ( .a(TIMEBOOST_net_17523), .b(FE_OFN1253_n_4143), .c(g62631_sb), .o(n_6292) );
in01m01 g65036_u0 ( .a(FE_OFN618_n_4490), .o(g65036_sb) );
na03s02 TIMEBOOST_cell_72464 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q), .b(g65853_sb), .c(g65853_db), .o(n_1583) );
na02s01 TIMEBOOST_cell_45249 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q), .o(TIMEBOOST_net_13519) );
na02m02 TIMEBOOST_cell_43508 ( .a(TIMEBOOST_net_12648), .b(g65724_db), .o(n_1610) );
in01m02 g65037_u0 ( .a(FE_OFN684_n_4417), .o(g65037_sb) );
na02f02 TIMEBOOST_cell_49900 ( .a(TIMEBOOST_net_15167), .b(g63049_sb), .o(n_5153) );
na04f04 TIMEBOOST_cell_73643 ( .a(TIMEBOOST_net_22889), .b(TIMEBOOST_net_675), .c(n_3131), .d(g62031_sb), .o(n_13509) );
in01m01 g65038_u0 ( .a(FE_OFN633_n_4454), .o(g65038_sb) );
na04f04 TIMEBOOST_cell_47205 ( .a(TIMEBOOST_net_13490), .b(FE_OFN2198_n_10256), .c(g52616_sb), .d(TIMEBOOST_net_695), .o(n_11854) );
na02s02 TIMEBOOST_cell_62646 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q), .b(FE_OFN227_n_9841), .o(TIMEBOOST_net_20270) );
na03f02 TIMEBOOST_cell_73264 ( .a(TIMEBOOST_net_17296), .b(FE_OFN2212_n_8407), .c(g61825_sb), .o(n_8137) );
in01m01 g65039_u0 ( .a(FE_OFN623_n_4409), .o(g65039_sb) );
in01s01 TIMEBOOST_cell_73950 ( .a(wbm_dat_i_25_), .o(TIMEBOOST_net_23515) );
in01m02 g65040_u0 ( .a(FE_OFN1809_n_4454), .o(g65040_sb) );
na02m10 TIMEBOOST_cell_38112 ( .a(g64273_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q), .o(TIMEBOOST_net_10668) );
na02s01 TIMEBOOST_cell_70435 ( .a(TIMEBOOST_net_22425), .b(FE_OFN577_n_9902), .o(TIMEBOOST_net_14935) );
na02f04 TIMEBOOST_cell_70204 ( .a(TIMEBOOST_net_14864), .b(FE_OFN1148_n_13249), .o(TIMEBOOST_net_22310) );
in01m01 g65041_u0 ( .a(FE_OFN625_n_4409), .o(g65041_sb) );
na04f02 TIMEBOOST_cell_73198 ( .a(TIMEBOOST_net_14946), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q), .c(FE_OFN1095_g64577_p), .d(g61957_sb), .o(n_6958) );
na02m06 TIMEBOOST_cell_52754 ( .a(TIMEBOOST_net_16594), .b(g65921_sb), .o(TIMEBOOST_net_14325) );
na03m04 TIMEBOOST_cell_72489 ( .a(n_3783), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q), .c(TIMEBOOST_net_16156), .o(TIMEBOOST_net_17047) );
in01m01 g65042_u0 ( .a(FE_OFN649_n_4497), .o(g65042_sb) );
na02s02 TIMEBOOST_cell_62915 ( .a(TIMEBOOST_net_20404), .b(g58073_sb), .o(TIMEBOOST_net_9523) );
in01m01 g65043_u0 ( .a(FE_OFN647_n_4497), .o(g65043_sb) );
na02s02 TIMEBOOST_cell_68619 ( .a(TIMEBOOST_net_21517), .b(FE_OFN1017_n_2053), .o(TIMEBOOST_net_16291) );
na02s02 TIMEBOOST_cell_48827 ( .a(g58035_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q), .o(TIMEBOOST_net_14631) );
na02m01 TIMEBOOST_cell_62952 ( .a(g57923_sb), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_20423) );
in01m01 g65044_u0 ( .a(FE_OFN625_n_4409), .o(g65044_sb) );
na02m02 TIMEBOOST_cell_49170 ( .a(TIMEBOOST_net_14802), .b(g61791_sb), .o(n_8218) );
na02s02 TIMEBOOST_cell_71365 ( .a(TIMEBOOST_net_22890), .b(g57904_sb), .o(TIMEBOOST_net_15212) );
na02m02 TIMEBOOST_cell_68300 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q), .b(n_4669), .o(TIMEBOOST_net_21358) );
in01m02 g65045_u0 ( .a(FE_OFN1810_n_4454), .o(g65045_sb) );
na04f04 TIMEBOOST_cell_67931 ( .a(n_2293), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q), .c(FE_OFN720_n_8060), .d(g61701_sb), .o(n_8426) );
na03f01 TIMEBOOST_cell_72463 ( .a(n_8884), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q), .c(wbu_addr_in_252), .o(TIMEBOOST_net_12386) );
in01m01 g65046_u0 ( .a(FE_OFN624_n_4409), .o(g65046_sb) );
na02f02 TIMEBOOST_cell_52460 ( .a(TIMEBOOST_net_16447), .b(g60626_sb), .o(n_5712) );
na03f02 TIMEBOOST_cell_34790 ( .a(TIMEBOOST_net_9543), .b(FE_OFN1420_n_8567), .c(g57274_sb), .o(n_11480) );
in01m01 g65047_u0 ( .a(FE_OFN631_n_4454), .o(g65047_sb) );
na03f02 TIMEBOOST_cell_34853 ( .a(TIMEBOOST_net_9509), .b(FE_OFN1380_n_8567), .c(g57293_sb), .o(n_10410) );
na02s01 TIMEBOOST_cell_39786 ( .a(g58063_sb), .b(FE_OFN245_n_9114), .o(TIMEBOOST_net_11505) );
in01m01 g65048_u0 ( .a(FE_OFN646_n_4497), .o(g65048_sb) );
na02m10 TIMEBOOST_cell_68094 ( .a(n_2078), .b(n_16690), .o(TIMEBOOST_net_21255) );
in01m01 g65049_u0 ( .a(FE_OFN687_n_4417), .o(g65049_sb) );
na02m04 TIMEBOOST_cell_31353 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(g65786_sb), .o(TIMEBOOST_net_9781) );
na02s01 TIMEBOOST_cell_52756 ( .a(TIMEBOOST_net_16595), .b(g57968_db), .o(TIMEBOOST_net_9501) );
na03f02 TIMEBOOST_cell_72851 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q), .b(g64971_sb), .c(TIMEBOOST_net_14421), .o(TIMEBOOST_net_17118) );
in01m01 g65050_u0 ( .a(FE_OFN687_n_4417), .o(g65050_sb) );
na02f02 TIMEBOOST_cell_52852 ( .a(TIMEBOOST_net_16643), .b(g61913_sb), .o(n_7995) );
na02m02 TIMEBOOST_cell_50022 ( .a(TIMEBOOST_net_15228), .b(g63194_sb), .o(n_4798) );
na03m02 TIMEBOOST_cell_70880 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q), .b(FE_OFN561_n_9895), .c(FE_OFN231_n_9839), .o(TIMEBOOST_net_22648) );
in01m01 g65051_u0 ( .a(FE_OFN648_n_4497), .o(g65051_sb) );
na02m08 TIMEBOOST_cell_69700 ( .a(FE_OFN1680_n_4655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q), .o(TIMEBOOST_net_22058) );
na03f02 TIMEBOOST_cell_47415 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q), .b(n_12066), .c(n_11831), .o(n_12486) );
in01m01 g65052_u0 ( .a(FE_OFN666_n_4495), .o(g65052_sb) );
na02s02 TIMEBOOST_cell_70723 ( .a(TIMEBOOST_net_22569), .b(FE_OFN1671_n_9477), .o(TIMEBOOST_net_20945) );
in01s01 TIMEBOOST_cell_73951 ( .a(TIMEBOOST_net_23515), .o(TIMEBOOST_net_23516) );
in01m08 g65053_u0 ( .a(FE_OFN620_n_4490), .o(g65053_sb) );
na03f04 TIMEBOOST_cell_73579 ( .a(TIMEBOOST_net_17522), .b(FE_OFN1085_n_13221), .c(g54197_sb), .o(n_13421) );
na03s01 TIMEBOOST_cell_64738 ( .a(pci_target_unit_del_sync_addr_in_232), .b(g66415_sb), .c(g66422_db), .o(n_2505) );
in01m01 g65054_u0 ( .a(FE_OFN618_n_4490), .o(g65054_sb) );
na02m01 TIMEBOOST_cell_69284 ( .a(n_4465), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q), .o(TIMEBOOST_net_21850) );
na03f02 TIMEBOOST_cell_65917 ( .a(TIMEBOOST_net_20433), .b(FE_OFN1166_n_5615), .c(g62129_sb), .o(n_5567) );
in01s04 TIMEBOOST_cell_67098 ( .a(TIMEBOOST_net_21132), .o(FE_OFN533_n_9823) );
in01m01 g65055_u0 ( .a(FE_OFN620_n_4490), .o(g65055_sb) );
na02f02 TIMEBOOST_cell_53651 ( .a(TIMEBOOST_net_13240), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_17043) );
na02m02 TIMEBOOST_cell_70409 ( .a(TIMEBOOST_net_22412), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_15133) );
in01m01 g65056_u0 ( .a(FE_OFN624_n_4409), .o(g65056_sb) );
na02f02 TIMEBOOST_cell_52290 ( .a(TIMEBOOST_net_16362), .b(g52627_sb), .o(TIMEBOOST_net_14894) );
na02s02 TIMEBOOST_cell_49292 ( .a(TIMEBOOST_net_14863), .b(TIMEBOOST_net_10853), .o(TIMEBOOST_net_9541) );
in01m01 g65057_u0 ( .a(n_4460), .o(g65057_sb) );
na02m04 g52469_u1 ( .a(wbs_adr_i_23_), .b(g52458_sb), .o(g52469_da) );
na02m01 g65057_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q), .b(n_4460), .o(g65057_db) );
in01m01 g65058_u0 ( .a(FE_OFN619_n_4490), .o(g65058_sb) );
na02s02 TIMEBOOST_cell_69287 ( .a(TIMEBOOST_net_21851), .b(g65771_sb), .o(n_1602) );
na02m01 g65058_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q), .b(FE_OFN619_n_4490), .o(g65058_db) );
na04m10 TIMEBOOST_cell_67419 ( .a(g58161_sb), .b(FE_OFN239_n_9832), .c(FE_OFN515_n_9697), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q), .o(n_9627) );
in01m04 g65059_u0 ( .a(FE_OFN1663_n_4490), .o(g65059_sb) );
na02s02 TIMEBOOST_cell_53272 ( .a(TIMEBOOST_net_16853), .b(TIMEBOOST_net_12872), .o(TIMEBOOST_net_9564) );
na02m02 TIMEBOOST_cell_69970 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q), .b(g64314_sb), .o(TIMEBOOST_net_22193) );
na02f01 TIMEBOOST_cell_70411 ( .a(TIMEBOOST_net_22413), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_15122) );
in01m04 g65060_u0 ( .a(FE_OFN667_n_4495), .o(g65060_sb) );
na02f01 TIMEBOOST_cell_30961 ( .a(n_2488), .b(wbu_addr_in_255), .o(TIMEBOOST_net_9585) );
in01m04 g65061_u0 ( .a(FE_OFN1663_n_4490), .o(g65061_sb) );
na02m02 TIMEBOOST_cell_49689 ( .a(n_3506), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q), .o(TIMEBOOST_net_15062) );
na02m02 TIMEBOOST_cell_68328 ( .a(n_14), .b(n_4669), .o(TIMEBOOST_net_21372) );
na02m02 TIMEBOOST_cell_69296 ( .a(n_4476), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q), .o(TIMEBOOST_net_21856) );
in01m04 g65062_u0 ( .a(FE_OFN1663_n_4490), .o(g65062_sb) );
na02f01 TIMEBOOST_cell_68306 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q), .b(n_4460), .o(TIMEBOOST_net_21361) );
in01m02 g65063_u0 ( .a(FE_OFN681_n_4460), .o(g65063_sb) );
na02s02 TIMEBOOST_cell_43797 ( .a(FE_OFN233_n_9876), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q), .o(TIMEBOOST_net_12793) );
na02m04 g65063_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q), .b(FE_OFN681_n_4460), .o(g65063_db) );
na03f02 TIMEBOOST_cell_65919 ( .a(TIMEBOOST_net_20436), .b(FE_OFN1170_n_5592), .c(g62126_sb), .o(n_5570) );
in01m02 g65064_u0 ( .a(FE_OFN1810_n_4454), .o(g65064_sb) );
na02s02 TIMEBOOST_cell_54618 ( .a(TIMEBOOST_net_17526), .b(g58178_sb), .o(TIMEBOOST_net_9436) );
in01m01 g65065_u0 ( .a(FE_OFN662_n_4392), .o(g65065_sb) );
na02m01 g65065_u2 ( .a(FE_OFN662_n_4392), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q), .o(g65065_db) );
na02m01 TIMEBOOST_cell_53881 ( .a(pci_target_unit_pcit_if_strd_addr_in_716), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80), .o(TIMEBOOST_net_17158) );
in01m01 g65066_u0 ( .a(FE_OFN620_n_4490), .o(g65066_sb) );
na04m04 TIMEBOOST_cell_67933 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q), .b(FE_OFN1812_n_7845), .c(n_2152), .d(g62020_sb), .o(n_7855) );
in01m01 g65067_u0 ( .a(FE_OFN1663_n_4490), .o(g65067_sb) );
na02m01 TIMEBOOST_cell_50033 ( .a(configuration_pci_err_addr_484), .b(wbm_adr_o_14_), .o(TIMEBOOST_net_15234) );
na02m06 TIMEBOOST_cell_45251 ( .a(n_263), .b(n_323), .o(TIMEBOOST_net_13520) );
in01m01 g65068_u0 ( .a(FE_OFN618_n_4490), .o(g65068_sb) );
na04f02 TIMEBOOST_cell_67948 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q), .b(FE_OFN1115_g64577_p), .c(n_3843), .d(g63131_sb), .o(n_4988) );
na03f02 TIMEBOOST_cell_73525 ( .a(TIMEBOOST_net_17485), .b(n_6554), .c(g62382_sb), .o(n_6837) );
in01m01 g65069_u0 ( .a(n_4460), .o(g65069_sb) );
na02s01 TIMEBOOST_cell_49469 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_14952) );
na02m01 g65069_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q), .b(n_4460), .o(g65069_db) );
na02m10 TIMEBOOST_cell_49017 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_121), .o(TIMEBOOST_net_14726) );
in01m04 g65070_u0 ( .a(FE_OFN665_n_4495), .o(g65070_sb) );
na02m01 TIMEBOOST_cell_68305 ( .a(TIMEBOOST_net_21360), .b(g60689_sb), .o(n_3204) );
na02s01 TIMEBOOST_cell_30963 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_15__Q), .b(n_9856), .o(TIMEBOOST_net_9586) );
in01m02 g65071_u0 ( .a(FE_OFN631_n_4454), .o(g65071_sb) );
na02m10 TIMEBOOST_cell_52661 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q), .o(TIMEBOOST_net_16548) );
na02m04 TIMEBOOST_cell_44057 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_141), .o(TIMEBOOST_net_12923) );
in01m01 g65072_u0 ( .a(FE_OFN681_n_4460), .o(g65072_sb) );
na02m02 g65072_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q), .b(FE_OFN681_n_4460), .o(g65072_db) );
na03m02 TIMEBOOST_cell_73014 ( .a(TIMEBOOST_net_23180), .b(g65031_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q), .o(TIMEBOOST_net_16771) );
in01m01 g65073_u0 ( .a(FE_OFN660_n_4392), .o(g65073_sb) );
na03m04 TIMEBOOST_cell_72931 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q), .b(g65284_sb), .c(TIMEBOOST_net_23256), .o(TIMEBOOST_net_17426) );
na03f20 TIMEBOOST_cell_34640 ( .a(n_8747), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q), .c(n_8657), .o(n_15515) );
na02m02 TIMEBOOST_cell_50146 ( .a(TIMEBOOST_net_15290), .b(g60667_sb), .o(n_5651) );
in01m01 g65074_u0 ( .a(FE_OFN681_n_4460), .o(g65074_sb) );
in01m08 g65075_u0 ( .a(FE_OFN666_n_4495), .o(g65075_sb) );
na02m02 TIMEBOOST_cell_62520 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q), .o(TIMEBOOST_net_20207) );
na02m01 TIMEBOOST_cell_68178 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_407), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q), .o(TIMEBOOST_net_21297) );
in01m01 g65076_u0 ( .a(FE_OFN662_n_4392), .o(g65076_sb) );
na03m08 TIMEBOOST_cell_65112 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q), .c(FE_OFN618_n_4490), .o(TIMEBOOST_net_10615) );
na03f02 TIMEBOOST_cell_68024 ( .a(TIMEBOOST_net_17033), .b(FE_OFN1207_n_6356), .c(g63011_sb), .o(n_5862) );
in01m01 g65077_u0 ( .a(n_4460), .o(g65077_sb) );
na02m01 TIMEBOOST_cell_68526 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q), .b(n_3761), .o(TIMEBOOST_net_21471) );
na02m01 g65077_u2 ( .a(n_4460), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q), .o(g65077_db) );
na02s01 TIMEBOOST_cell_42839 ( .a(wbu_addr_in_263), .b(g58772_sb), .o(TIMEBOOST_net_12314) );
in01m01 g65078_u0 ( .a(FE_OFN681_n_4460), .o(g65078_sb) );
na02f04 TIMEBOOST_cell_44992 ( .a(TIMEBOOST_net_13390), .b(g54185_db), .o(g53939_db) );
na03m02 TIMEBOOST_cell_72750 ( .a(n_4465), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q), .c(TIMEBOOST_net_12543), .o(TIMEBOOST_net_21038) );
in01m01 g65079_u0 ( .a(FE_OFN631_n_4454), .o(g65079_sb) );
na02m02 g65079_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q), .b(FE_OFN631_n_4454), .o(g65079_db) );
in01m04 g65080_u0 ( .a(FE_OFN682_n_4460), .o(g65080_sb) );
na03f02 TIMEBOOST_cell_68023 ( .a(TIMEBOOST_net_17026), .b(FE_OFN1260_n_4143), .c(g62522_sb), .o(n_6532) );
na02m02 TIMEBOOST_cell_52908 ( .a(TIMEBOOST_net_16671), .b(g58097_db), .o(TIMEBOOST_net_9348) );
in01m01 g65081_u0 ( .a(FE_OFN624_n_4409), .o(g65081_sb) );
na02s02 TIMEBOOST_cell_30863 ( .a(n_9680), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q), .o(TIMEBOOST_net_9536) );
in01m02 g65082_u0 ( .a(FE_OFN678_n_4460), .o(g65082_sb) );
na02f02 TIMEBOOST_cell_70581 ( .a(TIMEBOOST_net_22498), .b(g63116_sb), .o(n_5023) );
in01s01 TIMEBOOST_cell_63602 ( .a(TIMEBOOST_net_20782), .o(TIMEBOOST_net_20723) );
in01m01 g65083_u0 ( .a(FE_OFN624_n_4409), .o(g65083_sb) );
na03s01 TIMEBOOST_cell_64739 ( .a(pci_target_unit_del_sync_addr_in_227), .b(g66415_sb), .c(g66424_db), .o(n_2502) );
na02m04 TIMEBOOST_cell_68962 ( .a(g65313_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q), .o(TIMEBOOST_net_21689) );
in01m04 g65084_u0 ( .a(FE_OFN682_n_4460), .o(g65084_sb) );
na02m01 TIMEBOOST_cell_38221 ( .a(TIMEBOOST_net_10722), .b(TIMEBOOST_net_5435), .o(n_2643) );
in01m01 g65085_u0 ( .a(FE_OFN662_n_4392), .o(g65085_sb) );
na03m02 TIMEBOOST_cell_73425 ( .a(TIMEBOOST_net_17147), .b(FE_OFN1219_n_6886), .c(g62347_sb), .o(n_6905) );
in01s01 TIMEBOOST_cell_73952 ( .a(wbm_dat_i_26_), .o(TIMEBOOST_net_23517) );
in01m01 g65086_u0 ( .a(FE_OFN682_n_4460), .o(g65086_sb) );
na02f02 TIMEBOOST_cell_39575 ( .a(TIMEBOOST_net_11399), .b(g62796_sb), .o(n_5393) );
na02s01 TIMEBOOST_cell_48397 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q), .b(FE_OFN225_n_9122), .o(TIMEBOOST_net_14416) );
na02f02 TIMEBOOST_cell_69989 ( .a(TIMEBOOST_net_22202), .b(g61792_sb), .o(n_8215) );
in01m01 g65087_u0 ( .a(FE_OFN662_n_4392), .o(g65087_sb) );
in01m01 g65088_u0 ( .a(FE_OFN659_n_4392), .o(g65088_sb) );
na02s02 TIMEBOOST_cell_54543 ( .a(g58216_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q), .o(TIMEBOOST_net_17489) );
na02m02 TIMEBOOST_cell_69615 ( .a(TIMEBOOST_net_22015), .b(FE_OFN1032_n_4732), .o(TIMEBOOST_net_20417) );
in01m01 g65089_u0 ( .a(FE_OFN669_n_4505), .o(g65089_sb) );
na03m02 TIMEBOOST_cell_72863 ( .a(TIMEBOOST_net_21719), .b(g64751_sb), .c(TIMEBOOST_net_21952), .o(TIMEBOOST_net_17560) );
na02m04 TIMEBOOST_cell_48216 ( .a(TIMEBOOST_net_14325), .b(g65921_db), .o(TIMEBOOST_net_13394) );
na02f01 TIMEBOOST_cell_48218 ( .a(TIMEBOOST_net_14326), .b(g64977_db), .o(n_3650) );
in01m01 g65090_u0 ( .a(FE_OFN666_n_4495), .o(g65090_sb) );
na02m02 TIMEBOOST_cell_69008 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q), .b(FE_OFN651_n_4508), .o(TIMEBOOST_net_21712) );
na04f04 TIMEBOOST_cell_72641 ( .a(TIMEBOOST_net_21482), .b(g53939_sb), .c(wishbone_slave_unit_pcim_if_wbw_cbe_in_417), .d(FE_OFN1083_n_13221), .o(TIMEBOOST_net_23365) );
na02m01 TIMEBOOST_cell_48681 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q), .o(TIMEBOOST_net_14558) );
in01m01 g65091_u0 ( .a(FE_OFN667_n_4495), .o(g65091_sb) );
na02s01 TIMEBOOST_cell_53634 ( .a(TIMEBOOST_net_17034), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_11116) );
na02s01 TIMEBOOST_cell_42805 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q), .o(TIMEBOOST_net_12297) );
in01m01 g65092_u0 ( .a(FE_OFN618_n_4490), .o(g65092_sb) );
na04f04 TIMEBOOST_cell_24195 ( .a(n_9793), .b(g57128_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q), .d(FE_OFN1417_n_8567), .o(n_11617) );
na03f02 TIMEBOOST_cell_73265 ( .a(TIMEBOOST_net_12968), .b(g61958_sb), .c(g61958_db), .o(n_6956) );
in01m04 g65093_u0 ( .a(FE_OFN686_n_4417), .o(g65093_sb) );
in01s01 TIMEBOOST_cell_73832 ( .a(pci_rst_oe_o), .o(TIMEBOOST_net_23397) );
na02m06 g65093_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q), .b(FE_OFN686_n_4417), .o(g65093_db) );
na03f02 TIMEBOOST_cell_65673 ( .a(TIMEBOOST_net_20387), .b(FE_OFN2128_n_16497), .c(g54306_sb), .o(n_13026) );
in01m01 g65094_u0 ( .a(FE_OFN625_n_4409), .o(g65094_sb) );
na03f02 TIMEBOOST_cell_73825 ( .a(n_13891), .b(TIMEBOOST_net_16557), .c(FE_OFN1593_n_13741), .o(g53234_p) );
na03s01 TIMEBOOST_cell_70412 ( .a(FE_OFN223_n_9844), .b(FE_OFN1649_n_9428), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q), .o(TIMEBOOST_net_22414) );
na02f01 TIMEBOOST_cell_44354 ( .a(TIMEBOOST_net_13071), .b(FE_OFN1121_g64577_p), .o(TIMEBOOST_net_11389) );
in01m04 g65095_u0 ( .a(FE_OFN679_n_4460), .o(g65095_sb) );
na03f02 TIMEBOOST_cell_23121 ( .a(TIMEBOOST_net_343), .b(n_5743), .c(TIMEBOOST_net_5720), .o(n_7722) );
na02m01 TIMEBOOST_cell_53027 ( .a(configuration_pci_err_addr_495), .b(wbm_adr_o_25_), .o(TIMEBOOST_net_16731) );
na03f02 TIMEBOOST_cell_73470 ( .a(TIMEBOOST_net_17492), .b(FE_OFN1250_n_4093), .c(g62393_sb), .o(n_6812) );
in01m01 g65096_u0 ( .a(n_4417), .o(g65096_sb) );
na03m02 TIMEBOOST_cell_72865 ( .a(TIMEBOOST_net_21756), .b(g64861_sb), .c(TIMEBOOST_net_21971), .o(TIMEBOOST_net_17074) );
na02m01 g65096_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q), .b(n_4417), .o(g65096_db) );
in01m01 g65097_u0 ( .a(FE_OFN679_n_4460), .o(g65097_sb) );
na02s01 TIMEBOOST_cell_63258 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q), .b(FE_OFN516_n_9697), .o(TIMEBOOST_net_20576) );
in01m04 g65098_u0 ( .a(FE_OFN1660_n_4490), .o(g65098_sb) );
na02m02 TIMEBOOST_cell_68307 ( .a(TIMEBOOST_net_21361), .b(g64821_sb), .o(TIMEBOOST_net_12590) );
na02f01 TIMEBOOST_cell_44330 ( .a(TIMEBOOST_net_13059), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_11345) );
in01m01 g65099_u0 ( .a(FE_OFN669_n_4505), .o(g65099_sb) );
na02f02 TIMEBOOST_cell_70616 ( .a(TIMEBOOST_net_8324), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_22516) );
na02m02 g65099_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q), .b(FE_OFN669_n_4505), .o(g65099_db) );
na02f01 TIMEBOOST_cell_49698 ( .a(TIMEBOOST_net_15066), .b(FE_OFN1128_g64577_p), .o(TIMEBOOST_net_13174) );
ao22f02 g65101_u0 ( .a(configuration_wb_err_addr_547), .b(n_15444), .c(n_16000), .d(n_2831), .o(n_3072) );
in01f02 g65102_u0 ( .a(n_2871), .o(n_3071) );
ao22f06 g65103_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_517), .c(configuration_wb_err_data_586), .d(FE_OFN1069_n_15729), .o(n_2871) );
ao22f02 g65104_u0 ( .a(n_14919), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_525), .o(n_3070) );
ao22f02 g65105_u0 ( .a(configuration_wb_err_data_587), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2869), .o(n_2870) );
ao22f04 g65106_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_365), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_526), .o(n_3068) );
ao22f02 g65107_u0 ( .a(configuration_wb_err_addr_549), .b(n_15444), .c(n_16000), .d(n_2869), .o(n_3066) );
ao22f02 g65109_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_519), .c(n_14921), .d(n_16810), .o(n_2868) );
ao22f02 g65110_u0 ( .a(configuration_wb_err_data_588), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2866), .o(n_2867) );
ao22f02 g65111_u0 ( .a(configuration_wb_err_addr_550), .b(n_15444), .c(n_16000), .d(n_2866), .o(n_3064) );
ao22f02 g65112_u0 ( .a(configuration_wb_err_data_592), .b(FE_OFN1068_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2864), .o(n_2865) );
ao22f02 g65115_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_502), .c(n_3371), .d(wbu_pref_en_in_136), .o(n_3374) );
ao22f01 g65116_u0 ( .a(configuration_isr_bit_2975), .b(n_3246), .c(n_3248), .d(configuration_sync_command_bit1), .o(n_3245) );
ao22f04 g65117_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_521), .c(n_14923), .d(n_16810), .o(n_2775) );
ao22f04 g65118_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_368), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_529), .o(n_3062) );
ao22f02 g65119_u0 ( .a(configuration_wb_err_addr_552), .b(n_15444), .c(n_16000), .d(n_2835), .o(n_3061) );
ao22f02 g65120_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_522), .c(n_14924), .d(n_16810), .o(n_2860) );
ao22f02 g65121_u0 ( .a(n_3231), .b(pciu_bar0_in_370), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_531), .o(n_3060) );
ao22f01 g65122_u0 ( .a(configuration_wb_err_addr_554), .b(n_15444), .c(n_16000), .d(n_2864), .o(n_3059) );
ao22f04 g65125_u0 ( .a(FE_OFN1065_n_15808), .b(configuration_pci_err_data_523), .c(n_14925), .d(n_16810), .o(n_2859) );
ao22f02 g65126_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_518), .c(n_14920), .d(n_16810), .o(n_2858) );
ao22f02 g65127_u0 ( .a(configuration_wb_err_data_596), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2856), .o(n_2857) );
ao22f02 g65128_u0 ( .a(configuration_status_bit_435), .b(n_3248), .c(n_16000), .d(n_2841), .o(n_17048) );
ao22f02 g65129_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_529), .c(configuration_wb_err_cs_bit_567), .d(n_16543), .o(n_3241) );
ao22f02 g65130_u0 ( .a(configuration_status_bit_379), .b(n_3248), .c(n_16000), .d(n_2854), .o(n_17039) );
ao22f02 g65131_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_530), .c(configuration_wb_err_cs_bit_568), .d(n_16543), .o(n_17027) );
ao22f02 g65132_u0 ( .a(n_14932), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_538), .o(n_3058) );
ao22f02 g65133_u0 ( .a(configuration_wb_err_data_599), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2854), .o(n_2855) );
ao22f01 g65134_u0 ( .a(configuration_wb_err_data_573), .b(FE_OFN1071_n_15729), .c(configuration_wb_err_addr_535), .d(n_15445), .o(n_2853) );
ao22f02 g65135_u0 ( .a(n_3372), .b(n_14906), .c(n_3371), .d(n_14907), .o(n_3373) );
ao22f02 g65136_u0 ( .a(configuration_status_bit_351), .b(n_3248), .c(n_16000), .d(n_2851), .o(n_3238) );
ao22f02 g65137_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_531), .c(configuration_wb_err_cs_bit_569), .d(n_16543), .o(n_3237) );
ao22f02 g65138_u0 ( .a(n_14933), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_539), .o(n_3057) );
ao22f02 g65139_u0 ( .a(configuration_wb_err_data_600), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2851), .o(n_2852) );
ao22f02 g65141_u0 ( .a(configuration_wb_err_data_574), .b(FE_OFN1071_n_15729), .c(configuration_wb_err_addr_536), .d(n_15445), .o(n_2849) );
ao22f02 g65142_u0 ( .a(configuration_interrupt_line_40), .b(n_3295), .c(FE_OFN1695_n_3368), .d(wbu_cache_line_size_in_208), .o(n_3370) );
ao22f01 g65143_u0 ( .a(configuration_wb_err_data_575), .b(FE_OFN1071_n_15729), .c(configuration_wb_err_addr_537), .d(n_15445), .o(n_2848) );
ao22f02 g65144_u0 ( .a(configuration_wb_err_cs_bit_564), .b(n_16543), .c(n_3231), .d(pciu_bar0_in_373), .o(n_3236) );
ao22f04 g65145_u0 ( .a(configuration_wb_err_data_576), .b(FE_OFN1071_n_15729), .c(n_3248), .d(configuration_sync_command_bit6), .o(n_3235) );
ao22f08 g65146_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_507), .c(configuration_wb_err_addr_538), .d(n_15445), .o(n_2847) );
ao22f01 g65147_u0 ( .a(configuration_wb_err_data_577), .b(FE_OFN1071_n_15729), .c(configuration_wb_err_addr_539), .d(n_15445), .o(n_2846) );
ao22f02 g65148_u0 ( .a(configuration_interrupt_line_43), .b(n_3295), .c(FE_OFN1695_n_3368), .d(wbu_cache_line_size_in_211), .o(n_3367) );
ao22f01 g65151_u0 ( .a(configuration_wb_err_addr_546), .b(n_15444), .c(n_16000), .d(n_2809), .o(n_3055) );
ao22f04 g65152_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_366), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_527), .o(n_3054) );
ao22f02 g65153_u0 ( .a(configuration_status_bit_407), .b(n_3248), .c(n_16000), .d(n_2825), .o(n_3233) );
ao22f02 g65155_u0 ( .a(FE_OFN1065_n_15808), .b(configuration_pci_err_data_526), .c(n_16791), .d(pciu_bar0_in_373), .o(n_2843) );
ao22f02 g65156_u0 ( .a(configuration_wb_err_data_597), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2841), .o(n_2842) );
ao22f02 g65157_u0 ( .a(configuration_wb_err_cs_bit_565), .b(n_16543), .c(n_3231), .d(pciu_bar0_in_374), .o(n_3232) );
ao22f02 g65158_u0 ( .a(configuration_status_bit_322), .b(n_3504), .c(n_16000), .d(n_3592), .o(n_3593) );
ao22f02 g65159_u0 ( .a(FE_OFN1066_n_15808), .b(configuration_pci_err_data_528), .c(configuration_wb_err_cs_bit_566), .d(n_16543), .o(n_17034) );
ao22f02 g65160_u0 ( .a(FE_OFN1065_n_15808), .b(configuration_pci_err_data_527), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_535), .o(n_3053) );
ao22f06 g65161_u0 ( .a(configuration_wb_err_data_601), .b(FE_OFN1070_n_15729), .c(n_16810), .d(n_14934), .o(n_2840) );
ao22f01 g65162_u0 ( .a(n_3231), .b(pciu_bar0_in_379), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_540), .o(n_3052) );
ao22f01 g65163_u0 ( .a(n_16000), .b(n_2838), .c(n_15444), .d(configuration_wb_err_addr_541), .o(n_3051) );
ao22f02 g65164_u0 ( .a(n_14930), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_536), .o(n_3050) );
ao22f02 g65165_u0 ( .a(n_15808), .b(configuration_pci_err_data_532), .c(configuration_wb_err_cs_bit_570), .d(n_16543), .o(n_3229) );
ao22f02 g65166_u0 ( .a(FE_OCPN1845_n_16427), .b(n_2838), .c(FE_OFN1068_n_15729), .d(configuration_wb_err_data_579), .o(n_2839) );
ao22f01 g65168_u0 ( .a(n_3252), .b(configuration_pci_err_cs_bit9), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_243), .o(n_2969) );
ao22f02 g65169_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_363), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_524), .o(n_3049) );
ao22f04 g65170_u0 ( .a(configuration_wb_err_data_590), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2835), .o(n_2836) );
ao22f02 g65171_u0 ( .a(configuration_wb_err_data_595), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2833), .o(n_2834) );
ao22f04 g65173_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_369), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_530), .o(n_3048) );
ao22f02 g65174_u0 ( .a(n_14929), .b(n_16810), .c(n_16791), .d(pciu_bar0_in_374), .o(n_2830) );
ao22f02 g65175_u0 ( .a(configuration_wb_err_data_591), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2828), .o(n_2829) );
ao22f10 g65177_u0 ( .a(n_1724), .b(parchk_pci_trdy_en_in), .c(n_2804), .d(conf_wb_err_bc_in), .o(n_3047) );
ao22f02 g65178_u0 ( .a(configuration_wb_err_data_598), .b(FE_OFN1070_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2825), .o(n_2826) );
ao22f02 g65179_u0 ( .a(n_3371), .b(wbu_mrl_en_in_141), .c(FE_OCPN1845_n_16427), .d(pciu_am1_in_540), .o(n_3366) );
ao22f02 g65180_u0 ( .a(configuration_wb_err_cs_bit0), .b(n_16543), .c(n_3372), .d(wbu_mrl_en_in_142), .o(n_3228) );
ao22f01 g65181_u0 ( .a(configuration_cache_line_size_reg), .b(FE_OFN1695_n_3368), .c(n_16000), .d(pciu_am1_in_540), .o(n_3046) );
ao22f01 g65182_u0 ( .a(n_3252), .b(configuration_pci_err_cs_bit0), .c(configuration_interrupt_line), .d(n_3295), .o(n_3365) );
ao22f02 g65183_u0 ( .a(configuration_wb_err_addr_553), .b(n_15445), .c(n_16000), .d(n_2828), .o(n_3045) );
ao22f04 g65184_u0 ( .a(n_3252), .b(configuration_pci_err_cs_bit10), .c(FE_OFN1694_n_3368), .d(wbu_latency_tim_val_in_244), .o(n_2824) );
ao22f02 g65185_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_511), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_519), .o(n_3044) );
ao22f02 g65186_u0 ( .a(configuration_wb_err_data_580), .b(FE_OFN1068_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2822), .o(n_2823) );
ao22f01 g65187_u0 ( .a(configuration_wb_err_addr_542), .b(n_15445), .c(n_16000), .d(n_2822), .o(n_3043) );
na03f06 TIMEBOOST_cell_18549 ( .a(n_4674), .b(n_4675), .c(n_4874), .o(TIMEBOOST_net_5638) );
in01f02 g65189_u0 ( .a(n_2821), .o(n_3042) );
ao22f04 g65190_u0 ( .a(FE_OFN1065_n_15808), .b(configuration_pci_err_data_524), .c(configuration_wb_err_data_593), .d(FE_OFN1068_n_15729), .o(n_2821) );
ao22f02 g65191_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_512), .c(n_14914), .d(n_16810), .o(n_2820) );
ao22f02 g65192_u0 ( .a(configuration_wb_err_data_581), .b(FE_OFN1068_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2818), .o(n_2819) );
in01f02 g65193_u0 ( .a(n_3041), .o(n_3227) );
ao22f01 g65194_u0 ( .a(configuration_wb_err_addr_543), .b(n_15445), .c(n_16000), .d(n_2818), .o(n_3041) );
ao22f02 g65195_u0 ( .a(n_14931), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_537), .o(n_3040) );
ao22f02 g65196_u0 ( .a(n_14926), .b(n_16810), .c(FE_OFN2129_n_16720), .d(pciu_am1_in_532), .o(n_3039) );
ao22f02 g65201_u0 ( .a(n_14915), .b(n_16810), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_521), .o(n_3037) );
ao22f01 g65202_u0 ( .a(configuration_wb_err_addr_544), .b(n_15445), .c(n_16000), .d(n_16428), .o(n_3036) );
ao22f02 g65203_u0 ( .a(FE_OFN1063_n_15808), .b(configuration_pci_err_data_514), .c(n_14916), .d(n_16810), .o(n_2814) );
ao22f04 g65204_u0 ( .a(configuration_wb_err_data_583), .b(FE_OFN1069_n_15729), .c(FE_OCPN1845_n_16427), .d(n_2812), .o(n_2813) );
ao22f02 g65205_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_361), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_522), .o(n_3034) );
ao22f01 g65206_u0 ( .a(configuration_wb_err_addr_545), .b(n_15445), .c(n_16000), .d(n_2812), .o(n_3033) );
ao22f02 g65209_u0 ( .a(FE_OCPN1898_n_3231), .b(pciu_bar0_in_362), .c(FE_OFN1061_n_16720), .d(pciu_am1_in_523), .o(n_3032) );
in01f01 g65210_u0 ( .a(FE_OFN785_n_2678), .o(g65210_sb) );
na03f02 TIMEBOOST_cell_34877 ( .a(TIMEBOOST_net_9334), .b(FE_OFN1386_n_8567), .c(g57262_sb), .o(n_11492) );
na02s01 TIMEBOOST_cell_38593 ( .a(TIMEBOOST_net_10908), .b(g58066_db), .o(n_9726) );
in01f02 g65211_u0 ( .a(FE_OFN786_n_2678), .o(g65211_sb) );
na02f02 TIMEBOOST_cell_72153 ( .a(TIMEBOOST_net_23284), .b(g64366_sb), .o(TIMEBOOST_net_9986) );
na03f02 TIMEBOOST_cell_34911 ( .a(TIMEBOOST_net_9488), .b(FE_OFN1377_n_8567), .c(g57435_sb), .o(n_10357) );
na02s02 TIMEBOOST_cell_29146 ( .a(TIMEBOOST_net_8677), .b(g58002_sb), .o(n_9106) );
no02f04 TIMEBOOST_cell_51525 ( .a(FE_RN_734_0), .b(n_13725), .o(TIMEBOOST_net_15980) );
na02f01 g65212_u2 ( .a(pci_target_unit_wbm_sm_pci_tar_burst_ok), .b(n_2678), .o(g65212_db) );
in01s08 TIMEBOOST_cell_47505 ( .a(TIMEBOOST_net_13968), .o(FE_OFN597_n_9694) );
in01m01 g65213_u0 ( .a(FE_OFN789_n_2678), .o(g65213_sb) );
na03m08 TIMEBOOST_cell_65125 ( .a(n_3777), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q), .c(FE_OFN639_n_4669), .o(TIMEBOOST_net_14436) );
na02f02 TIMEBOOST_cell_63311 ( .a(TIMEBOOST_net_20602), .b(TIMEBOOST_net_13115), .o(TIMEBOOST_net_9415) );
in01f01 g65214_u0 ( .a(FE_OFN785_n_2678), .o(g65214_sb) );
na02f01 TIMEBOOST_cell_70333 ( .a(TIMEBOOST_net_22374), .b(g62111_db), .o(n_5587) );
na02m02 TIMEBOOST_cell_53882 ( .a(TIMEBOOST_net_17158), .b(n_16748), .o(TIMEBOOST_net_15944) );
na02m10 TIMEBOOST_cell_45617 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q), .o(TIMEBOOST_net_13703) );
in01f04 g65215_u0 ( .a(FE_OFN787_n_2678), .o(g65215_sb) );
na02m02 g64241_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_141), .b(FE_OFN917_n_4725), .o(g64241_db) );
na02s01 TIMEBOOST_cell_38587 ( .a(TIMEBOOST_net_10905), .b(g58089_db), .o(n_9707) );
in01s01 g65216_u0 ( .a(FE_OFN786_n_2678), .o(g65216_sb) );
na02f04 g54239_u2 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q), .b(FE_OFN1150_n_13249), .o(g54239_db) );
na03f02 TIMEBOOST_cell_35045 ( .a(TIMEBOOST_net_9589), .b(FE_OFN1439_n_9372), .c(g58464_sb), .o(n_9387) );
na03f20 TIMEBOOST_cell_41281 ( .a(n_1014), .b(n_709), .c(n_7705), .o(n_8569) );
in01f01 g65217_u0 ( .a(FE_OFN785_n_2678), .o(g65217_sb) );
na02s02 TIMEBOOST_cell_52451 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q), .b(g58295_sb), .o(TIMEBOOST_net_16443) );
na04f04 TIMEBOOST_cell_67633 ( .a(TIMEBOOST_net_20549), .b(g52443_sb), .c(n_3134), .d(FE_OFN1700_n_5751), .o(g52443_da) );
na03f02 TIMEBOOST_cell_35047 ( .a(TIMEBOOST_net_9597), .b(FE_OFN1441_n_9372), .c(g58457_sb), .o(n_9398) );
in01f01 g65218_u0 ( .a(FE_OFN785_n_2678), .o(g65218_sb) );
na02m01 g52467_u1 ( .a(wbs_adr_i_21_), .b(g52457_sb), .o(g52467_da) );
na02f02 TIMEBOOST_cell_68723 ( .a(TIMEBOOST_net_21569), .b(g65669_sb), .o(n_2029) );
in01f01 g65219_u0 ( .a(FE_OFN785_n_2678), .o(g65219_sb) );
na02m01 TIMEBOOST_cell_69026 ( .a(n_3774), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q), .o(TIMEBOOST_net_21721) );
na04f04 TIMEBOOST_cell_67470 ( .a(n_4265), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q), .c(FE_OFN1311_n_6624), .d(g63008_sb), .o(n_5866) );
na02s02 TIMEBOOST_cell_48789 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q), .b(g58344_sb), .o(TIMEBOOST_net_14612) );
in01f02 g65220_u0 ( .a(FE_OFN784_n_2678), .o(g65220_sb) );
na03f02 TIMEBOOST_cell_72518 ( .a(TIMEBOOST_net_14147), .b(g64135_sb), .c(g64135_db), .o(TIMEBOOST_net_9946) );
na03f02 TIMEBOOST_cell_66793 ( .a(TIMEBOOST_net_17164), .b(FE_OFN1230_n_6391), .c(g62985_sb), .o(n_5912) );
in01f01 g65221_u0 ( .a(FE_OFN789_n_2678), .o(g65221_sb) );
na03f06 TIMEBOOST_cell_66018 ( .a(TIMEBOOST_net_20926), .b(FE_OFN882_g64577_p), .c(g63051_sb), .o(n_5149) );
na03f02 TIMEBOOST_cell_34927 ( .a(TIMEBOOST_net_9496), .b(FE_OFN1399_n_8567), .c(g57202_sb), .o(n_11553) );
na03s02 TIMEBOOST_cell_48847 ( .a(g58256_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q), .c(TIMEBOOST_net_12904), .o(TIMEBOOST_net_14641) );
in01m01 g65222_u0 ( .a(FE_OFN784_n_2678), .o(g65222_sb) );
na02s01 TIMEBOOST_cell_47791 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q), .b(FE_OFN205_n_9140), .o(TIMEBOOST_net_14113) );
na02s01 TIMEBOOST_cell_38589 ( .a(TIMEBOOST_net_10906), .b(g58138_db), .o(n_9658) );
na02s02 TIMEBOOST_cell_38567 ( .a(TIMEBOOST_net_10895), .b(g57912_db), .o(n_9898) );
in01f01 g65223_u0 ( .a(FE_OFN785_n_2678), .o(g65223_sb) );
na02f02 TIMEBOOST_cell_49442 ( .a(TIMEBOOST_net_14938), .b(FE_OFN272_n_9828), .o(TIMEBOOST_net_9365) );
na02s01 TIMEBOOST_cell_38569 ( .a(TIMEBOOST_net_10896), .b(g58112_db), .o(n_9683) );
na02s01 TIMEBOOST_cell_38571 ( .a(TIMEBOOST_net_10897), .b(g58044_db), .o(n_9094) );
in01f02 g65224_u0 ( .a(FE_OFN784_n_2678), .o(g65224_sb) );
na02s01 TIMEBOOST_cell_38573 ( .a(TIMEBOOST_net_10898), .b(g58038_db), .o(n_9751) );
na02s01 TIMEBOOST_cell_38575 ( .a(TIMEBOOST_net_10899), .b(g58142_db), .o(n_9653) );
in01f02 g65225_u0 ( .a(FE_OFN786_n_2678), .o(g65225_sb) );
na02m02 TIMEBOOST_cell_68998 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q), .b(g65380_sb), .o(TIMEBOOST_net_21707) );
na02s01 TIMEBOOST_cell_48881 ( .a(FE_OFN601_n_9687), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q), .o(TIMEBOOST_net_14658) );
na03f02 TIMEBOOST_cell_73826 ( .a(TIMEBOOST_net_13806), .b(n_13903), .c(FE_OFN1596_n_13741), .o(n_14434) );
in01f01 g65226_u0 ( .a(FE_OFN785_n_2678), .o(g65226_sb) );
na02f02 g65905_u2 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(FE_OFN1059_n_4727), .o(g65905_db) );
na02m02 TIMEBOOST_cell_30551 ( .a(n_9006), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q), .o(TIMEBOOST_net_9380) );
na04m02 TIMEBOOST_cell_64989 ( .a(n_4470), .b(g65065_sb), .c(g65065_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q), .o(TIMEBOOST_net_17057) );
in01f02 g65227_u0 ( .a(FE_OFN785_n_2678), .o(g65227_sb) );
na02m02 TIMEBOOST_cell_68175 ( .a(TIMEBOOST_net_21295), .b(TIMEBOOST_net_14036), .o(TIMEBOOST_net_16795) );
na03s02 TIMEBOOST_cell_72532 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .b(n_8503), .c(FE_OFN2079_n_8069), .o(n_8504) );
in01f01 g65228_u0 ( .a(FE_OFN785_n_2678), .o(g65228_sb) );
na02f02 TIMEBOOST_cell_54604 ( .a(TIMEBOOST_net_17519), .b(FE_OFN1272_n_4096), .o(TIMEBOOST_net_15527) );
na02s01 TIMEBOOST_cell_70119 ( .a(TIMEBOOST_net_22267), .b(FE_OFN1795_n_9904), .o(TIMEBOOST_net_16380) );
in01m01 g65229_u0 ( .a(FE_OFN785_n_2678), .o(g65229_sb) );
na02s01 TIMEBOOST_cell_38807 ( .a(TIMEBOOST_net_11015), .b(g65858_sb), .o(n_2593) );
na02f02 TIMEBOOST_cell_70563 ( .a(TIMEBOOST_net_22489), .b(g62727_sb), .o(n_5526) );
in01f02 g65230_u0 ( .a(FE_OFN786_n_2678), .o(g65230_sb) );
na03f02 TIMEBOOST_cell_617 ( .a(n_4024), .b(g62777_sb), .c(g62777_db), .o(n_5438) );
na02f02 TIMEBOOST_cell_70627 ( .a(TIMEBOOST_net_22521), .b(g63100_sb), .o(n_5054) );
in01m01 g65231_u0 ( .a(FE_OFN784_n_2678), .o(g65231_sb) );
na02m02 TIMEBOOST_cell_68040 ( .a(pci_target_unit_del_sync_comp_cycle_count_2_), .b(pci_target_unit_del_sync_comp_cycle_count_1_), .o(TIMEBOOST_net_21228) );
na04f04 TIMEBOOST_cell_67093 ( .a(n_14055), .b(n_14226), .c(n_13982), .d(TIMEBOOST_net_16135), .o(n_16220) );
na03f02 TIMEBOOST_cell_34929 ( .a(TIMEBOOST_net_9519), .b(FE_OFN1404_n_8567), .c(g57422_sb), .o(n_10362) );
in01m01 g65232_u0 ( .a(FE_OFN789_n_2678), .o(g65232_sb) );
na02s03 TIMEBOOST_cell_47971 ( .a(pci_target_unit_fifos_pcir_data_in_188), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q), .o(TIMEBOOST_net_14203) );
na02s01 TIMEBOOST_cell_39192 ( .a(g57961_sb), .b(FE_OFN268_n_9880), .o(TIMEBOOST_net_11208) );
na02s02 TIMEBOOST_cell_39194 ( .a(g57948_sb), .b(FE_OFN260_n_9860), .o(TIMEBOOST_net_11209) );
in01f02 g65233_u0 ( .a(FE_OFN784_n_2678), .o(g65233_sb) );
na03f40 TIMEBOOST_cell_41569 ( .a(TIMEBOOST_net_10377), .b(n_2447), .c(n_4743), .o(g74576_p) );
na02s02 TIMEBOOST_cell_39196 ( .a(g57956_sb), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_11210) );
na03f02 TIMEBOOST_cell_68025 ( .a(TIMEBOOST_net_17025), .b(FE_OFN1253_n_4143), .c(g62895_sb), .o(n_6087) );
in01s01 TIMEBOOST_cell_73989 ( .a(TIMEBOOST_net_23553), .o(TIMEBOOST_net_23554) );
na02m02 TIMEBOOST_cell_68119 ( .a(TIMEBOOST_net_21267), .b(g61880_sb), .o(TIMEBOOST_net_17288) );
in01s01 g65235_u0 ( .a(FE_OFN786_n_2678), .o(g65235_sb) );
na04f02 TIMEBOOST_cell_25262 ( .a(n_14566), .b(n_14475), .c(n_14957), .d(n_14956), .o(n_14611) );
na02m10 TIMEBOOST_cell_45465 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q), .o(TIMEBOOST_net_13627) );
in01s01 g65236_u0 ( .a(FE_OFN786_n_2678), .o(g65236_sb) );
na03f02 TIMEBOOST_cell_53141 ( .a(n_5230), .b(n_3370), .c(n_2849), .o(TIMEBOOST_net_16788) );
na04f04 TIMEBOOST_cell_67928 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q), .b(FE_OFN2212_n_8407), .c(n_2184), .d(g61991_sb), .o(n_7913) );
in01f01 g65237_u0 ( .a(FE_OFN785_n_2678), .o(g65237_sb) );
in01f10 TIMEBOOST_cell_25263 ( .a(TIMEBOOST_net_6735), .o(n_16748) );
na03f02 TIMEBOOST_cell_66497 ( .a(TIMEBOOST_net_17118), .b(FE_OFN1312_n_6624), .c(g62547_sb), .o(n_6473) );
na02m02 TIMEBOOST_cell_53065 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(n_5769), .o(TIMEBOOST_net_16750) );
in01m01 g65238_u0 ( .a(FE_OFN789_n_2678), .o(g65238_sb) );
in01f08 TIMEBOOST_cell_25264 ( .a(TIMEBOOST_net_6736), .o(TIMEBOOST_net_6735) );
in01s01 g65240_u0 ( .a(FE_OFN786_n_2678), .o(g65240_sb) );
na02m01 TIMEBOOST_cell_68330 ( .a(n_4669), .b(n_12), .o(TIMEBOOST_net_21373) );
na03m06 TIMEBOOST_cell_69738 ( .a(g65362_sb), .b(FE_OFN1677_n_4655), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q), .o(TIMEBOOST_net_22077) );
in01f01 g65241_u0 ( .a(FE_OFN789_n_2678), .o(g65241_sb) );
na02s01 TIMEBOOST_cell_45595 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q), .o(TIMEBOOST_net_13692) );
na02s02 TIMEBOOST_cell_48032 ( .a(TIMEBOOST_net_14233), .b(g58024_sb), .o(TIMEBOOST_net_10379) );
in01f02 g65242_u0 ( .a(FE_OFN789_n_2678), .o(g65242_sb) );
na02m01 TIMEBOOST_cell_52833 ( .a(pci_target_unit_fifos_pciw_addr_data_in_150), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q), .o(TIMEBOOST_net_16634) );
in01f02 g65243_u0 ( .a(FE_OFN784_n_2678), .o(g65243_sb) );
na02s01 TIMEBOOST_cell_53029 ( .a(configuration_pci_err_data_530), .b(wbm_dat_o_29_), .o(TIMEBOOST_net_16732) );
in01f01 g65244_u0 ( .a(FE_OFN785_n_2678), .o(g65244_sb) );
na02s01 TIMEBOOST_cell_63009 ( .a(TIMEBOOST_net_20451), .b(g57968_sb), .o(TIMEBOOST_net_16595) );
na03m04 TIMEBOOST_cell_72484 ( .a(n_3792), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q), .c(TIMEBOOST_net_21533), .o(TIMEBOOST_net_17512) );
na04m10 TIMEBOOST_cell_67513 ( .a(g58017_sb), .b(FE_OFN262_n_9851), .c(FE_OFN527_n_9899), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q), .o(n_9775) );
in01f01 g65245_u0 ( .a(FE_OFN789_n_2678), .o(g65245_sb) );
na04f04 TIMEBOOST_cell_24197 ( .a(n_9097), .b(g57169_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q), .d(FE_OFN1416_n_8567), .o(n_10455) );
na02f02 TIMEBOOST_cell_70684 ( .a(TIMEBOOST_net_8322), .b(FE_OFN1120_g64577_p), .o(TIMEBOOST_net_22550) );
in01f01 g65246_u0 ( .a(FE_OFN785_n_2678), .o(g65246_sb) );
na02f02 TIMEBOOST_cell_70613 ( .a(TIMEBOOST_net_22514), .b(g63102_sb), .o(n_5050) );
in01f01 g65247_u0 ( .a(FE_OFN785_n_2678), .o(g65247_sb) );
na04f04 TIMEBOOST_cell_24199 ( .a(n_9745), .b(g57180_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q), .d(FE_OFN1406_n_8567), .o(n_11575) );
na02m20 TIMEBOOST_cell_53391 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q), .o(TIMEBOOST_net_16913) );
in01f01 g65248_u0 ( .a(FE_OFN785_n_2678), .o(g65248_sb) );
na04f04 TIMEBOOST_cell_24200 ( .a(n_9093), .b(g57188_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q), .d(FE_OFN1389_n_8567), .o(n_10449) );
na02m01 TIMEBOOST_cell_69800 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q), .o(TIMEBOOST_net_22108) );
in01f01 g65249_u0 ( .a(FE_OFN784_n_2678), .o(g65249_sb) );
na04f04 TIMEBOOST_cell_24201 ( .a(n_1465), .b(g58620_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .d(FE_OFN1369_n_8567), .o(n_9182) );
na03m02 TIMEBOOST_cell_68856 ( .a(g65049_sb), .b(n_4470), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q), .o(TIMEBOOST_net_21636) );
na02s01 TIMEBOOST_cell_45811 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q), .o(TIMEBOOST_net_13800) );
in01f02 g65250_u0 ( .a(FE_OFN784_n_2678), .o(g65250_sb) );
na02s01 TIMEBOOST_cell_31013 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_25__Q), .b(FE_OFN229_n_9120), .o(TIMEBOOST_net_9611) );
na02f02 TIMEBOOST_cell_40419 ( .a(TIMEBOOST_net_11821), .b(g59109_sb), .o(n_8709) );
in01m02 g65251_u0 ( .a(FE_OFN923_n_4740), .o(g65251_sb) );
na02s01 TIMEBOOST_cell_49299 ( .a(FE_OFN533_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q), .o(TIMEBOOST_net_14867) );
na02m10 TIMEBOOST_cell_51677 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q), .o(TIMEBOOST_net_16056) );
na02m02 TIMEBOOST_cell_49452 ( .a(TIMEBOOST_net_14943), .b(g58071_db), .o(TIMEBOOST_net_9559) );
in01s01 g65252_u0 ( .a(FE_OFN1046_n_16657), .o(g65252_sb) );
in01s01 TIMEBOOST_cell_35489 ( .a(TIMEBOOST_net_10080), .o(TIMEBOOST_net_10079) );
na02m06 TIMEBOOST_cell_72340 ( .a(TIMEBOOST_net_20765), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q), .o(TIMEBOOST_net_23378) );
na02s01 TIMEBOOST_cell_48222 ( .a(TIMEBOOST_net_14328), .b(g64225_sb), .o(n_4517) );
ao12f01 g65253_u0 ( .a(n_2469), .b(n_2468), .c(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_2979) );
no02s01 g65254_u0 ( .a(conf_wb_err_addr_in_945), .b(n_568), .o(g65254_p) );
ao12s01 g65254_u1 ( .a(g65254_p), .b(conf_wb_err_addr_in_945), .c(n_568), .o(n_1673) );
no02s01 g65255_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q), .b(n_1224), .o(g65255_p) );
ao12s01 g65255_u1 ( .a(g65255_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q), .c(n_1224), .o(n_2269) );
na02m06 TIMEBOOST_cell_68468 ( .a(g64806_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q), .o(TIMEBOOST_net_21442) );
no02m04 g65257_u0 ( .a(n_1674), .b(wbm_adr_o_4_), .o(g65257_p) );
ao12m02 g65257_u1 ( .a(g65257_p), .b(wbm_adr_o_4_), .c(n_1674), .o(n_1675) );
no02f01 g65258_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .b(n_1418), .o(g65258_p) );
ao12f01 g65258_u1 ( .a(g65258_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .c(n_1418), .o(n_1678) );
no02f01 g65259_u0 ( .a(n_2225), .b(wbu_addr_in_256), .o(g65259_p) );
ao12f01 g65259_u1 ( .a(g65259_p), .b(wbu_addr_in_256), .c(n_2225), .o(n_2226) );
no02s01 g65260_u0 ( .a(n_1679), .b(wbu_addr_in_253), .o(g65260_p) );
ao12s01 g65260_u1 ( .a(g65260_p), .b(wbu_addr_in_253), .c(n_1679), .o(n_1680) );
no02m06 g65261_u0 ( .a(n_1985), .b(wbm_adr_o_7_), .o(g65261_p) );
ao12m02 g65261_u1 ( .a(g65261_p), .b(wbm_adr_o_7_), .c(n_1985), .o(n_2224) );
in01f01 g65262_u0 ( .a(FE_OFN1012_n_4734), .o(g65262_sb) );
na02s01 TIMEBOOST_cell_48891 ( .a(FE_OFN235_n_9834), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q), .o(TIMEBOOST_net_14663) );
na02m08 TIMEBOOST_cell_62458 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q), .b(TIMEBOOST_net_12332), .o(TIMEBOOST_net_20176) );
no02s01 g65263_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_2_), .b(n_733), .o(g65263_p) );
ao12s01 g65263_u1 ( .a(g65263_p), .b(pci_target_unit_del_sync_comp_cycle_count_2_), .c(n_733), .o(n_1424) );
no02m02 g65264_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_), .b(n_554), .o(g65264_p) );
ao12m02 g65264_u1 ( .a(g65264_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_), .c(n_554), .o(n_1423) );
no02f03 g65265_u0 ( .a(conf_wb_err_addr_in_948), .b(n_1561), .o(g65265_p) );
ao12f02 g65265_u1 ( .a(g65265_p), .b(conf_wb_err_addr_in_948), .c(n_1561), .o(n_2395) );
no02s01 g65266_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .b(n_566), .o(g65266_p) );
ao12s01 g65266_u1 ( .a(g65266_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .c(n_566), .o(n_1422) );
no02f01 g65267_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .b(n_1215), .o(g65267_p) );
ao12f01 g65267_u1 ( .a(g65267_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .c(n_1215), .o(n_1421) );
in01s01 g65268_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(g65268_sb) );
na02s01 g65268_u1 ( .a(n_1109), .b(g65268_sb), .o(g65268_da) );
na02s01 g65268_u2 ( .a(n_8953), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(g65268_db) );
in01m01 g65269_u0 ( .a(FE_OCPN1839_n_1238), .o(g65269_sb) );
na04f04 TIMEBOOST_cell_73330 ( .a(n_4739), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q), .c(FE_OFN1119_g64577_p), .d(g62753_sb), .o(n_7134) );
na02m01 TIMEBOOST_cell_52713 ( .a(pci_target_unit_fifos_pciw_addr_data_in_135), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q), .o(TIMEBOOST_net_16574) );
in01f02 g65270_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .o(g65270_sb) );
na04f04 TIMEBOOST_cell_67684 ( .a(n_2797), .b(n_5230), .c(n_2820), .d(n_2819), .o(n_4167) );
na02s02 TIMEBOOST_cell_49436 ( .a(TIMEBOOST_net_14935), .b(g58070_sb), .o(TIMEBOOST_net_9581) );
in01m01 g65271_u0 ( .a(FE_OFN652_n_4508), .o(g65271_sb) );
na02m02 TIMEBOOST_cell_25396 ( .a(TIMEBOOST_net_6802), .b(n_4725), .o(TIMEBOOST_net_219) );
na03f10 TIMEBOOST_cell_37338 ( .a(n_2475), .b(n_2458), .c(n_2457), .o(TIMEBOOST_net_10281) );
in01m02 g65272_u0 ( .a(n_4677), .o(g65272_sb) );
na02s01 TIMEBOOST_cell_48719 ( .a(FE_OFN551_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q), .o(TIMEBOOST_net_14577) );
na02f02 TIMEBOOST_cell_18339 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q), .b(FE_OCPN1847_n_14981), .o(TIMEBOOST_net_5533) );
in01m04 g65273_u0 ( .a(FE_OFN643_n_4677), .o(g65273_sb) );
in01s01 TIMEBOOST_cell_45936 ( .a(TIMEBOOST_net_13897), .o(TIMEBOOST_net_13896) );
na02s01 TIMEBOOST_cell_52825 ( .a(pci_target_unit_fifos_pciw_addr_data_in_139), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q), .o(TIMEBOOST_net_16630) );
in01m02 g65274_u0 ( .a(FE_OFN1642_n_4671), .o(g65274_sb) );
na02s01 TIMEBOOST_cell_43657 ( .a(pci_target_unit_del_sync_addr_in_232), .b(parchk_pci_ad_reg_in_1233), .o(TIMEBOOST_net_12723) );
na02m10 TIMEBOOST_cell_31079 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .b(pci_target_unit_fifos_pcir_flush_in), .o(TIMEBOOST_net_9644) );
in01m02 g65275_u0 ( .a(FE_OFN643_n_4677), .o(g65275_sb) );
na02m01 TIMEBOOST_cell_48969 ( .a(TIMEBOOST_net_12678), .b(FE_OFN1055_n_4727), .o(TIMEBOOST_net_14702) );
in01m01 g65276_u0 ( .a(FE_OFN643_n_4677), .o(g65276_sb) );
na04f02 TIMEBOOST_cell_36827 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q), .b(FE_OFN1394_n_8567), .c(n_9499), .d(g57451_sb), .o(n_11283) );
na02s01 TIMEBOOST_cell_49453 ( .a(FE_OFN262_n_9851), .b(FE_RN_484_0), .o(TIMEBOOST_net_14944) );
na02m10 TIMEBOOST_cell_44031 ( .a(g58422_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q), .o(TIMEBOOST_net_12910) );
in01m02 g65277_u0 ( .a(FE_OFN642_n_4677), .o(g65277_sb) );
in01s01 TIMEBOOST_cell_67789 ( .a(TIMEBOOST_net_21216), .o(TIMEBOOST_net_21215) );
na04f02 TIMEBOOST_cell_68026 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q), .b(FE_OCPN1847_n_14981), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q), .d(g59112_sb), .o(n_8701) );
na02f01 TIMEBOOST_cell_68764 ( .a(n_2350), .b(pciu_pref_en_in_320), .o(TIMEBOOST_net_21590) );
in01m02 g65278_u0 ( .a(FE_OFN642_n_4677), .o(g65278_sb) );
na02s02 TIMEBOOST_cell_44033 ( .a(FE_OFN1789_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q), .o(TIMEBOOST_net_12911) );
na03m06 TIMEBOOST_cell_69730 ( .a(g65385_sb), .b(FE_OFN1677_n_4655), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q), .o(TIMEBOOST_net_22073) );
na03f02 TIMEBOOST_cell_42227 ( .a(n_3178), .b(g63550_sb), .c(TIMEBOOST_net_5550), .o(n_4607) );
in01m02 g65279_u0 ( .a(FE_OFN643_n_4677), .o(g65279_sb) );
na02m02 TIMEBOOST_cell_71979 ( .a(TIMEBOOST_net_23197), .b(g65329_sb), .o(TIMEBOOST_net_12545) );
na02f02 TIMEBOOST_cell_71525 ( .a(TIMEBOOST_net_22970), .b(FE_OFN1566_n_12502), .o(n_12507) );
in01m01 g65280_u0 ( .a(FE_OFN643_n_4677), .o(g65280_sb) );
na03f01 TIMEBOOST_cell_68218 ( .a(g57795_sb), .b(n_16070), .c(n_1083), .o(TIMEBOOST_net_21317) );
in01m01 g65281_u0 ( .a(FE_OFN643_n_4677), .o(g65281_sb) );
na02f01 TIMEBOOST_cell_44356 ( .a(TIMEBOOST_net_13072), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_11392) );
na02m02 TIMEBOOST_cell_44357 ( .a(n_4524), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q), .o(TIMEBOOST_net_13073) );
na02s01 TIMEBOOST_cell_44036 ( .a(TIMEBOOST_net_12912), .b(g58265_db), .o(n_9534) );
in01m02 g65282_u0 ( .a(FE_OFN644_n_4677), .o(g65282_sb) );
in01s02 TIMEBOOST_cell_45937 ( .a(TIMEBOOST_net_13898), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_101) );
in01m01 g65283_u0 ( .a(FE_OFN642_n_4677), .o(g65283_sb) );
in01m02 g65284_u0 ( .a(FE_OFN642_n_4677), .o(g65284_sb) );
na03f02 TIMEBOOST_cell_66494 ( .a(TIMEBOOST_net_13377), .b(n_6319), .c(g62348_sb), .o(n_6903) );
in01m04 g65285_u0 ( .a(FE_OFN644_n_4677), .o(g65285_sb) );
na03f02 TIMEBOOST_cell_73471 ( .a(TIMEBOOST_net_17416), .b(FE_OFN1206_n_6356), .c(g62712_sb), .o(n_6146) );
na03f02 TIMEBOOST_cell_66442 ( .a(TIMEBOOST_net_17132), .b(FE_OFN1317_n_6624), .c(g62481_sb), .o(n_6626) );
na02s01 TIMEBOOST_cell_37617 ( .a(TIMEBOOST_net_10420), .b(g58145_db), .o(n_9649) );
in01m06 g65286_u0 ( .a(n_4677), .o(g65286_sb) );
na02f02 TIMEBOOST_cell_51473 ( .a(n_14733), .b(n_8757), .o(TIMEBOOST_net_15954) );
na02m02 TIMEBOOST_cell_54098 ( .a(TIMEBOOST_net_17266), .b(FE_OFN215_n_9856), .o(n_9719) );
na02m02 TIMEBOOST_cell_52453 ( .a(wbm_adr_o_28_), .b(g59797_sb), .o(TIMEBOOST_net_16444) );
in01m01 g65287_u0 ( .a(FE_OFN643_n_4677), .o(g65287_sb) );
na02f01 TIMEBOOST_cell_68244 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_387), .o(TIMEBOOST_net_21330) );
in01m01 g65288_u0 ( .a(FE_OFN644_n_4677), .o(g65288_sb) );
na02m01 g65288_u2 ( .a(n_3739), .b(FE_OFN644_n_4677), .o(g65288_db) );
in01s01 TIMEBOOST_cell_73850 ( .a(n_7400), .o(TIMEBOOST_net_23415) );
in01m02 g65289_u0 ( .a(FE_OFN644_n_4677), .o(g65289_sb) );
na02s02 TIMEBOOST_cell_49455 ( .a(FE_OFN264_n_9849), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q), .o(TIMEBOOST_net_14945) );
na02m01 TIMEBOOST_cell_68932 ( .a(n_4645), .b(n_50), .o(TIMEBOOST_net_21674) );
na02f02 TIMEBOOST_cell_51516 ( .a(TIMEBOOST_net_15975), .b(n_16853), .o(n_4858) );
no03f06 TIMEBOOST_cell_67095 ( .a(FE_RN_805_0), .b(FE_RN_807_0), .c(FE_RN_806_0), .o(n_14273) );
na02s01 TIMEBOOST_cell_49269 ( .a(FE_OFN555_n_9864), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q), .o(TIMEBOOST_net_14852) );
in01m02 g65291_u0 ( .a(n_4677), .o(g65291_sb) );
na04f04 TIMEBOOST_cell_73426 ( .a(n_4406), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q), .c(FE_OFN1203_n_4090), .d(g62594_sb), .o(n_6364) );
na02s02 TIMEBOOST_cell_69157 ( .a(TIMEBOOST_net_21786), .b(FE_OFN1042_n_2037), .o(TIMEBOOST_net_16625) );
na03f02 TIMEBOOST_cell_73560 ( .a(TIMEBOOST_net_17077), .b(FE_OFN1230_n_6391), .c(g63000_sb), .o(n_5882) );
in01m01 g65292_u0 ( .a(FE_OFN642_n_4677), .o(g65292_sb) );
in01s01 TIMEBOOST_cell_73953 ( .a(TIMEBOOST_net_23517), .o(TIMEBOOST_net_23518) );
na03f02 TIMEBOOST_cell_73580 ( .a(TIMEBOOST_net_7616), .b(FE_OFN1085_n_13221), .c(TIMEBOOST_net_15683), .o(n_13490) );
na03f02 TIMEBOOST_cell_73526 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q), .b(n_4901), .c(n_6431), .o(TIMEBOOST_net_22815) );
in01m01 g65293_u0 ( .a(FE_OFN644_n_4677), .o(g65293_sb) );
na03m02 TIMEBOOST_cell_73172 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q), .b(g64319_sb), .c(g64319_db), .o(n_3857) );
na03m02 TIMEBOOST_cell_72636 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q), .c(TIMEBOOST_net_16208), .o(TIMEBOOST_net_17531) );
in01m01 g65294_u0 ( .a(FE_OFN636_n_4669), .o(g65294_sb) );
na02s01 TIMEBOOST_cell_43653 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q), .b(FE_OFN205_n_9140), .o(TIMEBOOST_net_12721) );
na03s02 TIMEBOOST_cell_73187 ( .a(TIMEBOOST_net_10046), .b(g62066_sb), .c(TIMEBOOST_net_5644), .o(n_7833) );
na04m02 TIMEBOOST_cell_73113 ( .a(TIMEBOOST_net_8271), .b(g65788_db), .c(g61807_sb), .d(TIMEBOOST_net_21051), .o(n_8180) );
in01m06 g65295_u0 ( .a(FE_OFN640_n_4669), .o(g65295_sb) );
na02s02 TIMEBOOST_cell_44600 ( .a(TIMEBOOST_net_13194), .b(g58297_sb), .o(n_9216) );
na02m01 TIMEBOOST_cell_49002 ( .a(TIMEBOOST_net_14718), .b(n_4672), .o(n_4358) );
na02s02 TIMEBOOST_cell_53556 ( .a(TIMEBOOST_net_16995), .b(g57994_sb), .o(TIMEBOOST_net_9388) );
in01m06 g65296_u0 ( .a(FE_OFN639_n_4669), .o(g65296_sb) );
na02m06 TIMEBOOST_cell_68858 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q), .b(n_4482), .o(TIMEBOOST_net_21637) );
in01s01 TIMEBOOST_cell_45893 ( .a(wbu_sel_in_313), .o(TIMEBOOST_net_13854) );
in01m01 g65297_u0 ( .a(FE_OFN639_n_4669), .o(g65297_sb) );
na02f01 TIMEBOOST_cell_70332 ( .a(TIMEBOOST_net_5267), .b(g62111_sb), .o(TIMEBOOST_net_22374) );
in01m01 g65298_u0 ( .a(FE_OFN640_n_4669), .o(g65298_sb) );
na03m02 TIMEBOOST_cell_72776 ( .a(n_4447), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q), .c(TIMEBOOST_net_12550), .o(TIMEBOOST_net_20972) );
na02f01 g65298_u2 ( .a(n_3744), .b(FE_OFN640_n_4669), .o(g65298_db) );
in01m02 g65299_u0 ( .a(FE_OFN640_n_4669), .o(g65299_sb) );
na03f02 TIMEBOOST_cell_66751 ( .a(TIMEBOOST_net_16832), .b(FE_OFN1306_n_13124), .c(g54349_sb), .o(n_13093) );
in01m01 g65300_u0 ( .a(FE_OFN640_n_4669), .o(g65300_sb) );
na03f02 TIMEBOOST_cell_72282 ( .a(TIMEBOOST_net_20994), .b(FE_OFN1670_n_9477), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q), .o(TIMEBOOST_net_23349) );
in01m02 g65301_u0 ( .a(FE_OFN640_n_4669), .o(g65301_sb) );
na04f04 TIMEBOOST_cell_24956 ( .a(n_16836), .b(n_10547), .c(n_16837), .d(n_9962), .o(n_12130) );
na02m02 TIMEBOOST_cell_68177 ( .a(TIMEBOOST_net_21296), .b(TIMEBOOST_net_14037), .o(TIMEBOOST_net_16804) );
na02s02 TIMEBOOST_cell_48720 ( .a(TIMEBOOST_net_14577), .b(TIMEBOOST_net_10516), .o(TIMEBOOST_net_9361) );
in01m04 g65302_u0 ( .a(FE_OFN639_n_4669), .o(g65302_sb) );
in01s01 TIMEBOOST_cell_72361 ( .a(TIMEBOOST_net_23393), .o(TIMEBOOST_net_23394) );
na03f02 TIMEBOOST_cell_34792 ( .a(TIMEBOOST_net_9556), .b(FE_OFN1409_n_8567), .c(g57167_sb), .o(n_11586) );
in01m02 g65303_u0 ( .a(FE_OFN642_n_4677), .o(g65303_sb) );
na02s02 TIMEBOOST_cell_44601 ( .a(FE_OFN201_n_9230), .b(g58446_sb), .o(TIMEBOOST_net_13195) );
na02m02 TIMEBOOST_cell_68837 ( .a(TIMEBOOST_net_21626), .b(TIMEBOOST_net_14276), .o(TIMEBOOST_net_17454) );
in01m02 g65304_u0 ( .a(FE_OFN639_n_4669), .o(g65304_sb) );
na04m02 TIMEBOOST_cell_67267 ( .a(n_3752), .b(g64986_sb), .c(g64986_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q), .o(TIMEBOOST_net_17102) );
na03f02 TIMEBOOST_cell_65883 ( .a(TIMEBOOST_net_14971), .b(g62757_sb), .c(g62757_db), .o(n_5474) );
na02s01 TIMEBOOST_cell_51565 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q), .o(TIMEBOOST_net_16000) );
in01m06 g65305_u0 ( .a(FE_OFN640_n_4669), .o(g65305_sb) );
in01s01 TIMEBOOST_cell_73936 ( .a(wbm_dat_i_19_), .o(TIMEBOOST_net_23501) );
in01m04 g65306_u0 ( .a(FE_OFN636_n_4669), .o(g65306_sb) );
na02s01 TIMEBOOST_cell_43785 ( .a(FE_OFN207_n_9865), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q), .o(TIMEBOOST_net_12787) );
na02s01 TIMEBOOST_cell_48877 ( .a(FE_OFN239_n_9832), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q), .o(TIMEBOOST_net_14656) );
na02f02 TIMEBOOST_cell_71091 ( .a(TIMEBOOST_net_22753), .b(g62670_sb), .o(n_6199) );
in01m01 g65307_u0 ( .a(FE_OFN640_n_4669), .o(g65307_sb) );
na02m02 TIMEBOOST_cell_50628 ( .a(TIMEBOOST_net_15531), .b(g62456_sb), .o(n_6684) );
na02m02 TIMEBOOST_cell_70155 ( .a(TIMEBOOST_net_22285), .b(g64086_sb), .o(n_4069) );
na03f02 TIMEBOOST_cell_73644 ( .a(TIMEBOOST_net_17468), .b(FE_OFN1250_n_4093), .c(g62957_sb), .o(n_5967) );
in01m02 g65308_u0 ( .a(FE_OFN636_n_4669), .o(g65308_sb) );
na02s01 TIMEBOOST_cell_43777 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q), .b(FE_OFN239_n_9832), .o(TIMEBOOST_net_12783) );
na03s01 TIMEBOOST_cell_64741 ( .a(pci_target_unit_del_sync_addr_in_218), .b(g66406_sb), .c(g66428_db), .o(n_2498) );
na02s01 TIMEBOOST_cell_43153 ( .a(FE_OFN243_n_9116), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q), .o(TIMEBOOST_net_12471) );
in01m01 g65309_u0 ( .a(n_4669), .o(g65309_sb) );
na02m02 g65309_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q), .b(g65309_sb), .o(g65309_da) );
in01m01 g65310_u0 ( .a(n_4669), .o(g65310_sb) );
na04m04 TIMEBOOST_cell_67318 ( .a(g64803_sb), .b(n_4493), .c(g64803_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q), .o(TIMEBOOST_net_17438) );
na03f02 TIMEBOOST_cell_66694 ( .a(TIMEBOOST_net_17150), .b(FE_OFN1313_n_6624), .c(g62562_sb), .o(n_6435) );
in01m01 g65311_u0 ( .a(FE_OFN636_n_4669), .o(g65311_sb) );
na02m02 TIMEBOOST_cell_54376 ( .a(TIMEBOOST_net_17405), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_15414) );
na03f02 TIMEBOOST_cell_66832 ( .a(TIMEBOOST_net_13487), .b(n_14839), .c(g59797_db), .o(TIMEBOOST_net_16007) );
in01s01 g65312_u0 ( .a(FE_OFN636_n_4669), .o(g65312_sb) );
na02s02 TIMEBOOST_cell_44602 ( .a(TIMEBOOST_net_13195), .b(g58446_db), .o(n_9199) );
na02f02 TIMEBOOST_cell_70253 ( .a(TIMEBOOST_net_22334), .b(g62780_sb), .o(n_5431) );
na02s01 TIMEBOOST_cell_51567 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q), .o(TIMEBOOST_net_16001) );
in01m02 g65313_u0 ( .a(FE_OFN1642_n_4671), .o(g65313_sb) );
na02s01 TIMEBOOST_cell_45253 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q), .o(TIMEBOOST_net_13521) );
na02s01 TIMEBOOST_cell_43761 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q), .b(FE_OFN239_n_9832), .o(TIMEBOOST_net_12775) );
in01m01 g65314_u0 ( .a(FE_OFN1643_n_4671), .o(g65314_sb) );
na04s02 TIMEBOOST_cell_46579 ( .a(TIMEBOOST_net_10785), .b(g65833_sb), .c(g61743_sb), .d(g61898_db), .o(n_8030) );
na02f02 TIMEBOOST_cell_71012 ( .a(TIMEBOOST_net_17426), .b(FE_OFN1202_n_4090), .o(TIMEBOOST_net_22714) );
in01m02 g65315_u0 ( .a(FE_OFN1642_n_4671), .o(g65315_sb) );
na03m06 TIMEBOOST_cell_72985 ( .a(FE_OFN1628_n_4438), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q), .c(g64991_sb), .o(TIMEBOOST_net_14718) );
na02m01 TIMEBOOST_cell_69926 ( .a(n_4645), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q), .o(TIMEBOOST_net_22171) );
in01s01 TIMEBOOST_cell_73954 ( .a(wbm_dat_i_27_), .o(TIMEBOOST_net_23519) );
in01m06 g65316_u0 ( .a(FE_OFN1642_n_4671), .o(g65316_sb) );
na02m02 TIMEBOOST_cell_68121 ( .a(TIMEBOOST_net_21268), .b(g61880_sb), .o(TIMEBOOST_net_17287) );
na03m02 TIMEBOOST_cell_65449 ( .a(TIMEBOOST_net_10760), .b(TIMEBOOST_net_9820), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q), .o(TIMEBOOST_net_20978) );
in01m01 g65317_u0 ( .a(FE_OFN1642_n_4671), .o(g65317_sb) );
na04m02 TIMEBOOST_cell_67271 ( .a(n_3749), .b(g64929_sb), .c(g64929_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q), .o(TIMEBOOST_net_17130) );
na02m01 g64963_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q), .b(FE_OFN618_n_4490), .o(g64963_db) );
in01m02 g65318_u0 ( .a(FE_OFN1642_n_4671), .o(g65318_sb) );
na04f02 TIMEBOOST_cell_68027 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q), .b(FE_OCPN1847_n_14981), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q), .d(g59111_sb), .o(n_8697) );
na02s01 TIMEBOOST_cell_52235 ( .a(FE_OFN211_n_9858), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q), .o(TIMEBOOST_net_16335) );
na03f02 TIMEBOOST_cell_73266 ( .a(TIMEBOOST_net_22199), .b(FE_OFN2081_n_8176), .c(g61910_sb), .o(n_8001) );
in01m04 g65319_u0 ( .a(FE_OFN1643_n_4671), .o(g65319_sb) );
na03f02 TIMEBOOST_cell_32959 ( .a(TIMEBOOST_net_8725), .b(n_5633), .c(g62090_sb), .o(n_5617) );
na02f02 TIMEBOOST_cell_68647 ( .a(TIMEBOOST_net_21531), .b(TIMEBOOST_net_20198), .o(TIMEBOOST_net_17372) );
in01s01 TIMEBOOST_cell_45943 ( .a(wbu_sel_in_312), .o(TIMEBOOST_net_13904) );
in01m06 g65320_u0 ( .a(FE_OFN1644_n_4671), .o(g65320_sb) );
na03f01 TIMEBOOST_cell_68122 ( .a(TIMEBOOST_net_13995), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q), .o(TIMEBOOST_net_21269) );
na03s02 TIMEBOOST_cell_72735 ( .a(TIMEBOOST_net_13895), .b(g65749_sb), .c(g65749_db), .o(n_1924) );
in01s01 TIMEBOOST_cell_45971 ( .a(pci_target_unit_fifos_pcir_data_in_187), .o(TIMEBOOST_net_13932) );
in01m01 g65321_u0 ( .a(FE_OFN1642_n_4671), .o(g65321_sb) );
na02m02 TIMEBOOST_cell_71882 ( .a(TIMEBOOST_net_20214), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q), .o(TIMEBOOST_net_23149) );
in01s01 TIMEBOOST_cell_45894 ( .a(TIMEBOOST_net_13854), .o(TIMEBOOST_net_13855) );
na02m02 TIMEBOOST_cell_68203 ( .a(TIMEBOOST_net_21309), .b(g56934_sb), .o(TIMEBOOST_net_14192) );
in01m02 g65322_u0 ( .a(FE_OFN1640_n_4671), .o(g65322_sb) );
na02s01 TIMEBOOST_cell_54101 ( .a(FE_OFN239_n_9832), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q), .o(TIMEBOOST_net_17268) );
in01s01 TIMEBOOST_cell_73913 ( .a(TIMEBOOST_net_23477), .o(TIMEBOOST_net_23478) );
na03f02 TIMEBOOST_cell_66160 ( .a(TIMEBOOST_net_20948), .b(FE_OFN1180_n_3476), .c(g60622_sb), .o(n_4832) );
in01m01 g65323_u0 ( .a(FE_OFN1640_n_4671), .o(g65323_sb) );
na04f04 TIMEBOOST_cell_67471 ( .a(n_4374), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q), .c(FE_OFN1250_n_4093), .d(g62352_sb), .o(n_6897) );
na02m02 TIMEBOOST_cell_49664 ( .a(TIMEBOOST_net_15049), .b(g61737_sb), .o(n_8344) );
in01m02 g65324_u0 ( .a(FE_OFN1645_n_4671), .o(g65324_sb) );
na02m02 g65324_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q), .b(g65324_sb), .o(g65324_da) );
na03f02 TIMEBOOST_cell_73267 ( .a(TIMEBOOST_net_12961), .b(g63141_sb), .c(g63141_db), .o(n_4965) );
in01f01 g65325_u0 ( .a(n_4671), .o(g65325_sb) );
na02m02 g65325_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q), .b(g65325_sb), .o(g65325_da) );
na03s02 TIMEBOOST_cell_289 ( .a(n_1565), .b(g61732_sb), .c(g61938_db), .o(n_7947) );
na04s02 TIMEBOOST_cell_32479 ( .a(FE_OFN209_n_9126), .b(g58141_sb), .c(g58141_db), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q), .o(TIMEBOOST_net_9551) );
in01m01 g65326_u0 ( .a(FE_OFN1644_n_4671), .o(g65326_sb) );
na02s01 TIMEBOOST_cell_43817 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q), .b(FE_OFN211_n_9858), .o(TIMEBOOST_net_12803) );
in01s01 TIMEBOOST_cell_45984 ( .a(TIMEBOOST_net_13944), .o(TIMEBOOST_net_13945) );
na03m02 TIMEBOOST_cell_72736 ( .a(g64329_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q), .c(TIMEBOOST_net_14301), .o(TIMEBOOST_net_13066) );
in01m01 g65327_u0 ( .a(FE_OFN654_n_4508), .o(g65327_sb) );
na04f10 TIMEBOOST_cell_31946 ( .a(n_1698), .b(n_2648), .c(n_8511), .d(n_3030), .o(n_2380) );
na02m02 TIMEBOOST_cell_51330 ( .a(TIMEBOOST_net_15882), .b(g62779_sb), .o(n_5433) );
in01s01 TIMEBOOST_cell_63561 ( .a(TIMEBOOST_net_20741), .o(TIMEBOOST_net_20740) );
in01m01 g65328_u0 ( .a(FE_OFN652_n_4508), .o(g65328_sb) );
na02f02 TIMEBOOST_cell_72157 ( .a(TIMEBOOST_net_23286), .b(TIMEBOOST_net_14754), .o(TIMEBOOST_net_17329) );
in01s01 TIMEBOOST_cell_73972 ( .a(wbm_dat_i_6_), .o(TIMEBOOST_net_23537) );
in01m01 g65329_u0 ( .a(FE_OFN653_n_4508), .o(g65329_sb) );
na03m02 TIMEBOOST_cell_72717 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q), .b(g63565_sb), .c(g63565_db), .o(TIMEBOOST_net_14946) );
na02m10 TIMEBOOST_cell_45553 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q), .o(TIMEBOOST_net_13671) );
in01m02 g65330_u0 ( .a(FE_OFN654_n_4508), .o(g65330_sb) );
na02s01 TIMEBOOST_cell_43665 ( .a(pci_target_unit_del_sync_addr_in_216), .b(parchk_pci_ad_reg_in_1217), .o(TIMEBOOST_net_12727) );
na02s01 TIMEBOOST_cell_45255 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q), .o(TIMEBOOST_net_13522) );
na02m08 TIMEBOOST_cell_52869 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q), .b(wbs_dat_i_26_), .o(TIMEBOOST_net_16652) );
in01m01 g65331_u0 ( .a(FE_OFN654_n_4508), .o(g65331_sb) );
na03m04 TIMEBOOST_cell_72491 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q), .b(n_3755), .c(TIMEBOOST_net_22077), .o(TIMEBOOST_net_17077) );
in01m01 g65332_u0 ( .a(FE_OFN654_n_4508), .o(g65332_sb) );
na02m02 g65332_u2 ( .a(n_3774), .b(FE_OFN654_n_4508), .o(g65332_db) );
na02m02 TIMEBOOST_cell_69087 ( .a(TIMEBOOST_net_21751), .b(g65058_db), .o(TIMEBOOST_net_17406) );
in01m01 g65333_u0 ( .a(FE_OFN651_n_4508), .o(g65333_sb) );
na02s01 TIMEBOOST_cell_43673 ( .a(pci_target_unit_del_sync_addr_in_224), .b(parchk_pci_ad_reg_in_1225), .o(TIMEBOOST_net_12731) );
na03m02 TIMEBOOST_cell_72737 ( .a(g64992_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q), .c(TIMEBOOST_net_16196), .o(TIMEBOOST_net_17019) );
in01m01 g65334_u0 ( .a(FE_OFN653_n_4508), .o(g65334_sb) );
na02s02 TIMEBOOST_cell_52236 ( .a(TIMEBOOST_net_16335), .b(FE_OFN1687_n_9528), .o(TIMEBOOST_net_11525) );
na02m02 TIMEBOOST_cell_63987 ( .a(TIMEBOOST_net_20979), .b(FE_OFN1279_n_4097), .o(TIMEBOOST_net_15473) );
na02s01 TIMEBOOST_cell_43661 ( .a(pci_target_unit_del_sync_addr_in_226), .b(parchk_pci_ad_reg_in_1227), .o(TIMEBOOST_net_12725) );
in01m01 g65335_u0 ( .a(FE_OFN653_n_4508), .o(g65335_sb) );
na02m01 g65335_u2 ( .a(n_3785), .b(FE_OFN653_n_4508), .o(g65335_db) );
na03f02 TIMEBOOST_cell_66954 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_16505), .c(FE_OFN1568_n_11027), .o(n_12644) );
in01m04 g65336_u0 ( .a(FE_OFN654_n_4508), .o(g65336_sb) );
na02f01 TIMEBOOST_cell_31115 ( .a(n_3030), .b(g67051_sb), .o(TIMEBOOST_net_9662) );
in01m01 g65337_u0 ( .a(FE_OFN652_n_4508), .o(g65337_sb) );
na02m04 TIMEBOOST_cell_43685 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q), .b(FE_OFN685_n_4417), .o(TIMEBOOST_net_12737) );
na02f01 TIMEBOOST_cell_31117 ( .a(g67051_sb), .b(parchk_pci_trdy_reg_in), .o(TIMEBOOST_net_9663) );
na04f04 TIMEBOOST_cell_73645 ( .a(n_1881), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q), .c(FE_OFN706_n_8119), .d(g61905_sb), .o(n_8012) );
in01m01 g65338_u0 ( .a(FE_OFN654_n_4508), .o(g65338_sb) );
na02s02 TIMEBOOST_cell_51401 ( .a(g58240_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q), .o(TIMEBOOST_net_15918) );
na02f02 g65338_u2 ( .a(n_3770), .b(FE_OFN654_n_4508), .o(g65338_db) );
in01s01 TIMEBOOST_cell_73901 ( .a(TIMEBOOST_net_23465), .o(TIMEBOOST_net_23466) );
in01m04 g65339_u0 ( .a(FE_OFN644_n_4677), .o(g65339_sb) );
na02f02 TIMEBOOST_cell_71397 ( .a(TIMEBOOST_net_22906), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_16642) );
in01m01 g65340_u0 ( .a(FE_OFN651_n_4508), .o(g65340_sb) );
na02f02 TIMEBOOST_cell_49391 ( .a(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74), .b(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(TIMEBOOST_net_14913) );
in01s02 TIMEBOOST_cell_67097 ( .a(TIMEBOOST_net_21131), .o(TIMEBOOST_net_21130) );
in01m04 g65341_u0 ( .a(FE_OFN651_n_4508), .o(g65341_sb) );
na03f06 TIMEBOOST_cell_73490 ( .a(n_3290), .b(pciu_bar0_in), .c(n_2905), .o(TIMEBOOST_net_8004) );
na04f04 TIMEBOOST_cell_24562 ( .a(n_9229), .b(g57095_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q), .d(FE_OFN1417_n_8567), .o(n_10843) );
in01m02 g65342_u0 ( .a(FE_OFN652_n_4508), .o(g65342_sb) );
na02f01 TIMEBOOST_cell_49690 ( .a(TIMEBOOST_net_15062), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_13166) );
in01m02 g65343_u0 ( .a(FE_OFN652_n_4508), .o(g65343_sb) );
na02f02 TIMEBOOST_cell_50978 ( .a(TIMEBOOST_net_15706), .b(g62958_sb), .o(n_5966) );
na02m01 TIMEBOOST_cell_62644 ( .a(n_3739), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q), .o(TIMEBOOST_net_20269) );
na03f02 TIMEBOOST_cell_66611 ( .a(TIMEBOOST_net_17103), .b(FE_OFN1323_n_6436), .c(g62561_sb), .o(n_6438) );
na02f02 TIMEBOOST_cell_38855 ( .a(TIMEBOOST_net_11039), .b(g61785_sb), .o(n_8234) );
in01m02 g65345_u0 ( .a(FE_OFN1643_n_4671), .o(g65345_sb) );
na03m02 TIMEBOOST_cell_72587 ( .a(TIMEBOOST_net_21431), .b(g64790_sb), .c(TIMEBOOST_net_21639), .o(TIMEBOOST_net_17435) );
in01s01 TIMEBOOST_cell_73955 ( .a(TIMEBOOST_net_23519), .o(TIMEBOOST_net_23520) );
in01m02 g65346_u0 ( .a(FE_OFN640_n_4669), .o(g65346_sb) );
na03f02 TIMEBOOST_cell_24958 ( .a(n_10634), .b(FE_RN_474_0), .c(n_12574), .o(n_12836) );
in01m01 g65347_u0 ( .a(FE_OFN1676_n_4655), .o(g65347_sb) );
na02m04 TIMEBOOST_cell_62620 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_138), .o(TIMEBOOST_net_20257) );
na03m02 TIMEBOOST_cell_65095 ( .a(n_3770), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q), .c(FE_OFN1642_n_4671), .o(TIMEBOOST_net_16249) );
in01m01 g65348_u0 ( .a(FE_OFN1677_n_4655), .o(g65348_sb) );
na02s02 TIMEBOOST_cell_52319 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q), .b(g58299_sb), .o(TIMEBOOST_net_16377) );
in01s01 TIMEBOOST_cell_67714 ( .a(TIMEBOOST_net_21140), .o(TIMEBOOST_net_21141) );
in01m02 g65349_u0 ( .a(FE_OFN1679_n_4655), .o(g65349_sb) );
na02f02 TIMEBOOST_cell_71399 ( .a(TIMEBOOST_net_22907), .b(FE_OFN709_n_8232), .o(TIMEBOOST_net_16643) );
na02f06 TIMEBOOST_cell_48693 ( .a(FE_RN_47_0), .b(n_2409), .o(TIMEBOOST_net_14564) );
in01m06 g65350_u0 ( .a(FE_OFN1680_n_4655), .o(g65350_sb) );
na03f02 TIMEBOOST_cell_72913 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q), .b(g64282_sb), .c(TIMEBOOST_net_22098), .o(TIMEBOOST_net_20627) );
in01m04 g65351_u0 ( .a(FE_OFN1677_n_4655), .o(g65351_sb) );
in01s01 TIMEBOOST_cell_63551 ( .a(TIMEBOOST_net_20731), .o(TIMEBOOST_net_20730) );
na03f02 TIMEBOOST_cell_66520 ( .a(TIMEBOOST_net_16809), .b(FE_OFN1333_n_13547), .c(g53929_sb), .o(n_13516) );
in01m01 g65352_u0 ( .a(FE_OFN1677_n_4655), .o(g65352_sb) );
na02f02 TIMEBOOST_cell_70666 ( .a(TIMEBOOST_net_13055), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_22541) );
na02m02 TIMEBOOST_cell_71927 ( .a(TIMEBOOST_net_23171), .b(g64142_sb), .o(n_4523) );
in01m01 g65353_u0 ( .a(FE_OFN1677_n_4655), .o(g65353_sb) );
na02f02 TIMEBOOST_cell_70665 ( .a(TIMEBOOST_net_22540), .b(g62732_sb), .o(n_5515) );
na03m02 TIMEBOOST_cell_72605 ( .a(TIMEBOOST_net_21472), .b(FE_OFN1643_n_4671), .c(TIMEBOOST_net_21723), .o(TIMEBOOST_net_17022) );
na03s01 TIMEBOOST_cell_46921 ( .a(FE_OFN201_n_9230), .b(g57891_sb), .c(g57891_db), .o(n_9233) );
in01m01 g65354_u0 ( .a(FE_OFN1679_n_4655), .o(g65354_sb) );
in01s01 TIMEBOOST_cell_63545 ( .a(TIMEBOOST_net_20725), .o(TIMEBOOST_net_20724) );
in01m08 g65355_u0 ( .a(FE_OFN1676_n_4655), .o(g65355_sb) );
in01s01 TIMEBOOST_cell_45895 ( .a(TIMEBOOST_net_13856), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_81) );
in01m01 g65356_u0 ( .a(FE_OFN1680_n_4655), .o(g65356_sb) );
na02s01 TIMEBOOST_cell_63008 ( .a(FE_OFN237_n_9118), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q), .o(TIMEBOOST_net_20451) );
in01m06 g65357_u0 ( .a(FE_OFN1678_n_4655), .o(g65357_sb) );
na04f02 TIMEBOOST_cell_68020 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in), .b(g54172_sb), .c(g53946_da), .d(TIMEBOOST_net_645), .o(n_13497) );
in01m01 g65358_u0 ( .a(FE_OFN1680_n_4655), .o(g65358_sb) );
na02s01 TIMEBOOST_cell_49470 ( .a(TIMEBOOST_net_14952), .b(FE_OFN1650_n_9428), .o(TIMEBOOST_net_11175) );
na02s03 TIMEBOOST_cell_42887 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q), .o(TIMEBOOST_net_12338) );
in01m01 g65359_u0 ( .a(FE_OFN1676_n_4655), .o(g65359_sb) );
na02s02 TIMEBOOST_cell_49471 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q), .o(TIMEBOOST_net_14953) );
in01s01 TIMEBOOST_cell_67731 ( .a(pci_target_unit_fifos_pcir_data_in_175), .o(TIMEBOOST_net_21158) );
na02m06 TIMEBOOST_cell_42859 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_145), .o(TIMEBOOST_net_12324) );
in01m01 g65360_u0 ( .a(FE_OFN1678_n_4655), .o(g65360_sb) );
in01s01 TIMEBOOST_cell_63544 ( .a(TIMEBOOST_net_20724), .o(TIMEBOOST_net_10060) );
na03m04 TIMEBOOST_cell_72498 ( .a(n_3744), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q), .c(TIMEBOOST_net_22076), .o(TIMEBOOST_net_17076) );
na02m02 TIMEBOOST_cell_63983 ( .a(TIMEBOOST_net_20977), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_15404) );
in01m02 g65361_u0 ( .a(FE_OFN1676_n_4655), .o(g65361_sb) );
na02s01 TIMEBOOST_cell_42801 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q), .o(TIMEBOOST_net_12295) );
in01s01 TIMEBOOST_cell_67791 ( .a(TIMEBOOST_net_21218), .o(TIMEBOOST_net_21213) );
in01m04 g65362_u0 ( .a(FE_OFN1677_n_4655), .o(g65362_sb) );
na04m06 TIMEBOOST_cell_67426 ( .a(g58043_db), .b(FE_OFN211_n_9858), .c(g58043_sb), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q), .o(TIMEBOOST_net_16847) );
na02m02 TIMEBOOST_cell_69045 ( .a(TIMEBOOST_net_21730), .b(TIMEBOOST_net_20245), .o(TIMEBOOST_net_17448) );
in01m02 g65363_u0 ( .a(FE_OFN1676_n_4655), .o(g65363_sb) );
in01s01 TIMEBOOST_cell_73851 ( .a(TIMEBOOST_net_23415), .o(TIMEBOOST_net_23416) );
na02s02 TIMEBOOST_cell_38441 ( .a(TIMEBOOST_net_10832), .b(g57919_db), .o(n_9134) );
na02m01 TIMEBOOST_cell_47581 ( .a(n_8831), .b(g58770_sb), .o(TIMEBOOST_net_14008) );
in01m01 g65364_u0 ( .a(FE_OFN1676_n_4655), .o(g65364_sb) );
na02m02 TIMEBOOST_cell_68955 ( .a(TIMEBOOST_net_21685), .b(g65331_sb), .o(n_4265) );
in01m01 g65365_u0 ( .a(FE_OFN1676_n_4655), .o(g65365_sb) );
na03f02 TIMEBOOST_cell_73787 ( .a(TIMEBOOST_net_16540), .b(FE_OFN1601_n_13995), .c(FE_OFN1605_n_13997), .o(g53310_p) );
na02f02 TIMEBOOST_cell_49658 ( .a(TIMEBOOST_net_15046), .b(g61860_sb), .o(n_8118) );
na03s02 TIMEBOOST_cell_67906 ( .a(TIMEBOOST_net_7103), .b(FE_OFN775_n_15366), .c(g65893_sb), .o(n_2585) );
in01m02 g65366_u0 ( .a(FE_OFN1643_n_4671), .o(g65366_sb) );
na02m20 TIMEBOOST_cell_43677 ( .a(pci_target_unit_fifos_pciw_addr_data_in_130), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q), .o(TIMEBOOST_net_12733) );
na02f02 TIMEBOOST_cell_70165 ( .a(TIMEBOOST_net_22290), .b(g64222_sb), .o(n_3947) );
in01m01 g65367_u0 ( .a(FE_OFN1642_n_4671), .o(g65367_sb) );
na04f04 TIMEBOOST_cell_24564 ( .a(n_9199), .b(g57596_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q), .d(FE_OFN1402_n_8567), .o(n_10797) );
in01m02 g65368_u0 ( .a(FE_OFN644_n_4677), .o(g65368_sb) );
na03f02 TIMEBOOST_cell_65946 ( .a(g62108_sb), .b(FE_OFN1174_n_5592), .c(TIMEBOOST_net_16409), .o(n_5591) );
na02m02 TIMEBOOST_cell_68805 ( .a(TIMEBOOST_net_21610), .b(g64360_sb), .o(TIMEBOOST_net_13057) );
na02s01 TIMEBOOST_cell_38305 ( .a(TIMEBOOST_net_10764), .b(g52479_sb), .o(TIMEBOOST_net_745) );
in01m01 g65369_u0 ( .a(FE_OFN1640_n_4671), .o(g65369_sb) );
na03s02 TIMEBOOST_cell_22337 ( .a(FE_OFN254_n_9825), .b(g58140_sb), .c(g58168_db), .o(n_9623) );
in01m01 g65370_u0 ( .a(FE_OFN1644_n_4671), .o(g65370_sb) );
na03f02 TIMEBOOST_cell_73427 ( .a(TIMEBOOST_net_17362), .b(FE_OFN1282_n_4097), .c(g62360_sb), .o(n_6878) );
na02m02 TIMEBOOST_cell_64170 ( .a(wbm_adr_o_27_), .b(g60679_sb), .o(TIMEBOOST_net_21071) );
in01s01 TIMEBOOST_cell_45973 ( .a(TIMEBOOST_net_13933), .o(TIMEBOOST_net_13934) );
na02m01 g65371_u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q), .b(g65325_sb), .o(g65371_da) );
in01m02 g65372_u0 ( .a(FE_OFN642_n_4677), .o(g65372_sb) );
na04f02 TIMEBOOST_cell_23169 ( .a(n_2918), .b(n_5230), .c(n_3367), .d(n_2846), .o(n_5232) );
in01s01 g65373_u0 ( .a(n_4669), .o(g65373_sb) );
na02f01 TIMEBOOST_cell_62991 ( .a(TIMEBOOST_net_20442), .b(g62119_db), .o(n_5577) );
na03f02 TIMEBOOST_cell_73064 ( .a(TIMEBOOST_net_22033), .b(FE_OFN709_n_8232), .c(g62015_sb), .o(n_7865) );
in01m01 g65374_u0 ( .a(FE_OFN640_n_4669), .o(g65374_sb) );
na04m04 TIMEBOOST_cell_67888 ( .a(n_3785), .b(FE_OFN1643_n_4671), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q), .d(g65345_sb), .o(TIMEBOOST_net_7590) );
na02m06 TIMEBOOST_cell_45825 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q), .o(TIMEBOOST_net_13807) );
in01m01 g65375_u0 ( .a(FE_OFN653_n_4508), .o(g65375_sb) );
na04f02 TIMEBOOST_cell_67280 ( .a(TIMEBOOST_net_20226), .b(FE_OFN916_n_4725), .c(g64336_sb), .d(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q), .o(TIMEBOOST_net_15064) );
na02m01 g65375_u2 ( .a(n_4452), .b(FE_OFN653_n_4508), .o(g65375_db) );
in01m01 g65376_u0 ( .a(FE_OFN1059_n_4727), .o(g65376_sb) );
na02f02 TIMEBOOST_cell_37598 ( .a(g58081_sb), .b(FE_OFN223_n_9844), .o(TIMEBOOST_net_10411) );
in01s02 TIMEBOOST_cell_67733 ( .a(TIMEBOOST_net_21160), .o(pci_target_unit_fifos_pcir_data_in_162) );
na02f02 TIMEBOOST_cell_37599 ( .a(TIMEBOOST_net_10411), .b(g58081_db), .o(n_9713) );
in01m01 g65377_u0 ( .a(n_4669), .o(g65377_sb) );
na02m03 TIMEBOOST_cell_39794 ( .a(g58331_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q), .o(TIMEBOOST_net_11509) );
na02m02 TIMEBOOST_cell_49594 ( .a(TIMEBOOST_net_15014), .b(g63616_sb), .o(n_7153) );
in01m01 g65378_u0 ( .a(FE_OFN652_n_4508), .o(g65378_sb) );
na02s01 TIMEBOOST_cell_53397 ( .a(pci_target_unit_fifos_pcir_data_in_160), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q), .o(TIMEBOOST_net_16916) );
na03f04 TIMEBOOST_cell_23171 ( .a(FE_OCPN1823_n_16560), .b(FE_OCP_RBN2223_n_15347), .c(n_15376), .o(n_15377) );
na02s01 TIMEBOOST_cell_31129 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(g65760_sb), .o(TIMEBOOST_net_9669) );
in01m01 g65379_u0 ( .a(FE_OFN652_n_4508), .o(g65379_sb) );
na03m02 TIMEBOOST_cell_69140 ( .a(n_4488), .b(g64765_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q), .o(TIMEBOOST_net_21778) );
na02f01 TIMEBOOST_cell_70338 ( .a(TIMEBOOST_net_17286), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_22377) );
in01m01 g65380_u0 ( .a(FE_OFN1642_n_4671), .o(g65380_sb) );
na02f01 TIMEBOOST_cell_49692 ( .a(TIMEBOOST_net_15063), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_13167) );
na02s01 TIMEBOOST_cell_45259 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q), .o(TIMEBOOST_net_13524) );
in01m01 g65381_u0 ( .a(FE_OFN1680_n_4655), .o(g65381_sb) );
in01s01 TIMEBOOST_cell_73902 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .o(TIMEBOOST_net_23467) );
na02m02 TIMEBOOST_cell_44101 ( .a(g58380_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q), .o(TIMEBOOST_net_12945) );
in01m01 g65382_u0 ( .a(FE_OFN1677_n_4655), .o(g65382_sb) );
na03m06 TIMEBOOST_cell_48473 ( .a(n_4465), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q), .c(FE_OFN636_n_4669), .o(TIMEBOOST_net_14454) );
na03f20 TIMEBOOST_cell_64322 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q), .b(n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_399), .o(TIMEBOOST_net_20391) );
in01m02 g65383_u0 ( .a(FE_OFN1678_n_4655), .o(g65383_sb) );
na03s01 TIMEBOOST_cell_64394 ( .a(TIMEBOOST_net_12275), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_396), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q), .o(TIMEBOOST_net_16794) );
in01m01 g65384_u0 ( .a(FE_OFN1680_n_4655), .o(g65384_sb) );
na03s02 TIMEBOOST_cell_67935 ( .a(TIMEBOOST_net_20398), .b(FE_OFN563_n_9895), .c(g57918_sb), .o(TIMEBOOST_net_9430) );
in01m04 g65385_u0 ( .a(FE_OFN1677_n_4655), .o(g65385_sb) );
na02s02 TIMEBOOST_cell_63089 ( .a(TIMEBOOST_net_20491), .b(g58201_sb), .o(TIMEBOOST_net_17345) );
na02s01 TIMEBOOST_cell_53975 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q), .o(TIMEBOOST_net_17205) );
in01m01 g65387_u0 ( .a(FE_OFN1677_n_4655), .o(g65387_sb) );
na03f04 TIMEBOOST_cell_70314 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_403), .b(FE_OFN2247_n_2113), .c(g54138_sb), .o(TIMEBOOST_net_22365) );
na03s01 TIMEBOOST_cell_68034 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q), .b(FE_OFN540_n_9690), .c(FE_OFN268_n_9880), .o(TIMEBOOST_net_12984) );
na02m02 TIMEBOOST_cell_44102 ( .a(TIMEBOOST_net_12945), .b(g58380_db), .o(n_9008) );
in01m02 g65388_u0 ( .a(FE_OFN639_n_4669), .o(g65388_sb) );
na04s06 TIMEBOOST_cell_72558 ( .a(TIMEBOOST_net_14179), .b(FE_OFN952_n_2055), .c(g65722_sb), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q), .o(TIMEBOOST_net_22028) );
in01m02 g65389_u0 ( .a(FE_OFN1677_n_4655), .o(g65389_sb) );
na02m04 TIMEBOOST_cell_62632 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_136), .o(TIMEBOOST_net_20263) );
in01s01 TIMEBOOST_cell_73903 ( .a(TIMEBOOST_net_23467), .o(TIMEBOOST_net_23468) );
na03f02 TIMEBOOST_cell_73760 ( .a(TIMEBOOST_net_16055), .b(FE_OFN1774_n_13800), .c(FE_OFN1771_n_14054), .o(g74872_p) );
in01s01 g65390_u0 ( .a(n_2629), .o(g65390_sb) );
na02m01 TIMEBOOST_cell_68980 ( .a(n_4280), .b(FE_OFN636_n_4669), .o(TIMEBOOST_net_21698) );
na02s01 g65390_u2 ( .a(n_16307), .b(n_2629), .o(g65390_db) );
na02f03 TIMEBOOST_cell_18458 ( .a(n_16966), .b(TIMEBOOST_net_5592), .o(TIMEBOOST_net_449) );
in01m02 g65391_u0 ( .a(FE_OFN642_n_4677), .o(g65391_sb) );
na02m08 TIMEBOOST_cell_54121 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_125), .o(TIMEBOOST_net_17278) );
na02m08 TIMEBOOST_cell_52737 ( .a(pci_target_unit_pcit_if_strd_addr_in_692), .b(n_2541), .o(TIMEBOOST_net_16586) );
in01m01 g65392_u0 ( .a(FE_OFN1680_n_4655), .o(g65392_sb) );
na04f04 TIMEBOOST_cell_36098 ( .a(parchk_pci_ad_out_in_1176), .b(g62110_sb), .c(configuration_wb_err_data_579), .d(FE_OFN1165_n_5615), .o(n_5588) );
na02f02 TIMEBOOST_cell_50570 ( .a(TIMEBOOST_net_15502), .b(g62574_sb), .o(n_6405) );
na03f02 TIMEBOOST_cell_66748 ( .a(TIMEBOOST_net_16827), .b(FE_OFN1306_n_13124), .c(g54359_sb), .o(n_13083) );
in01m01 g65393_u0 ( .a(FE_OFN640_n_4669), .o(g65393_sb) );
no03f10 TIMEBOOST_cell_72511 ( .a(n_1403), .b(FE_OCP_RBN2000_n_1403), .c(n_1397), .o(TIMEBOOST_net_17208) );
in01m04 g65394_u0 ( .a(FE_OFN1677_n_4655), .o(g65394_sb) );
na04f04 TIMEBOOST_cell_24300 ( .a(n_9064), .b(g57303_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q), .d(FE_OFN1416_n_8567), .o(n_10405) );
in01s01 TIMEBOOST_cell_73852 ( .a(n_7400), .o(TIMEBOOST_net_23417) );
in01m02 g65395_u0 ( .a(FE_OFN1678_n_4655), .o(g65395_sb) );
no02f10 TIMEBOOST_cell_68164 ( .a(n_2866), .b(FE_RN_637_0), .o(TIMEBOOST_net_21290) );
na02f02 TIMEBOOST_cell_54624 ( .a(TIMEBOOST_net_17529), .b(FE_OFN1294_n_4098), .o(TIMEBOOST_net_15481) );
in01m04 g65396_u0 ( .a(FE_OFN1680_n_4655), .o(g65396_sb) );
na04f04 TIMEBOOST_cell_36100 ( .a(parchk_pci_ad_out_in_1173), .b(g62107_sb), .c(configuration_wb_err_data_576), .d(FE_OFN1174_n_5592), .o(n_5593) );
in01m06 g65397_u0 ( .a(FE_OFN1677_n_4655), .o(g65397_sb) );
in01s01 TIMEBOOST_cell_73853 ( .a(TIMEBOOST_net_23417), .o(TIMEBOOST_net_23418) );
in01m01 g65398_u0 ( .a(FE_OFN644_n_4677), .o(g65398_sb) );
na02s02 TIMEBOOST_cell_52765 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(g65708_sb), .o(TIMEBOOST_net_16600) );
in01m01 g65399_u0 ( .a(FE_OFN1643_n_4671), .o(g65399_sb) );
na02m01 TIMEBOOST_cell_47995 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q), .b(n_3747), .o(TIMEBOOST_net_14215) );
na02m01 TIMEBOOST_cell_52739 ( .a(pci_target_unit_pcit_if_strd_addr_in_697), .b(pci_target_unit_del_sync_addr_in_215), .o(TIMEBOOST_net_16587) );
in01m01 g65400_u0 ( .a(FE_OFN639_n_4669), .o(g65400_sb) );
na03m04 TIMEBOOST_cell_72752 ( .a(n_4444), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q), .c(TIMEBOOST_net_12544), .o(TIMEBOOST_net_17068) );
na03f02 TIMEBOOST_cell_66686 ( .a(TIMEBOOST_net_17124), .b(FE_OFN1322_n_6436), .c(g62504_sb), .o(n_6572) );
in01s01 TIMEBOOST_cell_63548 ( .a(pci_target_unit_fifos_pcir_data_in_186), .o(TIMEBOOST_net_20728) );
in01m01 g65401_u0 ( .a(FE_OFN1676_n_4655), .o(g65401_sb) );
na03f02 TIMEBOOST_cell_65006 ( .a(TIMEBOOST_net_14335), .b(g64357_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q), .o(TIMEBOOST_net_17327) );
na02s01 TIMEBOOST_cell_63060 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q), .o(TIMEBOOST_net_20477) );
in01m08 g65402_u0 ( .a(FE_OFN1643_n_4671), .o(g65402_sb) );
na03f02 TIMEBOOST_cell_68029 ( .a(TIMEBOOST_net_20535), .b(FE_OFN1270_n_4095), .c(g63148_sb), .o(n_5844) );
na02s01 TIMEBOOST_cell_52741 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q), .o(TIMEBOOST_net_16588) );
na02s01 TIMEBOOST_cell_52742 ( .a(TIMEBOOST_net_16588), .b(FE_OFN955_n_1699), .o(TIMEBOOST_net_14544) );
in01m02 g65403_u0 ( .a(FE_OFN1642_n_4671), .o(g65403_sb) );
na03f02 TIMEBOOST_cell_66409 ( .a(n_4592), .b(g61965_sb), .c(g61965_db), .o(n_6946) );
na04m04 TIMEBOOST_cell_67430 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q), .b(FE_OFN704_n_8069), .c(n_1949), .d(g61755_sb), .o(n_8304) );
in01m08 g65404_u0 ( .a(FE_OFN636_n_4669), .o(g65404_sb) );
na02s01 TIMEBOOST_cell_51569 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q), .o(TIMEBOOST_net_16002) );
na03s01 TIMEBOOST_cell_23181 ( .a(g58268_db), .b(g58268_sb), .c(FE_OFN201_n_9230), .o(n_9219) );
na03s02 TIMEBOOST_cell_23180 ( .a(FE_OFN203_n_9228), .b(g58269_sb), .c(g58269_db), .o(n_9218) );
in01m01 g65405_u0 ( .a(FE_OFN636_n_4669), .o(g65405_sb) );
na02m10 TIMEBOOST_cell_53311 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q), .o(TIMEBOOST_net_16873) );
na03m02 TIMEBOOST_cell_69002 ( .a(FE_OFN612_n_4501), .b(g64959_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q), .o(TIMEBOOST_net_21709) );
in01m01 g65406_u0 ( .a(FE_OFN1643_n_4671), .o(g65406_sb) );
na02f02 TIMEBOOST_cell_70543 ( .a(TIMEBOOST_net_22479), .b(g62786_sb), .o(n_5418) );
na02m08 TIMEBOOST_cell_52787 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q), .b(TIMEBOOST_net_12682), .o(TIMEBOOST_net_16611) );
in01m02 g65407_u0 ( .a(FE_OFN642_n_4677), .o(g65407_sb) );
na03m02 TIMEBOOST_cell_69850 ( .a(TIMEBOOST_net_14685), .b(TIMEBOOST_net_10709), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q), .o(TIMEBOOST_net_22133) );
in01m01 g65408_u0 ( .a(FE_OFN651_n_4508), .o(g65408_sb) );
na03f02 TIMEBOOST_cell_35104 ( .a(TIMEBOOST_net_10025), .b(FE_OFN2155_n_16439), .c(g58829_sb), .o(n_8609) );
na02f02 TIMEBOOST_cell_70527 ( .a(TIMEBOOST_net_22471), .b(g62769_sb), .o(n_5456) );
na02m02 TIMEBOOST_cell_68915 ( .a(TIMEBOOST_net_21665), .b(g64775_db), .o(TIMEBOOST_net_17399) );
in01m02 g65409_u0 ( .a(FE_OFN1642_n_4671), .o(g65409_sb) );
na02f01 TIMEBOOST_cell_63035 ( .a(TIMEBOOST_net_20464), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_15559) );
in01s01 TIMEBOOST_cell_73904 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .o(TIMEBOOST_net_23469) );
in01m01 g65410_u0 ( .a(FE_OFN643_n_4677), .o(g65410_sb) );
na02f02 TIMEBOOST_cell_62496 ( .a(g58093_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q), .o(TIMEBOOST_net_20195) );
na02f02 TIMEBOOST_cell_68413 ( .a(TIMEBOOST_net_21414), .b(n_2119), .o(TIMEBOOST_net_16638) );
na03m02 TIMEBOOST_cell_68834 ( .a(FE_OFN664_n_4495), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q), .c(n_4444), .o(TIMEBOOST_net_21625) );
na03m02 TIMEBOOST_cell_72574 ( .a(TIMEBOOST_net_14175), .b(g65715_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q), .o(TIMEBOOST_net_22319) );
in01m04 g65412_u0 ( .a(FE_OFN639_n_4669), .o(g65412_sb) );
na02s01 TIMEBOOST_cell_43749 ( .a(FE_OFN213_n_9124), .b(g58111_sb), .o(TIMEBOOST_net_12769) );
na03f08 TIMEBOOST_cell_32481 ( .a(TIMEBOOST_net_211), .b(FE_OCP_RBN2004_FE_OFN1026_n_16760), .c(n_16162), .o(TIMEBOOST_net_7587) );
in01m02 g65413_u0 ( .a(FE_OFN1640_n_4671), .o(g65413_sb) );
na04s02 TIMEBOOST_cell_67438 ( .a(wbs_dat_i_11_), .b(TIMEBOOST_net_575), .c(g63611_sb), .d(g63611_db), .o(n_7193) );
in01m01 g65414_u0 ( .a(FE_OFN651_n_4508), .o(g65414_sb) );
na03f04 TIMEBOOST_cell_32055 ( .a(n_2804), .b(n_2803), .c(FE_OFN2121_n_2687), .o(n_3260) );
na02s02 TIMEBOOST_cell_51876 ( .a(TIMEBOOST_net_16155), .b(g65750_sb), .o(n_1605) );
in01m02 g65415_u0 ( .a(FE_OFN1640_n_4671), .o(g65415_sb) );
na03f02 TIMEBOOST_cell_73527 ( .a(TIMEBOOST_net_15571), .b(TIMEBOOST_net_15653), .c(g54196_sb), .o(n_13422) );
na03s02 TIMEBOOST_cell_72513 ( .a(TIMEBOOST_net_12461), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q), .c(FE_OFN587_n_9692), .o(TIMEBOOST_net_14323) );
in01m08 g65416_u0 ( .a(FE_OFN1640_n_4671), .o(g65416_sb) );
na03s02 TIMEBOOST_cell_72660 ( .a(TIMEBOOST_net_12440), .b(FE_OFN1016_n_2053), .c(g65821_sb), .o(n_1895) );
na02f02 TIMEBOOST_cell_70671 ( .a(TIMEBOOST_net_22543), .b(g63081_sb), .o(n_5090) );
na02f02 TIMEBOOST_cell_50256 ( .a(TIMEBOOST_net_15345), .b(g62429_sb), .o(n_6741) );
in01m01 g65417_u0 ( .a(FE_OFN654_n_4508), .o(g65417_sb) );
na02f01 TIMEBOOST_cell_70996 ( .a(TIMEBOOST_net_20536), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_22706) );
na02m02 TIMEBOOST_cell_63059 ( .a(TIMEBOOST_net_20476), .b(g58097_sb), .o(TIMEBOOST_net_16671) );
na02s02 TIMEBOOST_cell_64169 ( .a(TIMEBOOST_net_21070), .b(g57946_sb), .o(TIMEBOOST_net_9396) );
in01m02 g65418_u0 ( .a(FE_OFN638_n_4669), .o(g65418_sb) );
na02m01 TIMEBOOST_cell_43745 ( .a(FE_OFN235_n_9834), .b(g57935_sb), .o(TIMEBOOST_net_12767) );
na02m01 TIMEBOOST_cell_52187 ( .a(configuration_wb_err_addr_555), .b(conf_wb_err_addr_in_964), .o(TIMEBOOST_net_16311) );
na04f04 TIMEBOOST_cell_73472 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q), .b(n_3627), .c(FE_OFN1222_n_6391), .d(g62480_sb), .o(n_6629) );
na03f02 TIMEBOOST_cell_73707 ( .a(TIMEBOOST_net_16480), .b(n_12313), .c(FE_OFN1566_n_12502), .o(n_12753) );
na02f02 g55235_u0 ( .a(FE_OCPN1827_n_14995), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q), .o(n_12116) );
na02s01 TIMEBOOST_cell_30983 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_12__Q), .b(FE_OFN209_n_9126), .o(TIMEBOOST_net_9596) );
na02s02 TIMEBOOST_cell_48722 ( .a(TIMEBOOST_net_14578), .b(TIMEBOOST_net_10527), .o(TIMEBOOST_net_9520) );
in01m02 g65421_u0 ( .a(FE_OFN653_n_4508), .o(g65421_sb) );
na02s01 TIMEBOOST_cell_54103 ( .a(FE_OFN239_n_9832), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q), .o(TIMEBOOST_net_17269) );
na02m01 TIMEBOOST_cell_68460 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q), .b(FE_OFN669_n_4505), .o(TIMEBOOST_net_21438) );
na02m02 TIMEBOOST_cell_54452 ( .a(TIMEBOOST_net_17443), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_15383) );
in01m06 g65422_u0 ( .a(FE_OFN653_n_4508), .o(g65422_sb) );
na02m08 TIMEBOOST_cell_52879 ( .a(wbs_dat_i_16_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q), .o(TIMEBOOST_net_16657) );
no04f08 TIMEBOOST_cell_23194 ( .a(n_7216), .b(wishbone_slave_unit_wbs_sm_wbr_control_in_190), .c(n_16456), .d(n_16455), .o(g75081_p) );
in01m01 g65423_u0 ( .a(FE_OFN644_n_4677), .o(g65423_sb) );
na02f01 TIMEBOOST_cell_49700 ( .a(TIMEBOOST_net_15067), .b(FE_OFN1129_g64577_p), .o(TIMEBOOST_net_13178) );
na03m02 TIMEBOOST_cell_72670 ( .a(TIMEBOOST_net_14265), .b(FE_OFN955_n_1699), .c(g65736_sb), .o(n_1607) );
na03s20 TIMEBOOST_cell_72462 ( .a(n_8884), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q), .c(wbu_addr_in_268), .o(TIMEBOOST_net_12391) );
in01m02 g65424_u0 ( .a(FE_OFN652_n_4508), .o(g65424_sb) );
na03s02 TIMEBOOST_cell_72674 ( .a(TIMEBOOST_net_12450), .b(FE_OFN956_n_1699), .c(g65783_sb), .o(n_1599) );
in01s01 TIMEBOOST_cell_45993 ( .a(TIMEBOOST_net_13953), .o(TIMEBOOST_net_13954) );
na03m02 TIMEBOOST_cell_73268 ( .a(pci_cbe_o_0_), .b(n_14389), .c(g52879_sb), .o(TIMEBOOST_net_665) );
in01s01 g65425_u0 ( .a(n_4725), .o(g65425_sb) );
na02s01 g65425_u2 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(n_4725), .o(g65425_db) );
na02s01 TIMEBOOST_cell_39796 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q), .b(g58439_sb), .o(TIMEBOOST_net_11510) );
in01m01 g65426_u0 ( .a(FE_OFN651_n_4508), .o(g65426_sb) );
na02f02 TIMEBOOST_cell_45414 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13601), .o(TIMEBOOST_net_12031) );
na02m08 TIMEBOOST_cell_52881 ( .a(wbs_dat_i_10_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q), .o(TIMEBOOST_net_16658) );
in01m01 g65427_u0 ( .a(FE_OFN651_n_4508), .o(g65427_sb) );
na03m02 TIMEBOOST_cell_70224 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(FE_OFN1034_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q), .o(TIMEBOOST_net_22320) );
na03s02 TIMEBOOST_cell_22352 ( .a(FE_OFN254_n_9825), .b(g58093_sb), .c(g58098_db), .o(n_9702) );
in01m06 g65428_u0 ( .a(FE_OFN652_n_4508), .o(g65428_sb) );
na02s02 TIMEBOOST_cell_39798 ( .a(g58438_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q), .o(TIMEBOOST_net_11511) );
na02m01 TIMEBOOST_cell_68618 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q), .o(TIMEBOOST_net_21517) );
in01m01 g65429_u0 ( .a(FE_OFN654_n_4508), .o(g65429_sb) );
na02m02 TIMEBOOST_cell_69228 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q), .b(n_3777), .o(TIMEBOOST_net_21822) );
na03f80 TIMEBOOST_cell_23201 ( .a(n_16436), .b(n_4686), .c(n_16438), .o(TIMEBOOST_net_414) );
in01m01 g65430_u0 ( .a(FE_OFN653_n_4508), .o(g65430_sb) );
na02s02 TIMEBOOST_cell_43731 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q), .b(g65828_sb), .o(TIMEBOOST_net_12760) );
na02m02 TIMEBOOST_cell_54394 ( .a(TIMEBOOST_net_17414), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_15667) );
in01m01 g65431_u0 ( .a(FE_OFN1036_n_4732), .o(g65431_sb) );
in01s01 TIMEBOOST_cell_67736 ( .a(TIMEBOOST_net_21162), .o(TIMEBOOST_net_21163) );
na02m10 TIMEBOOST_cell_45813 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q), .o(TIMEBOOST_net_13801) );
in01m01 g65432_u0 ( .a(FE_OFN1640_n_4671), .o(g65432_sb) );
na04s03 TIMEBOOST_cell_67432 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q), .b(FE_OFN704_n_8069), .c(n_1942), .d(g61754_sb), .o(n_8307) );
in01m01 g65433_u0 ( .a(FE_OFN653_n_4508), .o(g65433_sb) );
na03f02 TIMEBOOST_cell_73827 ( .a(TIMEBOOST_net_13802), .b(n_13903), .c(FE_OCP_RBN1962_FE_OFN1591_n_13741), .o(n_14291) );
na02f02 TIMEBOOST_cell_26216 ( .a(TIMEBOOST_net_7212), .b(FE_OFN1145_n_15261), .o(TIMEBOOST_net_675) );
na03f03 TIMEBOOST_cell_73646 ( .a(g58292_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q), .c(TIMEBOOST_net_15554), .o(TIMEBOOST_net_9385) );
in01m02 g65434_u0 ( .a(FE_OFN639_n_4669), .o(g65434_sb) );
na02m01 TIMEBOOST_cell_53325 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q), .b(FE_OCPN1839_n_1238), .o(TIMEBOOST_net_16880) );
in01m02 g65435_u0 ( .a(FE_OFN636_n_4669), .o(g65435_sb) );
na02s02 TIMEBOOST_cell_44440 ( .a(TIMEBOOST_net_13114), .b(TIMEBOOST_net_11196), .o(TIMEBOOST_net_9328) );
na02m02 TIMEBOOST_cell_25869 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q), .b(g65876_sb), .o(TIMEBOOST_net_7039) );
no02m04 g65436_u0 ( .a(pci_target_unit_wishbone_master_read_count_reg_2__Q), .b(n_987), .o(g65436_p) );
ao12m02 g65436_u1 ( .a(g65436_p), .b(pci_target_unit_wishbone_master_read_count_reg_2__Q), .c(n_987), .o(n_1180) );
no02m01 g65437_u0 ( .a(pci_target_unit_wishbone_master_read_count_0_), .b(n_1999), .o(g65437_p) );
ao12s01 g65437_u1 ( .a(g65437_p), .b(pci_target_unit_wishbone_master_read_count_0_), .c(n_1999), .o(n_3226) );
ao22f01 g65438_u0 ( .a(n_1281), .b(wbm_rty_i), .c(pci_target_unit_wishbone_master_rty_counter_1_), .d(n_705), .o(n_2223) );
no02f08 g65439_u0 ( .a(n_582), .b(n_588), .o(g65439_p) );
ao12f06 g65439_u1 ( .a(g65439_p), .b(n_582), .c(n_588), .o(n_1461) );
in01s03 g65440_u0 ( .a(pci_target_unit_fifos_pciw_control_in), .o(n_3806) );
no02f04 g65484_u0 ( .a(n_2747), .b(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .o(n_3795) );
na02f02 TIMEBOOST_cell_31045 ( .a(n_14671), .b(n_14839), .o(TIMEBOOST_net_9627) );
na02m02 g65486_u0 ( .a(n_1696), .b(wishbone_slave_unit_pcim_if_del_req_in), .o(g65486_p) );
in01m02 g65486_u1 ( .a(g65486_p), .o(n_1697) );
no02f10 g65487_u0 ( .a(n_978), .b(n_1554), .o(n_13820) );
na02f20 g65488_u0 ( .a(n_1679), .b(wbu_addr_in_253), .o(g65488_p) );
in01f10 g65488_u1 ( .a(g65488_p), .o(n_2013) );
na02f08 g65489_u0 ( .a(n_1331), .b(wbu_am1_in), .o(g65489_p) );
in01f06 g65489_u1 ( .a(g65489_p), .o(n_2699) );
na02f40 g65490_u0 ( .a(n_1413), .b(conf_wb_err_addr_in_945), .o(g65490_p) );
in01f40 g65490_u1 ( .a(g65490_p), .o(n_1669) );
no02f10 g65491_u0 ( .a(n_1371), .b(n_602), .o(g65491_p) );
in01f10 g65491_u1 ( .a(g65491_p), .o(n_2399) );
no02f08 g65492_u0 ( .a(n_1346), .b(n_668), .o(n_2409) );
no02f06 g65493_u0 ( .a(n_3023), .b(n_2803), .o(g65493_p) );
in01f04 g65493_u1 ( .a(g65493_p), .o(n_3163) );
na02f06 g65494_u0 ( .a(n_3386), .b(n_3022), .o(n_4084) );
na02f01 g65495_u0 ( .a(n_1418), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_), .o(g65495_p) );
in01f02 g65495_u1 ( .a(g65495_p), .o(n_1419) );
na02f40 g65497_u0 ( .a(n_1674), .b(wbm_adr_o_4_), .o(g65497_p) );
in01f20 g65497_u1 ( .a(g65497_p), .o(n_2012) );
no02f01 g65498_u0 ( .a(n_1215), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .o(g65498_p) );
in01f02 g65498_u1 ( .a(g65498_p), .o(n_1216) );
na03f02 TIMEBOOST_cell_73473 ( .a(TIMEBOOST_net_20596), .b(FE_OFN1285_n_4097), .c(g62452_sb), .o(n_6693) );
na02f02 g65505_u0 ( .a(configuration_wb_err_addr_557), .b(n_15445), .o(n_2625) );
no02m02 g65506_u0 ( .a(n_660), .b(wishbone_slave_unit_pci_initiator_if_read_count_2_), .o(n_1659) );
na02f01 g65507_u0 ( .a(n_3250), .b(pci_target_unit_wishbone_master_read_bound), .o(n_2807) );
no02s01 g65508_u0 ( .a(n_988), .b(n_3250), .o(n_2806) );
in01m01 g65509_u0 ( .a(n_1226), .o(n_1178) );
no02f08 g65510_u0 ( .a(n_1011), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(g65510_p) );
in01f04 g65510_u1 ( .a(g65510_p), .o(n_1226) );
na02f10 g65511_u0 ( .a(n_948), .b(pci_target_unit_del_sync_comp_cycle_count_2_), .o(g65511_p) );
in01f08 g65511_u1 ( .a(g65511_p), .o(n_1438) );
no02f02 g65512_u0 ( .a(n_1554), .b(pci_target_unit_pci_target_sm_cnf_progress), .o(n_14070) );
na02f08 g65513_u0 ( .a(n_1333), .b(wbu_am2_in), .o(g65513_p) );
in01f06 g65513_u1 ( .a(g65513_p), .o(n_2698) );
na02f40 g65514_u0 ( .a(n_947), .b(wishbone_slave_unit_del_sync_comp_cycle_count_2_), .o(g65514_p) );
in01f20 g65514_u1 ( .a(g65514_p), .o(n_1476) );
no02f08 g65515_u0 ( .a(n_1345), .b(n_596), .o(g65515_p) );
in01f04 g65515_u1 ( .a(g65515_p), .o(n_1976) );
na02f03 g65516_u0 ( .a(FE_OFN1695_n_3368), .b(wbu_cache_line_size_in_207), .o(n_2624) );
no02f10 g65517_u0 ( .a(n_3123), .b(parchk_pci_frame_reg_in), .o(g65517_p) );
in01f08 g65517_u1 ( .a(g65517_p), .o(n_2623) );
na02f02 g65518_u0 ( .a(n_2347), .b(n_2556), .o(g65518_p) );
in01f02 g65518_u1 ( .a(g65518_p), .o(n_3027) );
no02f04 g65519_u0 ( .a(n_3026), .b(n_3295), .o(n_4880) );
no02f10 g65520_u0 ( .a(n_3231), .b(n_16791), .o(g65520_p) );
in01f10 g65520_u1 ( .a(g65520_p), .o(n_3290) );
na02f04 g65521_u0 ( .a(configuration_cache_line_size_reg_2996), .b(FE_OFN1695_n_3368), .o(n_2622) );
no02f02 g65522_u0 ( .a(n_1011), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .o(g65522_p1) );
no02f01 g65522_u1 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(g65522_p2) );
na02f02 g65522_u2 ( .a(g65522_p1), .b(g65522_p2), .o(n_1015) );
na02f20 g65523_u0 ( .a(n_1985), .b(n_1374), .o(g65523_p) );
in01f10 g65523_u1 ( .a(g65523_p), .o(n_2419) );
na02f02 g65524_u0 ( .a(n_16791), .b(pciu_bar0_in_379), .o(n_2621) );
na02f40 g65525_u0 ( .a(n_1027), .b(pci_target_unit_wishbone_master_rty_counter_4_), .o(n_1177) );
no02f08 g65526_u0 ( .a(n_1974), .b(n_1477), .o(n_1975) );
na02f01 g65528_u0 ( .a(n_1999), .b(n_3164), .o(n_3166) );
na02f02 g65529_u0 ( .a(FE_OFN1695_n_3368), .b(wbu_cache_line_size_in_209), .o(n_2620) );
no02m01 g65530_u0 ( .a(n_3223), .b(n_1999), .o(g65530_p) );
in01f02 g65530_u1 ( .a(FE_OFN147_g65530_p), .o(n_3224) );
na02f02 g65531_u0 ( .a(FE_OFN1061_n_16720), .b(pciu_am1_in_518), .o(n_2984) );
no02f06 g65532_u0 ( .a(n_1972), .b(n_1548), .o(n_1973) );
na02f08 g65533_u0 ( .a(n_1971), .b(n_1391), .o(g65533_p) );
in01f06 g65533_u1 ( .a(g65533_p), .o(n_2461) );
no02f01 g65534_u0 ( .a(n_3295), .b(n_3504), .o(n_3505) );
in01f06 g65536_u0 ( .a(n_2218), .o(n_2219) );
na02s01 TIMEBOOST_cell_18559 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q), .b(FE_OFN2079_n_8069), .o(TIMEBOOST_net_5643) );
na02s01 TIMEBOOST_cell_45415 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q), .o(TIMEBOOST_net_13602) );
no02f20 g65539_u0 ( .a(n_2750), .b(n_1639), .o(n_2457) );
na02f02 TIMEBOOST_cell_70497 ( .a(TIMEBOOST_net_22456), .b(g63061_sb), .o(n_5128) );
na02s01 TIMEBOOST_cell_49443 ( .a(g58147_sb), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_14939) );
na02f10 g65543_u0 ( .a(n_1415), .b(n_1679), .o(g65543_p) );
in01f10 g65543_u1 ( .a(g65543_p), .o(n_2256) );
na02f10 g65549_u0 ( .a(n_1478), .b(n_2225), .o(g65549_p) );
in01f08 g65549_u1 ( .a(g65549_p), .o(n_2694) );
na02f08 g65550_u0 ( .a(n_1969), .b(n_1968), .o(g65550_p) );
in01f04 g65550_u1 ( .a(g65550_p), .o(n_1970) );
in01f02 g65551_u0 ( .a(n_2049), .o(n_2406) );
ao12f04 g65552_u0 ( .a(n_692), .b(n_527), .c(n_1624), .o(n_2049) );
no02f08 g65555_u0 ( .a(n_15762), .b(n_3023), .o(g65555_p) );
in01f06 g65555_u1 ( .a(g65555_p), .o(n_3378) );
na02f20 g65556_u0 ( .a(n_1363), .b(n_1369), .o(n_2708) );
no02f06 g65557_u0 ( .a(n_1805), .b(pci_gnt_i), .o(g65557_p) );
in01f02 g65557_u1 ( .a(g65557_p), .o(n_3810) );
na02f04 g65558_u0 ( .a(n_3222), .b(n_3221), .o(n_3798) );
no02s01 g65559_u0 ( .a(n_3123), .b(output_backup_devsel_out_reg_Q), .o(g65559_p) );
in01s01 g65559_u1 ( .a(g65559_p), .o(n_2619) );
no02f06 g65561_u0 ( .a(n_3023), .b(n_3022), .o(n_4086) );
na02m06 g65562_u0 ( .a(n_1416), .b(n_1175), .o(g65562_p) );
in01m04 g65562_u1 ( .a(g65562_p), .o(n_1176) );
na02s01 g65563_u0 ( .a(n_1337), .b(n_1038), .o(n_2051) );
na02m02 g65564_u0 ( .a(n_1338), .b(n_1093), .o(n_1967) );
na03f02 TIMEBOOST_cell_34934 ( .a(TIMEBOOST_net_9523), .b(FE_OFN1374_n_8567), .c(g57213_sb), .o(n_11544) );
no02m02 g65566_u0 ( .a(n_2468), .b(pci_target_unit_del_sync_sync_comp_req_pending), .o(n_2469) );
na02f10 g65567_u0 ( .a(n_1414), .b(n_1413), .o(g65567_p) );
in01f10 g65567_u1 ( .a(g65567_p), .o(n_2260) );
na02f10 g65568_u0 ( .a(n_1966), .b(n_1965), .o(g65568_p) );
in01f08 g65568_u1 ( .a(g65568_p), .o(n_2691) );
na02f04 g65569_u0 ( .a(n_2214), .b(n_2390), .o(g65569_p) );
in01f04 g65569_u1 ( .a(g65569_p), .o(n_4675) );
na02f02 g65570_u0 ( .a(n_15762), .b(n_1471), .o(g65570_p) );
in01f02 g65570_u1 ( .a(g65570_p), .o(n_2065) );
na02f10 g65571_u0 ( .a(n_1412), .b(n_1674), .o(g65571_p) );
in01f10 g65571_u1 ( .a(g65571_p), .o(n_2258) );
no02f80 g65572_u0 ( .a(n_1016), .b(n_861), .o(g65572_p1) );
no02f80 g65572_u1 ( .a(n_845), .b(n_872), .o(g65572_p2) );
na02f80 g65572_u2 ( .a(g65572_p1), .b(g65572_p2), .o(n_4686) );
in01s01 g65573_u1 ( .a(g65573_p), .o(n_2801) );
no02f01 g65574_u0 ( .a(n_3123), .b(n_205), .o(n_2799) );
in01f08 g65576_u0 ( .a(FE_OFN2121_n_2687), .o(n_1964) );
na02f02 TIMEBOOST_cell_39515 ( .a(TIMEBOOST_net_11369), .b(g63027_sb), .o(n_5192) );
na02f02 TIMEBOOST_cell_45416 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13602), .o(TIMEBOOST_net_12032) );
na02f02 g65579_u0 ( .a(n_2001), .b(pci_target_unit_wishbone_master_rty_counter_6_), .o(n_2002) );
na02f08 g65580_u0 ( .a(n_1985), .b(n_1986), .o(n_1987) );
no02f04 g65582_u0 ( .a(n_1819), .b(n_15210), .o(n_3115) );
na02f02 g65583_u0 ( .a(n_15407), .b(pci_target_unit_pci_target_sm_rd_progress), .o(g65583_p) );
in01f02 g65583_u1 ( .a(g65583_p), .o(n_13745) );
na04f04 TIMEBOOST_cell_24208 ( .a(n_9516), .b(g57424_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q), .d(FE_OFN1424_n_8567), .o(n_11311) );
no02s01 g65585_u0 ( .a(n_3020), .b(n_1133), .o(n_3021) );
na02f06 g65586_u0 ( .a(n_16810), .b(n_14913), .o(n_2614) );
na02f04 g65587_u0 ( .a(FE_OFN1061_n_16720), .b(pciu_am1_in_520), .o(n_2797) );
na02f10 g65588_u0 ( .a(n_3018), .b(n_3019), .o(g65588_p) );
in01f08 g65588_u1 ( .a(g65588_p), .o(n_5230) );
no02s01 g65589_u0 ( .a(n_1696), .b(wishbone_slave_unit_del_sync_sync_comp_req_pending), .o(n_1635) );
na02f10 g65590_u0 ( .a(n_2392), .b(n_3107), .o(g65590_p) );
in01f08 g65590_u1 ( .a(g65590_p), .o(n_7110) );
in01m08 g65592_u0 ( .a(n_4512), .o(n_4904) );
no02f02 g65595_u0 ( .a(n_3001), .b(n_2685), .o(g65595_p) );
in01f04 g65595_u1 ( .a(g65595_p), .o(n_4512) );
na03f04 TIMEBOOST_cell_64456 ( .a(n_2235), .b(n_2258), .c(n_2426), .o(TIMEBOOST_net_142) );
na02m01 g65597_u0 ( .a(n_1329), .b(n_1283), .o(n_2057) );
in01f04 g65598_u0 ( .a(n_1632), .o(n_1633) );
no02f03 g65599_u0 ( .a(n_1425), .b(n_878), .o(n_1632) );
in01m02 g65600_u0 ( .a(n_1630), .o(n_1631) );
no02m04 g65601_u0 ( .a(n_883), .b(n_1426), .o(n_1630) );
na04f06 TIMEBOOST_cell_64455 ( .a(n_1387), .b(n_1351), .c(n_1799), .d(n_1486), .o(n_2876) );
ao12f02 g65603_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .b(n_1126), .c(pci_target_unit_pci_target_if_same_read_reg), .o(n_1961) );
na02s02 TIMEBOOST_cell_49425 ( .a(FE_OFN268_n_9880), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q), .o(TIMEBOOST_net_14930) );
oa12s01 g65605_u0 ( .a(n_2779), .b(pci_target_unit_del_sync_addr_in_204), .c(n_2301), .o(n_2794) );
oa12s01 g65606_u0 ( .a(g74689_p), .b(n_1698), .c(FE_OFN2214_n_15366), .o(n_2793) );
na02s01 TIMEBOOST_cell_37587 ( .a(TIMEBOOST_net_10405), .b(g58023_db), .o(n_9767) );
na02m10 TIMEBOOST_cell_69860 ( .a(FE_OFN1057_n_4727), .b(TIMEBOOST_net_14562), .o(TIMEBOOST_net_22138) );
oa12s01 g65609_u0 ( .a(n_2612), .b(pci_target_unit_del_sync_addr_in_212), .c(n_2301), .o(n_2613) );
na02s01 TIMEBOOST_cell_37600 ( .a(g58046_sb), .b(FE_OFN219_n_9853), .o(TIMEBOOST_net_10412) );
oa12s01 g65611_u0 ( .a(n_2610), .b(pci_target_unit_del_sync_addr_in_211), .c(n_2301), .o(n_2611) );
oa12s01 g65612_u0 ( .a(n_2790), .b(pci_target_unit_del_sync_addr_in_205), .c(n_2301), .o(n_2792) );
oa12s01 g65613_u0 ( .a(n_2788), .b(pci_target_unit_del_sync_addr_in_206), .c(n_2301), .o(n_2789) );
na02f08 g65614_u0 ( .a(n_3107), .b(n_2609), .o(g65614_p) );
in01f06 g65614_u1 ( .a(g65614_p), .o(n_3089) );
oa12s01 g65615_u0 ( .a(n_2783), .b(pci_target_unit_del_sync_addr_in_209), .c(n_2301), .o(n_2787) );
oa12s01 g65616_u0 ( .a(n_2790), .b(n_2742), .c(n_2301), .o(n_4214) );
na02f08 g65617_u0 ( .a(n_3108), .b(n_3107), .o(g65617_p) );
in01f06 g65617_u1 ( .a(g65617_p), .o(n_7108) );
na02s01 g65618_u0 ( .a(n_2361), .b(n_3217), .o(n_3220) );
na02s01 g65619_u0 ( .a(n_2356), .b(n_2610), .o(n_2786) );
na02s01 g65620_u0 ( .a(n_2366), .b(n_2612), .o(n_2785) );
na02s01 g65621_u0 ( .a(n_2363), .b(n_2783), .o(n_2784) );
na02s01 g65622_u0 ( .a(n_2362), .b(n_2604), .o(n_2782) );
na02s01 g65623_u0 ( .a(n_2364), .b(n_2732), .o(n_2781) );
no02f10 g65626_u0 ( .a(n_2345), .b(n_15805), .o(g65626_p) );
in01f08 g65626_u1 ( .a(g65626_p), .o(n_3314) );
oa12m01 g65627_u0 ( .a(n_2779), .b(n_16027), .c(n_2301), .o(n_2780) );
na02s01 g65628_u0 ( .a(n_2349), .b(n_2606), .o(n_2745) );
oa12s01 g65629_u0 ( .a(n_3217), .b(n_1724), .c(FE_OFN2093_n_2301), .o(n_3219) );
ao12s02 g65630_u0 ( .a(wbs_bte_i_0_), .b(n_1666), .c(wbs_bte_i_1_), .o(n_1667) );
oa12s01 g65631_u0 ( .a(n_2606), .b(pci_target_unit_del_sync_addr_in_210), .c(n_2301), .o(n_2608) );
na02s01 g65632_u0 ( .a(n_2767), .b(n_2788), .o(n_3216) );
ao12m08 g65633_u0 ( .a(n_1134), .b(n_1628), .c(pci_target_unit_pci_target_sm_n_3), .o(n_1629) );
oa12s01 g65634_u0 ( .a(n_2604), .b(pci_target_unit_del_sync_addr_in_208), .c(n_2301), .o(n_2605) );
no02s01 g65635_u0 ( .a(n_249), .b(pci_target_unit_del_sync_req_rty_exp_clr), .o(n_738) );
in01f02 g65636_u0 ( .a(n_2701), .o(n_2387) );
ao12m02 g65639_u0 ( .a(n_3386), .b(n_1322), .c(n_1686), .o(n_3361) );
ao12f02 g65641_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_transfer), .b(n_1436), .c(n_2043), .o(n_2726) );
ao12f08 g65642_u0 ( .a(n_2430), .b(wishbone_slave_unit_pcim_sm_be_in_558), .c(wishbone_slave_unit_pcim_sm_be_in_559), .o(n_1626) );
na02f10 g65643_u0 ( .a(n_2777), .b(n_2778), .o(n_3261) );
oa12s01 g65644_u0 ( .a(n_2601), .b(pci_target_unit_del_sync_addr_in), .c(n_2301), .o(n_2603) );
no02s01 g65646_u0 ( .a(n_1327), .b(wishbone_slave_unit_del_sync_req_rty_exp_clr), .o(n_2386) );
oa12s01 g65647_u0 ( .a(n_2601), .b(n_16390), .c(n_2301), .o(n_2602) );
oa12s01 g65648_u0 ( .a(n_2732), .b(pci_target_unit_del_sync_addr_in_207), .c(n_2301), .o(n_2734) );
ao12f02 g65649_u0 ( .a(n_15371), .b(n_1524), .c(n_1326), .o(n_2446) );
ao12s01 g65650_u0 ( .a(n_434), .b(n_802), .c(n_1624), .o(n_1625) );
ao22f01 g65651_u0 ( .a(n_15755), .b(n_1332), .c(n_16001), .d(wbu_am2_in), .o(n_3016) );
oa12m06 g65652_u0 ( .a(n_1453), .b(n_3415), .c(n_1316), .o(n_1623) );
oa12m08 g65653_u0 ( .a(n_1265), .b(n_8876), .c(n_1174), .o(n_1621) );
in01f08 g65654_u0 ( .a(n_1443), .o(n_1619) );
na02m02 TIMEBOOST_cell_64126 ( .a(g58390_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q), .o(TIMEBOOST_net_21049) );
ao22f01 g65658_u0 ( .a(n_2560), .b(n_14908), .c(n_15065), .d(n_1330), .o(n_2972) );
in01s01 g65661_u0 ( .a(n_2730), .o(n_2776) );
ao22s01 g65662_u0 ( .a(n_2671), .b(n_2599), .c(n_2597), .d(parchk_pci_ad_reg_in), .o(n_2730) );
in01s01 g65664_u0 ( .a(n_2600), .o(n_2973) );
ao22s01 g65665_u0 ( .a(n_2599), .b(n_2598), .c(n_2597), .d(parchk_pci_ad_reg_in_1205), .o(n_2600) );
na02f02 TIMEBOOST_cell_48451 ( .a(TIMEBOOST_net_12405), .b(FE_OFN1011_n_4734), .o(TIMEBOOST_net_14443) );
na04f04 TIMEBOOST_cell_24819 ( .a(n_10154), .b(n_10151), .c(n_9307), .d(n_9306), .o(n_12158) );
in01m02 g65668_u0 ( .a(FE_OFN672_n_4505), .o(g65668_sb) );
na02f02 TIMEBOOST_cell_71339 ( .a(TIMEBOOST_net_22877), .b(FE_OCPN1845_n_16427), .o(TIMEBOOST_net_20618) );
na02s01 TIMEBOOST_cell_45261 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q), .o(TIMEBOOST_net_13525) );
in01m01 g65669_u0 ( .a(FE_OFN1626_n_4438), .o(g65669_sb) );
na03m02 TIMEBOOST_cell_72809 ( .a(n_4488), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q), .c(TIMEBOOST_net_12690), .o(TIMEBOOST_net_20952) );
in01m04 g65670_u0 ( .a(FE_OFN648_n_4497), .o(g65670_sb) );
na03f02 TIMEBOOST_cell_73428 ( .a(TIMEBOOST_net_21028), .b(FE_OFN1212_n_4151), .c(g62445_sb), .o(n_6705) );
na02s01 TIMEBOOST_cell_63022 ( .a(FE_OFN223_n_9844), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q), .o(TIMEBOOST_net_20458) );
na02f04 TIMEBOOST_cell_38759 ( .a(TIMEBOOST_net_10991), .b(FE_OFN1142_n_15261), .o(TIMEBOOST_net_5664) );
in01m01 g65671_u0 ( .a(FE_OFN665_n_4495), .o(g65671_sb) );
na02s01 TIMEBOOST_cell_30973 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_9__Q), .b(n_9825), .o(TIMEBOOST_net_9591) );
na02m01 g65671_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q), .b(FE_OFN665_n_4495), .o(g65671_db) );
na03f02 TIMEBOOST_cell_70758 ( .a(n_2259), .b(FE_OFN1697_n_5751), .c(wbm_adr_o_8_), .o(TIMEBOOST_net_22587) );
in01m01 g65672_u0 ( .a(FE_OFN687_n_4417), .o(g65672_sb) );
na02f04 TIMEBOOST_cell_31027 ( .a(wbu_addr_in_267), .b(n_4210), .o(TIMEBOOST_net_9618) );
na03m02 TIMEBOOST_cell_73429 ( .a(TIMEBOOST_net_17560), .b(FE_OFN1219_n_6886), .c(g62541_sb), .o(n_6485) );
na03f02 TIMEBOOST_cell_66680 ( .a(TIMEBOOST_net_16774), .b(FE_OFN1313_n_6624), .c(g62498_sb), .o(n_6587) );
in01m01 g65673_u0 ( .a(FE_OFN623_n_4409), .o(g65673_sb) );
na02s02 TIMEBOOST_cell_70735 ( .a(TIMEBOOST_net_22575), .b(FE_OFN245_n_9114), .o(TIMEBOOST_net_15214) );
in01f01 g65674_u0 ( .a(FE_OFN938_n_2292), .o(g65674_sb) );
na02f02 TIMEBOOST_cell_44342 ( .a(TIMEBOOST_net_13065), .b(FE_OFN1126_g64577_p), .o(TIMEBOOST_net_11353) );
in01m01 g65675_u0 ( .a(FE_OFN1003_n_2047), .o(g65675_sb) );
na02f02 TIMEBOOST_cell_70125 ( .a(TIMEBOOST_net_22270), .b(FE_OFN1147_n_13249), .o(TIMEBOOST_net_15115) );
na04s02 TIMEBOOST_cell_33452 ( .a(g58018_sb), .b(FE_OFN264_n_9849), .c(g58018_db), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q), .o(TIMEBOOST_net_9397) );
in01s01 g65676_u0 ( .a(FE_OFN952_n_2055), .o(g65676_sb) );
na02f02 TIMEBOOST_cell_31029 ( .a(wbu_addr_in_275), .b(n_4708), .o(TIMEBOOST_net_9619) );
in01s01 TIMEBOOST_cell_63601 ( .a(TIMEBOOST_net_20781), .o(TIMEBOOST_net_20780) );
na02s01 TIMEBOOST_cell_70462 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q), .o(TIMEBOOST_net_22439) );
in01s02 g65677_u0 ( .a(FE_OFN936_n_2292), .o(g65677_sb) );
na02s02 TIMEBOOST_cell_63322 ( .a(FE_OFN260_n_9860), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q), .o(TIMEBOOST_net_20608) );
in01s01 g65678_u0 ( .a(FE_OFN936_n_2292), .o(g65678_sb) );
na02m02 TIMEBOOST_cell_68807 ( .a(TIMEBOOST_net_21611), .b(g64333_sb), .o(n_3844) );
in01s01 TIMEBOOST_cell_73956 ( .a(wbm_dat_i_28_), .o(TIMEBOOST_net_23521) );
na02m04 TIMEBOOST_cell_72070 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q), .b(FE_OFN956_n_1699), .o(TIMEBOOST_net_23243) );
in01s01 g65679_u0 ( .a(FE_OFN1003_n_2047), .o(g65679_sb) );
na02m02 TIMEBOOST_cell_43867 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q), .b(FE_OFN956_n_1699), .o(TIMEBOOST_net_12828) );
na02m02 TIMEBOOST_cell_69159 ( .a(TIMEBOOST_net_21787), .b(g65952_db), .o(n_1845) );
in01m01 g65680_u0 ( .a(FE_OFN1074_n_4740), .o(g65680_sb) );
in01m01 g65681_u0 ( .a(FE_OFN1046_n_16657), .o(g65681_sb) );
in01s01 TIMEBOOST_cell_35485 ( .a(TIMEBOOST_net_10076), .o(TIMEBOOST_net_10075) );
na02m01 g65681_u2 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q), .b(FE_OFN1046_n_16657), .o(g65681_db) );
na02m01 TIMEBOOST_cell_43036 ( .a(TIMEBOOST_net_12412), .b(FE_OFN908_n_4734), .o(TIMEBOOST_net_10599) );
in01s01 g65682_u0 ( .a(FE_OFN953_n_2055), .o(g65682_sb) );
na03s01 TIMEBOOST_cell_41893 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q), .b(g58346_sb), .c(g58346_db), .o(n_9017) );
na02f40 TIMEBOOST_cell_62395 ( .a(TIMEBOOST_net_20144), .b(n_562), .o(n_1477) );
na03m10 TIMEBOOST_cell_73129 ( .a(TIMEBOOST_net_22138), .b(g64259_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q), .o(TIMEBOOST_net_23312) );
in01m02 g65683_u0 ( .a(FE_OFN2108_n_2047), .o(g65683_sb) );
na03f10 TIMEBOOST_cell_23856 ( .a(g75178_da), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_), .c(n_16273), .o(n_16550) );
na03f02 TIMEBOOST_cell_34946 ( .a(TIMEBOOST_net_9475), .b(FE_OFN1409_n_8567), .c(g57473_sb), .o(n_11261) );
na03s02 TIMEBOOST_cell_32785 ( .a(n_2163), .b(g61997_sb), .c(g61997_db), .o(n_7901) );
in01s01 g65684_u0 ( .a(FE_OFN941_n_2047), .o(g65684_sb) );
na02s01 TIMEBOOST_cell_45547 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q), .o(TIMEBOOST_net_13668) );
na04f40 TIMEBOOST_cell_64426 ( .a(g58771_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q), .c(FE_OFN2055_n_8831), .d(wbu_addr_in_262), .o(n_9858) );
in01m01 g65685_u0 ( .a(FE_OFN938_n_2292), .o(g65685_sb) );
na03m02 TIMEBOOST_cell_64412 ( .a(TIMEBOOST_net_17202), .b(FE_OFN936_n_2292), .c(g65677_sb), .o(n_2212) );
in01s01 g65686_u0 ( .a(FE_OFN936_n_2292), .o(g65686_sb) );
na02m02 TIMEBOOST_cell_44394 ( .a(TIMEBOOST_net_13091), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_11426) );
na02f01 TIMEBOOST_cell_68326 ( .a(n_4501), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q), .o(TIMEBOOST_net_21371) );
in01m01 g65687_u0 ( .a(FE_OFN936_n_2292), .o(g65687_sb) );
na02m01 TIMEBOOST_cell_42867 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_127), .o(TIMEBOOST_net_12328) );
na03f02 TIMEBOOST_cell_67052 ( .a(FE_OCPN2218_n_13997), .b(TIMEBOOST_net_16544), .c(FE_OFN1600_n_13995), .o(n_14493) );
na02m02 TIMEBOOST_cell_71847 ( .a(TIMEBOOST_net_23131), .b(n_3761), .o(TIMEBOOST_net_17400) );
in01s01 g65688_u0 ( .a(FE_OFN936_n_2292), .o(g65688_sb) );
na02s02 TIMEBOOST_cell_30703 ( .a(n_9582), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q), .o(TIMEBOOST_net_9456) );
in01m01 g65689_u0 ( .a(FE_OFN937_n_2292), .o(g65689_sb) );
na02f04 TIMEBOOST_cell_63814 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_413), .b(FE_OFN2249_n_1790), .o(TIMEBOOST_net_20893) );
na02s01 TIMEBOOST_cell_62949 ( .a(TIMEBOOST_net_20421), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_11195) );
in01m04 g65690_u0 ( .a(FE_OFN2108_n_2047), .o(g65690_sb) );
na03f02 TIMEBOOST_cell_34948 ( .a(TIMEBOOST_net_9502), .b(FE_OFN1421_n_8567), .c(g57150_sb), .o(n_11600) );
na02m01 TIMEBOOST_cell_39181 ( .a(TIMEBOOST_net_11202), .b(g58078_db), .o(n_9716) );
in01f01 g65691_u0 ( .a(FE_OFN1003_n_2047), .o(g65691_sb) );
na03f02 TIMEBOOST_cell_34807 ( .a(TIMEBOOST_net_9380), .b(FE_OFN1400_n_8567), .c(g57533_sb), .o(n_10312) );
na02s01 g65691_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q), .b(FE_OFN1003_n_2047), .o(g65691_db) );
na03f02 TIMEBOOST_cell_65345 ( .a(TIMEBOOST_net_16311), .b(n_5633), .c(g62124_sb), .o(n_5572) );
in01m01 g65692_u0 ( .a(FE_OFN938_n_2292), .o(g65692_sb) );
na02s01 TIMEBOOST_cell_42991 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q), .o(TIMEBOOST_net_12390) );
na02m06 TIMEBOOST_cell_45339 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q), .o(TIMEBOOST_net_13564) );
in01s01 g65693_u0 ( .a(FE_OFN2108_n_2047), .o(g65693_sb) );
na03f02 TIMEBOOST_cell_34950 ( .a(TIMEBOOST_net_9498), .b(FE_OFN1414_n_8567), .c(g57295_sb), .o(n_11457) );
na04f02 TIMEBOOST_cell_36832 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q), .b(FE_OFN1394_n_8567), .c(n_9073), .d(g57270_sb), .o(n_10417) );
in01s01 g65694_u0 ( .a(FE_OFN950_n_2055), .o(g65694_sb) );
na03m02 TIMEBOOST_cell_64420 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q), .b(g65960_sb), .c(g65960_db), .o(n_2162) );
na03m02 TIMEBOOST_cell_48133 ( .a(n_3761), .b(FE_OFN1625_n_4438), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q), .o(TIMEBOOST_net_14284) );
in01s01 g65695_u0 ( .a(FE_OFN938_n_2292), .o(g65695_sb) );
na04m02 TIMEBOOST_cell_67916 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q), .b(FE_OFN1076_n_4740), .c(g64136_sb), .d(pci_target_unit_fifos_pciw_addr_data_in_127), .o(n_4026) );
na02s01 TIMEBOOST_cell_62948 ( .a(FE_OFN1651_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q), .o(TIMEBOOST_net_20421) );
na04f80 TIMEBOOST_cell_31924 ( .a(n_247), .b(n_104), .c(n_1416), .d(n_1715), .o(n_2218) );
in01s01 g65696_u0 ( .a(FE_OFN951_n_2055), .o(g65696_sb) );
na03f02 TIMEBOOST_cell_73647 ( .a(TIMEBOOST_net_17423), .b(FE_OFN1253_n_4143), .c(g62889_sb), .o(n_6099) );
na03s01 TIMEBOOST_cell_41857 ( .a(g58354_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q), .c(g58354_da), .o(TIMEBOOST_net_9347) );
in01s01 g65697_u0 ( .a(FE_OFN936_n_2292), .o(g65697_sb) );
na03m08 TIMEBOOST_cell_65100 ( .a(n_3777), .b(FE_OFN646_n_4497), .c(n_3672), .o(TIMEBOOST_net_14559) );
na02s01 g65697_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q), .b(FE_OFN936_n_2292), .o(g65697_db) );
in01s01 g65698_u0 ( .a(FE_OFN937_n_2292), .o(g65698_sb) );
in01s01 TIMEBOOST_cell_73905 ( .a(TIMEBOOST_net_23469), .o(TIMEBOOST_net_23470) );
na03s02 TIMEBOOST_cell_73184 ( .a(TIMEBOOST_net_10048), .b(g62069_sb), .c(TIMEBOOST_net_5643), .o(n_7830) );
in01s01 g65699_u0 ( .a(FE_OFN935_n_2292), .o(g65699_sb) );
na04f80 TIMEBOOST_cell_31927 ( .a(FE_OCP_RBN2290_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .b(n_16175), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_), .o(n_15824) );
in01s01 g65700_u0 ( .a(FE_OFN935_n_2292), .o(g65700_sb) );
na03m02 TIMEBOOST_cell_72811 ( .a(TIMEBOOST_net_21578), .b(g65005_sb), .c(TIMEBOOST_net_21855), .o(TIMEBOOST_net_17532) );
na02s01 TIMEBOOST_cell_49270 ( .a(TIMEBOOST_net_14852), .b(TIMEBOOST_net_10827), .o(TIMEBOOST_net_9381) );
in01s01 g65701_u0 ( .a(FE_OFN937_n_2292), .o(g65701_sb) );
na03f02 TIMEBOOST_cell_47306 ( .a(FE_OFN1553_n_12104), .b(TIMEBOOST_net_13591), .c(FE_OCPN1827_n_14995), .o(n_12511) );
na02s01 g65701_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN937_n_2292), .o(g65701_db) );
in01s01 TIMEBOOST_cell_67764 ( .a(TIMEBOOST_net_21190), .o(TIMEBOOST_net_21191) );
in01s01 g65702_u0 ( .a(FE_OFN2108_n_2047), .o(g65702_sb) );
na03f02 TIMEBOOST_cell_66415 ( .a(TIMEBOOST_net_17521), .b(FE_OFN1246_n_4093), .c(g62577_sb), .o(n_6400) );
in01s01 TIMEBOOST_cell_45938 ( .a(TIMEBOOST_net_13899), .o(TIMEBOOST_net_13898) );
in01s02 g65703_u0 ( .a(FE_OFN937_n_2292), .o(g65703_sb) );
na02s01 TIMEBOOST_cell_48836 ( .a(TIMEBOOST_net_14635), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_12761) );
na03f02 TIMEBOOST_cell_47308 ( .a(FE_OFN1554_n_12104), .b(TIMEBOOST_net_13593), .c(FE_OCP_RBN1979_n_10273), .o(n_12483) );
in01s02 g65704_u0 ( .a(FE_OFN955_n_1699), .o(g65704_sb) );
na04f04 TIMEBOOST_cell_73474 ( .a(n_3789), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q), .c(FE_OFN1207_n_6356), .d(g62374_sb), .o(n_6855) );
na03f02 TIMEBOOST_cell_34912 ( .a(TIMEBOOST_net_9532), .b(FE_OFN1411_n_8567), .c(g57139_sb), .o(n_11610) );
in01s01 g65705_u0 ( .a(FE_OFN951_n_2055), .o(g65705_sb) );
na02s01 g65705_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q), .b(FE_OFN951_n_2055), .o(g65705_db) );
in01s01 g65706_u0 ( .a(FE_OFN937_n_2292), .o(g65706_sb) );
na04m02 TIMEBOOST_cell_72493 ( .a(n_3764), .b(n_4671), .c(g65325_da), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q), .o(TIMEBOOST_net_17445) );
na03f02 TIMEBOOST_cell_64941 ( .a(g64367_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q), .c(TIMEBOOST_net_12478), .o(TIMEBOOST_net_13064) );
in01f01 g65707_u0 ( .a(FE_OFN938_n_2292), .o(g65707_sb) );
na03f02 TIMEBOOST_cell_73740 ( .a(TIMEBOOST_net_13587), .b(FE_OFN1741_n_11019), .c(FE_OFN1735_n_16317), .o(n_12750) );
na02m02 TIMEBOOST_cell_50055 ( .a(wbm_adr_o_18_), .b(g58799_sb), .o(TIMEBOOST_net_15245) );
in01s02 g65708_u0 ( .a(FE_OFN952_n_2055), .o(g65708_sb) );
na02m02 TIMEBOOST_cell_44398 ( .a(TIMEBOOST_net_13093), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_11430) );
na03m02 TIMEBOOST_cell_73269 ( .a(pci_cbe_o_3_), .b(n_14389), .c(g52881_sb), .o(TIMEBOOST_net_664) );
na02s01 TIMEBOOST_cell_68507 ( .a(TIMEBOOST_net_21461), .b(TIMEBOOST_net_12380), .o(TIMEBOOST_net_17297) );
in01m02 g65709_u0 ( .a(FE_OFN2109_n_2047), .o(g65709_sb) );
na02s02 TIMEBOOST_cell_48878 ( .a(TIMEBOOST_net_14656), .b(g58220_sb), .o(TIMEBOOST_net_10860) );
in01m02 g65710_u0 ( .a(FE_OFN1003_n_2047), .o(g65710_sb) );
na03m02 TIMEBOOST_cell_73270 ( .a(pci_cbe_o_2_), .b(n_14389), .c(g52880_sb), .o(TIMEBOOST_net_666) );
na02s02 TIMEBOOST_cell_53889 ( .a(g58224_sb), .b(FE_OFN245_n_9114), .o(TIMEBOOST_net_17162) );
in01m01 g65711_u0 ( .a(FE_OFN938_n_2292), .o(g65711_sb) );
na04f04 TIMEBOOST_cell_65126 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q), .b(FE_OFN1654_n_9502), .c(g58334_sb), .d(FE_OFN272_n_9828), .o(n_9483) );
na03f10 TIMEBOOST_cell_67937 ( .a(n_16485), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q), .c(n_13221), .o(g59331_p) );
na03f02 TIMEBOOST_cell_66700 ( .a(TIMEBOOST_net_17106), .b(FE_OFN1313_n_6624), .c(g62885_sb), .o(n_6107) );
in01m01 g65712_u0 ( .a(FE_OFN936_n_2292), .o(g65712_sb) );
na04f04 TIMEBOOST_cell_73430 ( .a(n_4307), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q), .c(FE_OFN1241_n_4092), .d(g62711_sb), .o(n_6148) );
na02m10 TIMEBOOST_cell_52991 ( .a(wishbone_slave_unit_pcim_sm_data_in_641), .b(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q), .o(TIMEBOOST_net_16713) );
in01s01 g65713_u0 ( .a(FE_OFN1786_n_1699), .o(g65713_sb) );
na03f02 TIMEBOOST_cell_42208 ( .a(conf_wb_err_addr_in_962), .b(g62122_sb), .c(TIMEBOOST_net_8823), .o(n_5574) );
na02s01 g65713_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q), .b(FE_OFN1786_n_1699), .o(g65713_db) );
in01s01 g65714_u0 ( .a(FE_OFN941_n_2047), .o(g65714_sb) );
na02m01 g52485_u1 ( .a(wbs_adr_i_9_), .b(g52470_sb), .o(g52485_da) );
na02m01 g65714_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q), .b(FE_OFN941_n_2047), .o(g65714_db) );
na03f02 TIMEBOOST_cell_35063 ( .a(TIMEBOOST_net_9601), .b(FE_OFN1436_n_9372), .c(g58455_sb), .o(n_9402) );
in01m01 g65715_u0 ( .a(FE_OFN1003_n_2047), .o(g65715_sb) );
na03m04 TIMEBOOST_cell_72637 ( .a(n_4473), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q), .c(TIMEBOOST_net_9755), .o(TIMEBOOST_net_17496) );
na03f02 TIMEBOOST_cell_66615 ( .a(TIMEBOOST_net_17084), .b(FE_OFN2063_n_6391), .c(g62367_sb), .o(n_6868) );
na02m02 TIMEBOOST_cell_43379 ( .a(g58313_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q), .o(TIMEBOOST_net_12584) );
na03m02 TIMEBOOST_cell_73130 ( .a(pci_target_unit_fifos_pciw_addr_data_in_131), .b(g64206_sb), .c(g64206_db), .o(n_3963) );
na02s01 g65716_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q), .b(FE_OFN1003_n_2047), .o(g65716_db) );
na03f02 TIMEBOOST_cell_73528 ( .a(TIMEBOOST_net_13287), .b(g52444_sb), .c(TIMEBOOST_net_22794), .o(n_14848) );
in01s01 g65717_u0 ( .a(FE_OFN1784_n_1699), .o(g65717_sb) );
na02s01 g65717_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q), .b(FE_OFN1784_n_1699), .o(g65717_db) );
na03f02 TIMEBOOST_cell_73761 ( .a(FE_OFN1774_n_13800), .b(TIMEBOOST_net_13706), .c(FE_OFN1768_n_14054), .o(n_14498) );
in01s01 g65718_u0 ( .a(FE_OFN935_n_2292), .o(g65718_sb) );
na02s02 TIMEBOOST_cell_53890 ( .a(TIMEBOOST_net_17162), .b(g58224_db), .o(n_9049) );
na02m08 TIMEBOOST_cell_45417 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q), .o(TIMEBOOST_net_13603) );
na04s02 TIMEBOOST_cell_67847 ( .a(TIMEBOOST_net_10339), .b(g65787_sb), .c(g61748_sb), .d(g61748_db), .o(n_8321) );
in01s01 g65719_u0 ( .a(FE_OFN936_n_2292), .o(g65719_sb) );
na02m04 TIMEBOOST_cell_72138 ( .a(n_4450), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q), .o(TIMEBOOST_net_23277) );
in01s01 g65720_u0 ( .a(FE_OFN2109_n_2047), .o(g65720_sb) );
na02f02 TIMEBOOST_cell_68961 ( .a(TIMEBOOST_net_21688), .b(TIMEBOOST_net_14429), .o(TIMEBOOST_net_17105) );
na03f02 TIMEBOOST_cell_66753 ( .a(TIMEBOOST_net_17516), .b(FE_OFN1234_n_6391), .c(g62473_sb), .o(n_6644) );
in01s02 g65721_u0 ( .a(FE_OFN953_n_2055), .o(g65721_sb) );
na02m02 TIMEBOOST_cell_52155 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q), .b(g65913_sb), .o(TIMEBOOST_net_16295) );
na04s02 TIMEBOOST_cell_72876 ( .a(TIMEBOOST_net_14149), .b(g61804_sb), .c(g65795_db), .d(g61804_db), .o(n_8186) );
na02f02 TIMEBOOST_cell_63383 ( .a(TIMEBOOST_net_20638), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_15364) );
in01m01 g65722_u0 ( .a(FE_OFN952_n_2055), .o(g65722_sb) );
na02s02 TIMEBOOST_cell_54736 ( .a(TIMEBOOST_net_17585), .b(TIMEBOOST_net_12987), .o(TIMEBOOST_net_9461) );
na02m02 TIMEBOOST_cell_62836 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q), .b(FE_OFN2257_n_8060), .o(TIMEBOOST_net_20365) );
na02m04 TIMEBOOST_cell_44971 ( .a(n_1959), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q), .o(TIMEBOOST_net_13380) );
in01s02 g65723_u0 ( .a(FE_OFN950_n_2055), .o(g65723_sb) );
in01s01 TIMEBOOST_cell_67735 ( .a(pci_target_unit_fifos_pcir_data_in_172), .o(TIMEBOOST_net_21162) );
na02f02 TIMEBOOST_cell_51174 ( .a(TIMEBOOST_net_15804), .b(g61871_sb), .o(n_8092) );
na03f02 TIMEBOOST_cell_35106 ( .a(TIMEBOOST_net_10027), .b(FE_OFN2155_n_16439), .c(g58826_sb), .o(n_8615) );
in01s02 g65724_u0 ( .a(FE_OFN956_n_1699), .o(g65724_sb) );
na02s01 g65724_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q), .b(FE_OFN956_n_1699), .o(g65724_db) );
na02m02 TIMEBOOST_cell_44951 ( .a(n_3676), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q), .o(TIMEBOOST_net_13370) );
in01s01 g65725_u0 ( .a(FE_OFN950_n_2055), .o(g65725_sb) );
na03f01 TIMEBOOST_cell_68106 ( .a(TIMEBOOST_net_14003), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q), .o(TIMEBOOST_net_21261) );
na02s01 TIMEBOOST_cell_62835 ( .a(TIMEBOOST_net_20364), .b(TIMEBOOST_net_11025), .o(TIMEBOOST_net_10023) );
na03f08 TIMEBOOST_cell_69918 ( .a(TIMEBOOST_net_16937), .b(FE_OFN1063_n_15808), .c(configuration_wb_err_cs_bit8), .o(TIMEBOOST_net_22167) );
in01s01 g65726_u0 ( .a(FE_OFN953_n_2055), .o(g65726_sb) );
na02m02 TIMEBOOST_cell_69230 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q), .b(FE_OFN1677_n_4655), .o(TIMEBOOST_net_21823) );
na03f02 TIMEBOOST_cell_73475 ( .a(TIMEBOOST_net_20950), .b(FE_OFN1284_n_4097), .c(g62372_sb), .o(n_6859) );
in01s01 g65727_u0 ( .a(FE_OFN955_n_1699), .o(g65727_sb) );
na02m10 TIMEBOOST_cell_51679 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q), .o(TIMEBOOST_net_16057) );
na03f02 TIMEBOOST_cell_34914 ( .a(TIMEBOOST_net_9518), .b(FE_OFN1413_n_8567), .c(g57170_sb), .o(n_10453) );
na02s01 TIMEBOOST_cell_48522 ( .a(TIMEBOOST_net_14478), .b(g65910_db), .o(n_1854) );
in01m02 g65728_u0 ( .a(FE_OFN953_n_2055), .o(g65728_sb) );
na02f01 TIMEBOOST_cell_62514 ( .a(n_8884), .b(wbu_addr_in_250), .o(TIMEBOOST_net_20204) );
na03f02 TIMEBOOST_cell_34880 ( .a(TIMEBOOST_net_9432), .b(FE_OFN1409_n_8567), .c(g57589_sb), .o(n_11162) );
no02m01 g65729_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .b(n_905), .o(g65729_p) );
ao12m01 g65729_u1 ( .a(g65729_p), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .c(n_905), .o(n_1609) );
in01m01 g65730_u0 ( .a(FE_OFN951_n_2055), .o(g65730_sb) );
na02f01 TIMEBOOST_cell_70262 ( .a(TIMEBOOST_net_9310), .b(FE_OFN1095_g64577_p), .o(TIMEBOOST_net_22339) );
in01s01 g65731_u0 ( .a(FE_OFN953_n_2055), .o(g65731_sb) );
in01s01 TIMEBOOST_cell_73906 ( .a(n_13611), .o(TIMEBOOST_net_23471) );
na02f02 TIMEBOOST_cell_71577 ( .a(TIMEBOOST_net_22996), .b(n_12362), .o(n_12783) );
in01s02 g65732_u0 ( .a(FE_OFN2109_n_2047), .o(g65732_sb) );
na02m02 TIMEBOOST_cell_42973 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_144), .o(TIMEBOOST_net_12381) );
in01s01 g65733_u0 ( .a(FE_OFN935_n_2292), .o(g65733_sb) );
na02s01 g65733_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q), .b(FE_OFN935_n_2292), .o(g65733_db) );
in01s01 g65734_u0 ( .a(FE_OFN1003_n_2047), .o(g65734_sb) );
na02s01 g65734_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q), .b(FE_OFN1003_n_2047), .o(g65734_db) );
in01s01 TIMEBOOST_cell_73957 ( .a(TIMEBOOST_net_23521), .o(TIMEBOOST_net_23522) );
in01s02 g65735_u0 ( .a(FE_OFN956_n_1699), .o(g65735_sb) );
na02f02 TIMEBOOST_cell_70499 ( .a(TIMEBOOST_net_22457), .b(g63135_sb), .o(n_4980) );
in01s02 g65736_u0 ( .a(FE_OFN955_n_1699), .o(g65736_sb) );
na02s02 TIMEBOOST_cell_63066 ( .a(FE_OFN250_n_9789), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q), .o(TIMEBOOST_net_20480) );
in01m01 g65737_u0 ( .a(FE_OFN941_n_2047), .o(g65737_sb) );
na02m01 TIMEBOOST_cell_42981 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_139), .o(TIMEBOOST_net_12385) );
na02m02 g65737_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q), .b(FE_OFN941_n_2047), .o(g65737_db) );
no02m08 TIMEBOOST_cell_45477 ( .a(FE_RN_722_0), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374), .o(TIMEBOOST_net_13633) );
in01m01 g65738_u0 ( .a(FE_OFN953_n_2055), .o(g65738_sb) );
na03f02 TIMEBOOST_cell_34881 ( .a(TIMEBOOST_net_9333), .b(FE_OFN1409_n_8567), .c(g57380_sb), .o(n_11367) );
na03f02 TIMEBOOST_cell_34936 ( .a(TIMEBOOST_net_9473), .b(FE_OFN1399_n_8567), .c(g57365_sb), .o(n_11382) );
in01f01 g65739_u0 ( .a(FE_OFN952_n_2055), .o(g65739_sb) );
na03f02 TIMEBOOST_cell_34937 ( .a(TIMEBOOST_net_9525), .b(FE_OFN1413_n_8567), .c(g57502_sb), .o(n_10327) );
in01s01 TIMEBOOST_cell_63573 ( .a(TIMEBOOST_net_20752), .o(TIMEBOOST_net_20753) );
in01m01 g65740_u0 ( .a(FE_OFN951_n_2055), .o(g65740_sb) );
na03f02 TIMEBOOST_cell_66470 ( .a(TIMEBOOST_net_17441), .b(FE_OFN1285_n_4097), .c(g62459_sb), .o(n_6678) );
na03f02 TIMEBOOST_cell_73476 ( .a(TIMEBOOST_net_16750), .b(FE_OFN1192_n_6935), .c(g63197_sb), .o(n_5770) );
in01s01 g65741_u0 ( .a(FE_OFN953_n_2055), .o(g65741_sb) );
na02m02 TIMEBOOST_cell_69545 ( .a(TIMEBOOST_net_21980), .b(TIMEBOOST_net_14418), .o(TIMEBOOST_net_16787) );
na02s01 g65741_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q), .b(FE_OFN953_n_2055), .o(g65741_db) );
in01s01 TIMEBOOST_cell_63572 ( .a(wishbone_slave_unit_wishbone_slave_map), .o(TIMEBOOST_net_20752) );
in01m01 g65742_u0 ( .a(FE_OFN952_n_2055), .o(g65742_sb) );
na03f02 TIMEBOOST_cell_73788 ( .a(TIMEBOOST_net_13744), .b(FE_OFN1600_n_13995), .c(FE_OCPN2218_n_13997), .o(n_14467) );
na03f10 TIMEBOOST_cell_41336 ( .a(TIMEBOOST_net_10177), .b(n_1629), .c(n_8801), .o(n_9177) );
in01s01 g65743_u0 ( .a(FE_OFN951_n_2055), .o(g65743_sb) );
na03f02 TIMEBOOST_cell_34938 ( .a(TIMEBOOST_net_9526), .b(FE_OFN1368_n_8567), .c(g57298_sb), .o(n_10408) );
na02s01 TIMEBOOST_cell_48814 ( .a(TIMEBOOST_net_14624), .b(FE_OFN596_n_9694), .o(TIMEBOOST_net_12763) );
in01s02 g65744_u0 ( .a(FE_OFN951_n_2055), .o(g65744_sb) );
na02m02 TIMEBOOST_cell_37427 ( .a(TIMEBOOST_net_10325), .b(g63537_sb), .o(n_4618) );
na03f02 TIMEBOOST_cell_66417 ( .a(TIMEBOOST_net_17502), .b(FE_OFN1234_n_6391), .c(g62625_sb), .o(n_6305) );
na03f02 TIMEBOOST_cell_34939 ( .a(TIMEBOOST_net_9533), .b(FE_OFN1388_n_8567), .c(g57462_sb), .o(n_11271) );
in01s01 g65745_u0 ( .a(FE_OFN937_n_2292), .o(g65745_sb) );
na02m10 TIMEBOOST_cell_53031 ( .a(configuration_pci_err_data_528), .b(wbm_dat_o_27_), .o(TIMEBOOST_net_16733) );
in01s01 g65746_u0 ( .a(FE_OFN950_n_2055), .o(g65746_sb) );
na03m02 TIMEBOOST_cell_73015 ( .a(TIMEBOOST_net_21838), .b(FE_OFN1809_n_4454), .c(TIMEBOOST_net_22118), .o(TIMEBOOST_net_17163) );
na02s01 TIMEBOOST_cell_43363 ( .a(FE_OFN225_n_9122), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q), .o(TIMEBOOST_net_12576) );
na04f02 TIMEBOOST_cell_35110 ( .a(wbs_dat_o_9_), .b(g52534_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_108), .d(FE_OFN1471_g52675_p), .o(n_13685) );
in01s02 g65747_u0 ( .a(FE_OFN2109_n_2047), .o(g65747_sb) );
na02s02 TIMEBOOST_cell_48820 ( .a(TIMEBOOST_net_14627), .b(FE_OFN2253_n_9687), .o(TIMEBOOST_net_12764) );
na03s01 TIMEBOOST_cell_72393 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_82), .b(FE_OFN2116_wishbone_slave_unit_pci_initiator_if_data_source), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q), .o(TIMEBOOST_net_20798) );
na04f06 TIMEBOOST_cell_73271 ( .a(g65884_db), .b(TIMEBOOST_net_14831), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q), .d(FE_OFN1812_n_7845), .o(TIMEBOOST_net_15097) );
in01s01 g65748_u0 ( .a(FE_OFN955_n_1699), .o(g65748_sb) );
na03m02 TIMEBOOST_cell_72998 ( .a(TIMEBOOST_net_23219), .b(g65009_sb), .c(TIMEBOOST_net_22091), .o(TIMEBOOST_net_17095) );
na03f02 TIMEBOOST_cell_34916 ( .a(TIMEBOOST_net_9452), .b(FE_OFN1374_n_8567), .c(g57263_sb), .o(n_11490) );
in01s01 g65749_u0 ( .a(FE_OFN951_n_2055), .o(g65749_sb) );
na04f02 TIMEBOOST_cell_35111 ( .a(wbs_dat_o_8_), .b(g52533_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_107), .d(FE_OFN1471_g52675_p), .o(n_13686) );
na02s01 g65749_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q), .b(FE_OFN951_n_2055), .o(g65749_db) );
na03f20 TIMEBOOST_cell_32047 ( .a(FE_RN_527_0), .b(FE_RN_528_0), .c(FE_RN_529_0), .o(FE_OFN1060_n_16720) );
in01s01 g65750_u0 ( .a(FE_OFN1786_n_1699), .o(g65750_sb) );
in01s03 TIMEBOOST_cell_45975 ( .a(pci_target_unit_fifos_pcir_data_in_187), .o(TIMEBOOST_net_13936) );
in01m01 g65751_u0 ( .a(FE_OFN2108_n_2047), .o(g65751_sb) );
in01s01 TIMEBOOST_cell_73958 ( .a(wbm_dat_i_29_), .o(TIMEBOOST_net_23523) );
na02m02 TIMEBOOST_cell_68811 ( .a(TIMEBOOST_net_21613), .b(g65082_sb), .o(TIMEBOOST_net_20288) );
in01m01 g65752_u0 ( .a(FE_OFN1012_n_4734), .o(g65752_sb) );
na02s01 TIMEBOOST_cell_53977 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q), .o(TIMEBOOST_net_17206) );
na03f02 TIMEBOOST_cell_47310 ( .a(FE_OFN1552_n_12104), .b(TIMEBOOST_net_13595), .c(FE_OCPN1827_n_14995), .o(n_12710) );
na02m01 TIMEBOOST_cell_43795 ( .a(pci_target_unit_fifos_pciw_addr_data_in_129), .b(FE_OFN928_n_4730), .o(TIMEBOOST_net_12792) );
in01s01 g65753_u0 ( .a(FE_OFN1003_n_2047), .o(g65753_sb) );
na02f02 TIMEBOOST_cell_71490 ( .a(g59231_db), .b(g52399_db), .o(TIMEBOOST_net_22953) );
na02s01 g65753_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q), .b(FE_OFN1003_n_2047), .o(g65753_db) );
na03f10 TIMEBOOST_cell_72434 ( .a(n_2228), .b(n_2229), .c(n_2260), .o(TIMEBOOST_net_10220) );
in01s01 g65754_u0 ( .a(FE_OFN950_n_2055), .o(g65754_sb) );
na02s01 g65754_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q), .b(FE_OFN950_n_2055), .o(g65754_db) );
in01s01 g65755_u0 ( .a(FE_OFN1785_n_1699), .o(g65755_sb) );
na02f02 TIMEBOOST_cell_71323 ( .a(TIMEBOOST_net_22869), .b(g59799_sb), .o(n_7714) );
na04f02 TIMEBOOST_cell_67526 ( .a(n_4061), .b(g62738_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q), .d(FE_OFN1097_g64577_p), .o(n_5503) );
in01s01 g65756_u0 ( .a(FE_OFN1783_n_1699), .o(g65756_sb) );
na02m02 TIMEBOOST_cell_68917 ( .a(TIMEBOOST_net_21666), .b(TIMEBOOST_net_12422), .o(TIMEBOOST_net_17383) );
na02m01 g65756_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q), .b(FE_OFN1783_n_1699), .o(g65756_db) );
na02m03 TIMEBOOST_cell_52883 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_140), .o(TIMEBOOST_net_16659) );
na03f02 TIMEBOOST_cell_73708 ( .a(TIMEBOOST_net_13532), .b(n_12313), .c(FE_OFN1566_n_12502), .o(n_17035) );
in01m01 g65758_u0 ( .a(FE_OFN952_n_2055), .o(g65758_sb) );
na02m02 TIMEBOOST_cell_54517 ( .a(TIMEBOOST_net_13227), .b(FE_OFN1193_n_6935), .o(TIMEBOOST_net_17476) );
in01s01 g65759_u0 ( .a(FE_OFN951_n_2055), .o(g65759_sb) );
na03f02 TIMEBOOST_cell_66570 ( .a(TIMEBOOST_net_17131), .b(FE_OFN1313_n_6624), .c(g62401_sb), .o(n_6797) );
na04f04 TIMEBOOST_cell_46530 ( .a(n_2205), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q), .c(FE_OFN713_n_8140), .d(g61723_sb), .o(n_8376) );
na04f02 TIMEBOOST_cell_35112 ( .a(wbs_dat_o_7_), .b(g52532_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_106), .d(FE_OFN1471_g52675_p), .o(n_13687) );
in01s01 g65760_u0 ( .a(FE_OFN1783_n_1699), .o(g65760_sb) );
na02s03 TIMEBOOST_cell_62982 ( .a(configuration_wb_err_cs_bit_565), .b(TIMEBOOST_net_13843), .o(TIMEBOOST_net_20438) );
na02s01 g65760_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q), .b(FE_OFN1783_n_1699), .o(g65760_db) );
na03m02 TIMEBOOST_cell_72505 ( .a(TIMEBOOST_net_21359), .b(g64953_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q), .o(TIMEBOOST_net_21622) );
in01f02 g65761_u0 ( .a(FE_OFN1003_n_2047), .o(g65761_sb) );
na02m02 TIMEBOOST_cell_68780 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q), .b(FE_OFN681_n_4460), .o(TIMEBOOST_net_21598) );
na02m10 TIMEBOOST_cell_45275 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q), .o(TIMEBOOST_net_13532) );
na02m01 TIMEBOOST_cell_69500 ( .a(n_4452), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q), .o(TIMEBOOST_net_21958) );
in01s01 g65762_u0 ( .a(FE_OFN950_n_2055), .o(g65762_sb) );
na03f02 TIMEBOOST_cell_73477 ( .a(TIMEBOOST_net_17456), .b(FE_OFN1215_n_4151), .c(g63153_sb), .o(n_5836) );
na03f02 TIMEBOOST_cell_66928 ( .a(FE_OFN1751_n_12086), .b(TIMEBOOST_net_13621), .c(FE_OFN1572_n_11027), .o(TIMEBOOST_net_16875) );
na04m01 TIMEBOOST_cell_67128 ( .a(TIMEBOOST_net_6765), .b(g54209_sb), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_412), .d(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q), .o(TIMEBOOST_net_16800) );
in01s04 TIMEBOOST_cell_67099 ( .a(TIMEBOOST_net_21133), .o(TIMEBOOST_net_21132) );
na02s01 g65763_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q), .b(FE_OFN1003_n_2047), .o(g65763_db) );
na02s01 g65763_u1 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(g65715_sb), .o(g65763_da) );
in01m01 g65764_u0 ( .a(FE_OFN941_n_2047), .o(g65764_sb) );
na03m02 TIMEBOOST_cell_72633 ( .a(g65041_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q), .c(TIMEBOOST_net_10638), .o(TIMEBOOST_net_17572) );
na02m02 g65764_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q), .b(FE_OFN941_n_2047), .o(g65764_db) );
na02f02 TIMEBOOST_cell_49892 ( .a(TIMEBOOST_net_15163), .b(g62741_sb), .o(n_5497) );
na03m02 TIMEBOOST_cell_72634 ( .a(g65010_sb), .b(n_3636), .c(TIMEBOOST_net_12426), .o(TIMEBOOST_net_20537) );
na02s01 g65765_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q), .b(FE_OFN1003_n_2047), .o(g65765_db) );
in01s01 g65766_u0 ( .a(FE_OFN955_n_1699), .o(g65766_sb) );
na02f04 TIMEBOOST_cell_30035 ( .a(TIMEBOOST_net_5471), .b(n_14839), .o(TIMEBOOST_net_9122) );
na03f02 TIMEBOOST_cell_34918 ( .a(TIMEBOOST_net_9514), .b(FE_OFN1383_n_8567), .c(g57498_sb), .o(n_11240) );
na02f02 TIMEBOOST_cell_70911 ( .a(TIMEBOOST_net_22663), .b(g60650_sb), .o(n_5675) );
in01s01 g65767_u0 ( .a(FE_OFN953_n_2055), .o(g65767_sb) );
na02m02 TIMEBOOST_cell_37423 ( .a(TIMEBOOST_net_10323), .b(g64172_sb), .o(n_3993) );
na03f02 TIMEBOOST_cell_34680 ( .a(TIMEBOOST_net_8552), .b(g60681_db), .c(TIMEBOOST_net_7661), .o(n_14822) );
na04f02 TIMEBOOST_cell_35113 ( .a(wbs_dat_o_6_), .b(g52531_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_105), .d(FE_OFN1471_g52675_p), .o(n_13792) );
in01s02 g65768_u0 ( .a(FE_OFN956_n_1699), .o(g65768_sb) );
na02f02 TIMEBOOST_cell_71749 ( .a(TIMEBOOST_net_23082), .b(FE_OCP_RBN1961_FE_OFN1591_n_13741), .o(n_16257) );
na02s03 TIMEBOOST_cell_69171 ( .a(TIMEBOOST_net_21793), .b(TIMEBOOST_net_20166), .o(n_7975) );
in01s01 g65769_u0 ( .a(FE_OFN941_n_2047), .o(g65769_sb) );
na02m02 TIMEBOOST_cell_44613 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q), .b(g58280_sb), .o(TIMEBOOST_net_13201) );
na02s01 TIMEBOOST_cell_45419 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q), .o(TIMEBOOST_net_13604) );
in01s01 g65770_u0 ( .a(FE_OFN941_n_2047), .o(g65770_sb) );
na02s01 g65770_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q), .b(FE_OFN941_n_2047), .o(g65770_db) );
na02m02 TIMEBOOST_cell_69458 ( .a(g65281_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q), .o(TIMEBOOST_net_21937) );
in01s02 g65771_u0 ( .a(FE_OFN956_n_1699), .o(g65771_sb) );
na02f02 TIMEBOOST_cell_71147 ( .a(TIMEBOOST_net_22781), .b(g62690_sb), .o(n_7364) );
in01s01 TIMEBOOST_cell_73854 ( .a(n_7400), .o(TIMEBOOST_net_23419) );
in01m02 g65772_u0 ( .a(FE_OFN935_n_2292), .o(g65772_sb) );
na02f02 TIMEBOOST_cell_54466 ( .a(TIMEBOOST_net_17450), .b(FE_OFN1276_n_4096), .o(TIMEBOOST_net_15471) );
na02f04 g55325_u0 ( .a(FE_OFN1551_n_12104), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q), .o(n_12369) );
na03s02 TIMEBOOST_cell_41911 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q), .b(g58305_sb), .c(g58305_db), .o(n_9506) );
in01m04 g65773_u0 ( .a(FE_OFN2108_n_2047), .o(g65773_sb) );
na02m10 TIMEBOOST_cell_45341 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q), .o(TIMEBOOST_net_13565) );
no02s01 TIMEBOOST_cell_45479 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358), .b(FE_RN_725_0), .o(TIMEBOOST_net_13634) );
in01s01 g65774_u0 ( .a(FE_OFN935_n_2292), .o(g65774_sb) );
in01s01 TIMEBOOST_cell_63592 ( .a(TIMEBOOST_net_20772), .o(TIMEBOOST_net_20739) );
na03s01 TIMEBOOST_cell_72790 ( .a(TIMEBOOST_net_20219), .b(g65902_db), .c(g65902_da), .o(n_7919) );
in01s01 g65775_u0 ( .a(FE_OFN937_n_2292), .o(g65775_sb) );
na04f04 TIMEBOOST_cell_67410 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q), .b(FE_OFN2257_n_8060), .c(n_1566), .d(g61942_sb), .o(n_7939) );
in01m02 TIMEBOOST_cell_67737 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .o(TIMEBOOST_net_21164) );
in01s01 g65776_u0 ( .a(FE_OFN936_n_2292), .o(g65776_sb) );
na03f02 TIMEBOOST_cell_35057 ( .a(TIMEBOOST_net_9615), .b(FE_OFN1441_n_9372), .c(g58470_sb), .o(n_9377) );
no04f80 TIMEBOOST_cell_31934 ( .a(FE_RN_797_0), .b(FE_RN_798_0), .c(parchk_pci_ad_out_in_1168), .d(parchk_pci_ad_out_in), .o(n_584) );
in01m01 g65777_u0 ( .a(FE_OFN1783_n_1699), .o(g65777_sb) );
na02s04 TIMEBOOST_cell_72046 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q), .b(g65836_sb), .o(TIMEBOOST_net_23231) );
na02s01 g65777_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q), .b(FE_OFN1783_n_1699), .o(g65777_db) );
in01s02 g65778_u0 ( .a(FE_OFN1784_n_1699), .o(g65778_sb) );
na02s04 TIMEBOOST_cell_63302 ( .a(FE_OFN260_n_9860), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q), .o(TIMEBOOST_net_20598) );
in01s01 g65779_u0 ( .a(FE_OFN950_n_2055), .o(g65779_sb) );
na04f02 TIMEBOOST_cell_35114 ( .a(wbs_dat_o_5_), .b(g52530_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_104), .d(FE_OFN1472_g52675_p), .o(n_13793) );
na02s02 TIMEBOOST_cell_63320 ( .a(FE_OFN264_n_9849), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q), .o(TIMEBOOST_net_20607) );
na04f02 TIMEBOOST_cell_35115 ( .a(wbs_dat_o_4_), .b(g52529_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_103), .d(FE_OFN1471_g52675_p), .o(n_13688) );
in01s01 g65780_u0 ( .a(FE_OFN935_n_2292), .o(g65780_sb) );
na02s01 TIMEBOOST_cell_49249 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q), .b(FE_OFN595_n_9694), .o(TIMEBOOST_net_14842) );
na02s01 g65780_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q), .b(FE_OFN935_n_2292), .o(g65780_db) );
na03m04 TIMEBOOST_cell_72770 ( .a(n_4479), .b(n_4273), .c(TIMEBOOST_net_12593), .o(TIMEBOOST_net_17484) );
in01s01 g65781_u0 ( .a(FE_OFN950_n_2055), .o(g65781_sb) );
na03f04 TIMEBOOST_cell_66619 ( .a(TIMEBOOST_net_16464), .b(n_16748), .c(g52624_sb), .o(n_14682) );
na02s01 g65781_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q), .b(FE_OFN950_n_2055), .o(g65781_db) );
na02s01 g65781_u1 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(g65781_sb), .o(g65781_da) );
in01s01 g65782_u0 ( .a(FE_OFN1784_n_1699), .o(g65782_sb) );
na03m02 TIMEBOOST_cell_72452 ( .a(TIMEBOOST_net_10203), .b(n_4730), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q), .o(TIMEBOOST_net_23135) );
na02s01 g65782_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q), .b(FE_OFN1784_n_1699), .o(g65782_db) );
na02s02 TIMEBOOST_cell_38493 ( .a(TIMEBOOST_net_10858), .b(g58252_sb), .o(n_9542) );
in01s02 g65783_u0 ( .a(FE_OFN956_n_1699), .o(g65783_sb) );
in01s02 TIMEBOOST_cell_67101 ( .a(TIMEBOOST_net_21135), .o(TIMEBOOST_net_21134) );
na02m02 TIMEBOOST_cell_48708 ( .a(TIMEBOOST_net_14571), .b(g65693_sb), .o(n_1952) );
na02m01 g64319_u2 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(FE_OFN1034_n_4732), .o(g64319_db) );
in01s01 g65784_u0 ( .a(FE_OFN941_n_2047), .o(g65784_sb) );
na03m04 TIMEBOOST_cell_72406 ( .a(TIMEBOOST_net_9644), .b(g56933_sb), .c(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q), .o(TIMEBOOST_net_22894) );
na02s01 TIMEBOOST_cell_62834 ( .a(wbs_adr_i_8_), .b(g52477_sb), .o(TIMEBOOST_net_20364) );
na03s01 TIMEBOOST_cell_22245 ( .a(FE_OFN254_n_9825), .b(g58041_sb), .c(g58067_db), .o(n_9725) );
in01m04 g65786_u0 ( .a(FE_OFN956_n_1699), .o(g65786_sb) );
na03f02 TIMEBOOST_cell_34922 ( .a(TIMEBOOST_net_9493), .b(FE_OFN1420_n_8567), .c(g57209_sb), .o(n_11547) );
in01s01 g65787_u0 ( .a(FE_OFN941_n_2047), .o(g65787_sb) );
na03f02 TIMEBOOST_cell_70648 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q), .b(FE_OFN1115_g64577_p), .c(n_4067), .o(TIMEBOOST_net_22532) );
na03m02 TIMEBOOST_cell_68880 ( .a(n_4493), .b(g64795_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q), .o(TIMEBOOST_net_21648) );
na02s01 TIMEBOOST_cell_44615 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q), .b(g58452_sb), .o(TIMEBOOST_net_13202) );
in01s01 g65788_u0 ( .a(FE_OFN955_n_1699), .o(g65788_sb) );
na02s02 g65788_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q), .b(FE_OFN955_n_1699), .o(g65788_db) );
na03f02 TIMEBOOST_cell_72975 ( .a(g64955_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q), .c(TIMEBOOST_net_14561), .o(TIMEBOOST_net_13379) );
in01s01 g65789_u0 ( .a(FE_OFN938_n_2292), .o(g65789_sb) );
na02m02 TIMEBOOST_cell_39824 ( .a(g58290_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q), .o(TIMEBOOST_net_11524) );
na02s02 TIMEBOOST_cell_62947 ( .a(TIMEBOOST_net_20420), .b(g58179_sb), .o(TIMEBOOST_net_17303) );
in01m01 g65790_u0 ( .a(FE_OFN1785_n_1699), .o(g65790_sb) );
na03f02 TIMEBOOST_cell_73561 ( .a(TIMEBOOST_net_17078), .b(FE_OFN1233_n_6391), .c(g62614_sb), .o(n_6329) );
na02f01 TIMEBOOST_cell_68765 ( .a(TIMEBOOST_net_21590), .b(n_2301), .o(TIMEBOOST_net_378) );
in01s01 TIMEBOOST_cell_67103 ( .a(TIMEBOOST_net_21137), .o(TIMEBOOST_net_21136) );
in01s02 g65791_u0 ( .a(FE_OFN955_n_1699), .o(g65791_sb) );
in01s01 TIMEBOOST_cell_73907 ( .a(TIMEBOOST_net_23471), .o(TIMEBOOST_net_23472) );
in01s01 TIMEBOOST_cell_73928 ( .a(wbm_dat_i_15_), .o(TIMEBOOST_net_23493) );
in01m01 g65792_u0 ( .a(FE_OFN1786_n_1699), .o(g65792_sb) );
na03f20 TIMEBOOST_cell_46065 ( .a(TIMEBOOST_net_12281), .b(n_15414), .c(n_16855), .o(n_15347) );
na02m02 TIMEBOOST_cell_54518 ( .a(TIMEBOOST_net_17476), .b(g62399_sb), .o(n_6801) );
in01s02 g65793_u0 ( .a(FE_OFN955_n_1699), .o(g65793_sb) );
na02m08 TIMEBOOST_cell_53991 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_150), .o(TIMEBOOST_net_17213) );
na03m02 TIMEBOOST_cell_72932 ( .a(FE_OFN1680_n_4655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q), .c(TIMEBOOST_net_22110), .o(TIMEBOOST_net_13375) );
in01m02 g65794_u0 ( .a(FE_OFN1786_n_1699), .o(g65794_sb) );
na02f08 TIMEBOOST_cell_47529 ( .a(wishbone_slave_unit_wishbone_slave_c_state), .b(wishbone_slave_unit_wishbone_slave_c_state_2), .o(TIMEBOOST_net_13982) );
na03s02 TIMEBOOST_cell_66303 ( .a(n_1612), .b(g61820_sb), .c(g61820_db), .o(n_8150) );
in01s01 g65795_u0 ( .a(FE_OFN1784_n_1699), .o(g65795_sb) );
na02s01 g65795_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q), .b(FE_OFN1784_n_1699), .o(g65795_db) );
na04s02 TIMEBOOST_cell_46177 ( .a(g58148_sb), .b(g58148_db), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q), .d(FE_OFN264_n_9849), .o(TIMEBOOST_net_9550) );
na03f02 TIMEBOOST_cell_34945 ( .a(TIMEBOOST_net_9474), .b(FE_OFN1400_n_8567), .c(g57593_sb), .o(n_11161) );
in01m01 g65797_u0 ( .a(FE_OFN956_n_1699), .o(g65797_sb) );
na04f04 TIMEBOOST_cell_73581 ( .a(TIMEBOOST_net_16767), .b(FE_OFN1082_n_13221), .c(FE_OFN2072_n_15978), .d(g54177_sb), .o(n_13434) );
na03f02 TIMEBOOST_cell_66874 ( .a(FE_OFN1564_n_12502), .b(TIMEBOOST_net_15986), .c(n_12313), .o(n_12643) );
in01s02 g65798_u0 ( .a(FE_OFN956_n_1699), .o(g65798_sb) );
na04m04 TIMEBOOST_cell_68006 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_28__Q), .b(FE_OFN1084_n_13221), .c(TIMEBOOST_net_13431), .d(g54192_sb), .o(n_13425) );
in01s02 g65799_u0 ( .a(FE_OFN956_n_1699), .o(g65799_sb) );
na02f01 TIMEBOOST_cell_68079 ( .a(TIMEBOOST_net_21247), .b(FE_OFN988_n_574), .o(n_1483) );
na03f02 TIMEBOOST_cell_66797 ( .a(n_3948), .b(g62818_sb), .c(TIMEBOOST_net_7524), .o(n_5339) );
na03f02 TIMEBOOST_cell_73562 ( .a(TIMEBOOST_net_17496), .b(FE_OFN1231_n_6391), .c(g62529_sb), .o(n_6516) );
in01m02 g65800_u0 ( .a(FE_OFN951_n_2055), .o(g65800_sb) );
na04f02 TIMEBOOST_cell_35117 ( .a(wbs_dat_o_2_), .b(g52525_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_101), .d(FE_OFN1472_g52675_p), .o(n_13734) );
na04f02 TIMEBOOST_cell_35116 ( .a(wbs_dat_o_3_), .b(g52528_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_102), .d(FE_OFN1472_g52675_p), .o(n_13693) );
no02f04 g65801_u0 ( .a(n_908), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(g65801_p) );
ao12f02 g65801_u1 ( .a(g65801_p), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .c(n_908), .o(n_6136) );
in01s01 g65802_u0 ( .a(FE_OFN935_n_2292), .o(g65802_sb) );
na02f02 TIMEBOOST_cell_50566 ( .a(TIMEBOOST_net_15500), .b(g63158_sb), .o(n_5822) );
na02f02 TIMEBOOST_cell_70913 ( .a(TIMEBOOST_net_22664), .b(g60611_sb), .o(n_4843) );
na02f02 TIMEBOOST_cell_39828 ( .a(g58306_db), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q), .o(TIMEBOOST_net_11526) );
in01m01 g65803_u0 ( .a(FE_OFN938_n_2292), .o(g65803_sb) );
na02s01 TIMEBOOST_cell_62946 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q), .b(FE_OFN266_n_9884), .o(TIMEBOOST_net_20420) );
in01m02 g65804_u0 ( .a(FE_OFN952_n_2055), .o(g65804_sb) );
na03m06 TIMEBOOST_cell_72933 ( .a(TIMEBOOST_net_21824), .b(g65372_sb), .c(TIMEBOOST_net_22025), .o(TIMEBOOST_net_20540) );
na02s01 TIMEBOOST_cell_44616 ( .a(TIMEBOOST_net_13202), .b(g58452_db), .o(n_9405) );
na02m10 TIMEBOOST_cell_53485 ( .a(pci_target_unit_pcit_if_strd_addr_in_706), .b(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70), .o(TIMEBOOST_net_16960) );
in01s01 g65805_u0 ( .a(FE_OFN1784_n_1699), .o(g65805_sb) );
na02f02 TIMEBOOST_cell_53652 ( .a(TIMEBOOST_net_17043), .b(g63181_sb), .o(n_5788) );
no03f02 TIMEBOOST_cell_66110 ( .a(FE_RN_361_0), .b(FE_OFN1706_n_4868), .c(FE_RN_362_0), .o(TIMEBOOST_net_776) );
na02s02 TIMEBOOST_cell_63221 ( .a(TIMEBOOST_net_20557), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_10890) );
in01s01 g65806_u0 ( .a(FE_OFN1785_n_1699), .o(g65806_sb) );
na02f01 TIMEBOOST_cell_44412 ( .a(TIMEBOOST_net_13100), .b(FE_OFN1124_g64577_p), .o(TIMEBOOST_net_11444) );
na04s04 TIMEBOOST_cell_72898 ( .a(TIMEBOOST_net_17239), .b(FE_OFN1044_n_2037), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q), .d(g65825_sb), .o(TIMEBOOST_net_22063) );
in01f02 g65807_u0 ( .a(FE_OFN2108_n_2047), .o(g65807_sb) );
na02f01 TIMEBOOST_cell_53895 ( .a(TIMEBOOST_net_13070), .b(FE_OFN1123_g64577_p), .o(TIMEBOOST_net_17165) );
na02m02 g65807_u2 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q), .b(FE_OFN2108_n_2047), .o(g65807_db) );
na02s01 TIMEBOOST_cell_52831 ( .a(pci_target_unit_fifos_pciw_addr_data_in_146), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q), .o(TIMEBOOST_net_16633) );
in01f10 g65808_u3 ( .a(g65808_p), .o(n_1588) );
in01s01 g65809_u0 ( .a(FE_OFN1017_n_2053), .o(g65809_sb) );
na02m01 g65809_u2 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(FE_OFN1017_n_2053), .o(g65809_db) );
na03m02 TIMEBOOST_cell_68312 ( .a(g65077_sb), .b(g65077_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q), .o(TIMEBOOST_net_21364) );
in01s01 g65810_u0 ( .a(n_2299), .o(g65810_sb) );
na04f04 TIMEBOOST_cell_73331 ( .a(n_4032), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q), .c(FE_OFN1119_g64577_p), .d(g62785_sb), .o(n_5421) );
na02f02 TIMEBOOST_cell_37602 ( .a(g58094_sb), .b(FE_OFN243_n_9116), .o(TIMEBOOST_net_10413) );
in01s01 g65811_u0 ( .a(FE_OFN1017_n_2053), .o(g65811_sb) );
na04f06 TIMEBOOST_cell_72986 ( .a(TIMEBOOST_net_21125), .b(FE_OFN948_n_2248), .c(g65859_sb), .d(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q), .o(TIMEBOOST_net_22360) );
in01s01 g65812_u0 ( .a(FE_OFN1017_n_2053), .o(g65812_sb) );
na02s02 TIMEBOOST_cell_68624 ( .a(FE_OFN217_n_9889), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q), .o(TIMEBOOST_net_21520) );
na02s01 g65812_u2 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(FE_OFN1017_n_2053), .o(g65812_db) );
in01m01 g65813_u0 ( .a(FE_OFN776_n_15366), .o(g65813_sb) );
na03m04 TIMEBOOST_cell_72934 ( .a(TIMEBOOST_net_21825), .b(g65273_sb), .c(TIMEBOOST_net_22017), .o(TIMEBOOST_net_20967) );
na03s02 TIMEBOOST_cell_64452 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q), .b(g65849_sb), .c(g65849_db), .o(n_1586) );
na02s01 TIMEBOOST_cell_49295 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q), .b(FE_OFN559_n_9895), .o(TIMEBOOST_net_14865) );
in01s01 g65814_u0 ( .a(FE_OFN1017_n_2053), .o(g65814_sb) );
na02f02 TIMEBOOST_cell_50558 ( .a(TIMEBOOST_net_15496), .b(g62415_sb), .o(n_6768) );
na02s01 g65814_u2 ( .a(pci_target_unit_fifos_pcir_data_in_179), .b(FE_OFN1017_n_2053), .o(g65814_db) );
in01m02 g65815_u0 ( .a(FE_OFN2113_n_2053), .o(g65815_sb) );
na03f02 TIMEBOOST_cell_72935 ( .a(pci_target_unit_del_sync_addr_in_232), .b(g65245_sb), .c(TIMEBOOST_net_7153), .o(n_2637) );
na02m02 g65815_u2 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(FE_OFN2113_n_2053), .o(g65815_db) );
na03f06 TIMEBOOST_cell_64328 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q), .b(n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_388), .o(TIMEBOOST_net_17285) );
in01s01 g65816_u0 ( .a(FE_OFN1016_n_2053), .o(g65816_sb) );
na02s01 g65816_u2 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(FE_OFN1016_n_2053), .o(g65816_db) );
na02s01 TIMEBOOST_cell_37652 ( .a(g57961_sb), .b(FE_OFN227_n_9841), .o(TIMEBOOST_net_10438) );
na02m02 g65817_u2 ( .a(TIMEBOOST_net_21197), .b(FE_OFN1017_n_2053), .o(g65817_db) );
na02f02 TIMEBOOST_cell_70505 ( .a(TIMEBOOST_net_22460), .b(g62816_sb), .o(n_5345) );
in01m01 g65818_u0 ( .a(FE_OFN1016_n_2053), .o(g65818_sb) );
na02s01 TIMEBOOST_cell_53693 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q), .b(g58358_sb), .o(TIMEBOOST_net_17064) );
na02s02 g65818_u2 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(FE_OFN1016_n_2053), .o(g65818_db) );
na02m02 TIMEBOOST_cell_44483 ( .a(n_3385), .b(n_696), .o(TIMEBOOST_net_13136) );
in01m01 g65819_u0 ( .a(FE_OFN1016_n_2053), .o(g65819_sb) );
in01s02 g65820_u0 ( .a(FE_OFN2113_n_2053), .o(g65820_sb) );
na02m02 g65820_u2 ( .a(TIMEBOOST_net_21145), .b(FE_OFN2113_n_2053), .o(g65820_db) );
na02f01 TIMEBOOST_cell_68439 ( .a(TIMEBOOST_net_21427), .b(g65710_sb), .o(n_1907) );
in01m01 g65821_u0 ( .a(FE_OFN1016_n_2053), .o(g65821_sb) );
na02m04 TIMEBOOST_cell_45237 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q), .o(TIMEBOOST_net_13513) );
na03f02 TIMEBOOST_cell_34850 ( .a(TIMEBOOST_net_9383), .b(FE_OFN1377_n_8567), .c(g57598_sb), .o(n_10285) );
in01s01 g65822_u0 ( .a(FE_OFN1016_n_2053), .o(g65822_sb) );
na03f02 TIMEBOOST_cell_34940 ( .a(TIMEBOOST_net_9534), .b(FE_OFN1390_n_8567), .c(g57333_sb), .o(n_11417) );
na02s01 g65822_u2 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(FE_OFN1016_n_2053), .o(g65822_db) );
na03f02 TIMEBOOST_cell_34941 ( .a(TIMEBOOST_net_9535), .b(FE_OFN1392_n_8567), .c(g57152_sb), .o(n_11598) );
in01m01 g65823_u0 ( .a(FE_OFN1016_n_2053), .o(g65823_sb) );
na03m02 TIMEBOOST_cell_65430 ( .a(TIMEBOOST_net_10761), .b(TIMEBOOST_net_9794), .c(FE_RN_720_0), .o(TIMEBOOST_net_17468) );
na02s01 g52457_u1 ( .a(wbs_adr_i_11_), .b(g52457_sb), .o(g52457_da) );
na02s02 TIMEBOOST_cell_43075 ( .a(FE_OFN223_n_9844), .b(g58210_sb), .o(TIMEBOOST_net_12432) );
in01s01 g65824_u0 ( .a(FE_OFN1043_n_2037), .o(g65824_sb) );
na04m04 TIMEBOOST_cell_73272 ( .a(n_1562), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q), .c(FE_OFN1812_n_7845), .d(g61936_sb), .o(n_7951) );
in01s02 g65825_u0 ( .a(FE_OFN1044_n_2037), .o(g65825_sb) );
na02m06 TIMEBOOST_cell_72216 ( .a(TIMEBOOST_net_10070), .b(configuration_wb_err_addr_546), .o(TIMEBOOST_net_23316) );
in01s01 g65826_u0 ( .a(FE_OFN1043_n_2037), .o(g65826_sb) );
na03m02 TIMEBOOST_cell_67824 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q), .b(n_3783), .c(FE_OFN659_n_4392), .o(TIMEBOOST_net_16196) );
in01s02 g65827_u0 ( .a(FE_OFN1043_n_2037), .o(g65827_sb) );
na02m02 TIMEBOOST_cell_69659 ( .a(TIMEBOOST_net_22037), .b(n_3126), .o(TIMEBOOST_net_14762) );
na02m02 TIMEBOOST_cell_68458 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q), .b(FE_OFN670_n_4505), .o(TIMEBOOST_net_21437) );
na03m02 TIMEBOOST_cell_68866 ( .a(g64980_sb), .b(n_4465), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q), .o(TIMEBOOST_net_21641) );
in01s02 g65828_u0 ( .a(FE_OFN1044_n_2037), .o(g65828_sb) );
na03m02 TIMEBOOST_cell_72936 ( .a(TIMEBOOST_net_21826), .b(g65293_sb), .c(TIMEBOOST_net_22018), .o(TIMEBOOST_net_20527) );
na02s02 g65828_u2 ( .a(TIMEBOOST_net_21163), .b(FE_OFN1044_n_2037), .o(g65828_db) );
na04f04 TIMEBOOST_cell_24303 ( .a(n_9626), .b(g57299_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q), .d(FE_OFN1417_n_8567), .o(n_11452) );
in01s01 g65829_u0 ( .a(FE_OFN1043_n_2037), .o(g65829_sb) );
na04f04 TIMEBOOST_cell_42523 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_780), .c(FE_OFN2134_n_13124), .d(g54344_sb), .o(n_13097) );
na03f02 TIMEBOOST_cell_66221 ( .a(TIMEBOOST_net_21038), .b(FE_OFN1258_n_4143), .c(g63007_sb), .o(n_5868) );
in01s01 g65830_u0 ( .a(FE_OFN1044_n_2037), .o(g65830_sb) );
na02s01 TIMEBOOST_cell_49521 ( .a(n_15569), .b(FE_OFN262_n_9851), .o(TIMEBOOST_net_14978) );
na02m02 TIMEBOOST_cell_68179 ( .a(TIMEBOOST_net_21297), .b(TIMEBOOST_net_14030), .o(TIMEBOOST_net_16805) );
na02f01 TIMEBOOST_cell_68081 ( .a(TIMEBOOST_net_21248), .b(FE_OFN988_n_574), .o(n_1634) );
in01m01 g65831_u0 ( .a(FE_OFN1043_n_2037), .o(g65831_sb) );
na02m02 TIMEBOOST_cell_62833 ( .a(TIMEBOOST_net_20363), .b(g58382_da), .o(TIMEBOOST_net_9574) );
na02m02 TIMEBOOST_cell_68446 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q), .b(FE_OFN669_n_4505), .o(TIMEBOOST_net_21431) );
in01s01 g65832_u0 ( .a(FE_OFN1044_n_2037), .o(g65832_sb) );
na02m01 TIMEBOOST_cell_62806 ( .a(pci_target_unit_fifos_pciw_control_in_156), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q), .o(TIMEBOOST_net_20350) );
na02s01 TIMEBOOST_cell_48869 ( .a(FE_OFN239_n_9832), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q), .o(TIMEBOOST_net_14652) );
na02s01 TIMEBOOST_cell_49522 ( .a(TIMEBOOST_net_14978), .b(FE_OFN1793_n_9904), .o(TIMEBOOST_net_12957) );
in01s01 g65833_u0 ( .a(FE_OFN1044_n_2037), .o(g65833_sb) );
na02f01 TIMEBOOST_cell_30177 ( .a(n_2274), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_), .o(TIMEBOOST_net_9193) );
na02m08 TIMEBOOST_cell_53993 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_132), .o(TIMEBOOST_net_17214) );
in01s01 g65834_u0 ( .a(FE_OFN1043_n_2037), .o(g65834_sb) );
na02s01 TIMEBOOST_cell_48887 ( .a(FE_OFN1650_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q), .o(TIMEBOOST_net_14661) );
in01m01 g65835_u0 ( .a(n_2299), .o(g65835_sb) );
na03m02 TIMEBOOST_cell_70114 ( .a(FE_OFN1676_n_4655), .b(n_3764), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q), .o(TIMEBOOST_net_22265) );
in01m01 g65836_u0 ( .a(FE_OFN1041_n_2037), .o(g65836_sb) );
na03f02 TIMEBOOST_cell_47420 ( .a(FE_OFN1586_n_13736), .b(TIMEBOOST_net_13732), .c(FE_OCP_RBN1999_n_13971), .o(n_14432) );
na02m02 g65836_u2 ( .a(pci_target_unit_fifos_pcir_data_in_180), .b(FE_OFN1041_n_2037), .o(g65836_db) );
na03f02 TIMEBOOST_cell_72508 ( .a(n_2247), .b(n_1293), .c(FE_OFN1117_g64577_p), .o(TIMEBOOST_net_22474) );
in01s01 g65837_u0 ( .a(FE_OFN1043_n_2037), .o(g65837_sb) );
na02m01 TIMEBOOST_cell_68625 ( .a(TIMEBOOST_net_21520), .b(FE_OFN1631_n_9531), .o(TIMEBOOST_net_20363) );
na02s01 TIMEBOOST_cell_48888 ( .a(TIMEBOOST_net_14661), .b(FE_OFN215_n_9856), .o(TIMEBOOST_net_10864) );
na02s01 TIMEBOOST_cell_63898 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q), .o(TIMEBOOST_net_20935) );
in01s02 g65838_u0 ( .a(FE_OFN1042_n_2037), .o(g65838_sb) );
na03s02 TIMEBOOST_cell_72907 ( .a(TIMEBOOST_net_12445), .b(g65908_sb), .c(FE_OFN1016_n_2053), .o(n_1855) );
na02m01 TIMEBOOST_cell_71884 ( .a(n_3744), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q), .o(TIMEBOOST_net_23150) );
in01m01 g65839_u0 ( .a(FE_OFN1041_n_2037), .o(g65839_sb) );
in01s01 TIMEBOOST_cell_73959 ( .a(TIMEBOOST_net_23523), .o(TIMEBOOST_net_23524) );
na02m02 g65839_u2 ( .a(pci_target_unit_fifos_pcir_data_in_184), .b(FE_OFN1041_n_2037), .o(g65839_db) );
no04f10 TIMEBOOST_cell_72421 ( .a(FE_RN_685_0), .b(n_2864), .c(n_436), .d(FE_RN_686_0), .o(TIMEBOOST_net_117) );
in01m01 g65840_u0 ( .a(FE_OFN1041_n_2037), .o(g65840_sb) );
na03f06 TIMEBOOST_cell_65786 ( .a(TIMEBOOST_net_20402), .b(FE_OFN1151_n_13249), .c(g54155_sb), .o(n_13444) );
na03m02 TIMEBOOST_cell_72607 ( .a(TIMEBOOST_net_21473), .b(FE_OFN636_n_4669), .c(TIMEBOOST_net_21734), .o(TIMEBOOST_net_16783) );
na03f04 TIMEBOOST_cell_65675 ( .a(TIMEBOOST_net_20386), .b(FE_OFN2128_n_16497), .c(g54304_sb), .o(n_13028) );
in01s01 g65841_u0 ( .a(FE_OFN1042_n_2037), .o(g65841_sb) );
na04f04 TIMEBOOST_cell_24306 ( .a(n_9631), .b(g57296_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q), .d(FE_OFN1419_n_8567), .o(n_11456) );
na03m04 TIMEBOOST_cell_72609 ( .a(TIMEBOOST_net_21474), .b(FE_OFN640_n_4669), .c(TIMEBOOST_net_21725), .o(TIMEBOOST_net_17510) );
na02m02 TIMEBOOST_cell_37340 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q), .b(n_3752), .o(TIMEBOOST_net_10282) );
in01s01 g65842_u0 ( .a(FE_OFN1041_n_2037), .o(g65842_sb) );
na04m01 TIMEBOOST_cell_72412 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_90), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .c(g54209_sb), .d(wishbone_slave_unit_pcim_if_wbw_addr_data_in_403), .o(n_13175) );
na03m02 TIMEBOOST_cell_72999 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q), .b(FE_OFN1049_n_16657), .c(TIMEBOOST_net_16631), .o(TIMEBOOST_net_23272) );
na03f02 TIMEBOOST_cell_73762 ( .a(TIMEBOOST_net_13699), .b(FE_OFN1774_n_13800), .c(FE_OFN1770_n_14054), .o(g53183_p) );
in01s02 g65843_u0 ( .a(FE_OFN1042_n_2037), .o(g65843_sb) );
na02s02 g65843_u2 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(FE_OFN1042_n_2037), .o(g65843_db) );
na03f02 TIMEBOOST_cell_72679 ( .a(TIMEBOOST_net_16184), .b(FE_OFN786_n_2678), .c(g65225_sb), .o(n_2662) );
in01s01 g65844_u0 ( .a(FE_OFN1042_n_2037), .o(g65844_sb) );
na04f04 TIMEBOOST_cell_24310 ( .a(n_9637), .b(g57292_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q), .d(FE_OFN1424_n_8567), .o(n_11460) );
na03s02 TIMEBOOST_cell_64449 ( .a(wbs_dat_i_9_), .b(TIMEBOOST_net_603), .c(g63616_db), .o(TIMEBOOST_net_15014) );
in01m02 g65845_u0 ( .a(FE_OFN1041_n_2037), .o(g65845_sb) );
na03f02 TIMEBOOST_cell_65676 ( .a(g58386_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q), .c(TIMEBOOST_net_11183), .o(TIMEBOOST_net_9544) );
na02m02 g65845_u2 ( .a(TIMEBOOST_net_21185), .b(FE_OFN1041_n_2037), .o(g65845_db) );
na03f02 TIMEBOOST_cell_66432 ( .a(TIMEBOOST_net_17049), .b(n_6431), .c(g62563_sb), .o(n_6433) );
in01s01 g65846_u0 ( .a(FE_OFN1044_n_2037), .o(g65846_sb) );
na03f02 TIMEBOOST_cell_73199 ( .a(TIMEBOOST_net_14835), .b(FE_OFN1092_g64577_p), .c(g63562_sb), .o(n_4112) );
in01s01 g65847_u0 ( .a(FE_OFN946_n_2248), .o(g65847_sb) );
na02f02 TIMEBOOST_cell_71045 ( .a(TIMEBOOST_net_22730), .b(g62890_sb), .o(n_6097) );
na02s01 g65847_u2 ( .a(pci_target_unit_fifos_pcir_data_in), .b(FE_OFN946_n_2248), .o(g65847_db) );
na02m02 TIMEBOOST_cell_69051 ( .a(TIMEBOOST_net_21733), .b(g65409_sb), .o(TIMEBOOST_net_10631) );
in01m02 g65848_u0 ( .a(FE_OFN948_n_2248), .o(g65848_sb) );
na03s01 TIMEBOOST_cell_72395 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_78), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .c(g54205_sb), .o(TIMEBOOST_net_20794) );
na02s02 TIMEBOOST_cell_63896 ( .a(FE_OFN209_n_9126), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q), .o(TIMEBOOST_net_20934) );
in01s01 g65849_u0 ( .a(FE_OFN945_n_2248), .o(g65849_sb) );
na02s01 TIMEBOOST_cell_29359 ( .a(parchk_pci_ad_out_in_1189), .b(configuration_wb_err_data_592), .o(TIMEBOOST_net_8784) );
na02s01 g65849_u2 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(FE_OFN945_n_2248), .o(g65849_db) );
na03f02 TIMEBOOST_cell_73273 ( .a(TIMEBOOST_net_23318), .b(FE_OFN1174_n_5592), .c(g62121_sb), .o(n_5575) );
in01s01 g65850_u0 ( .a(FE_OFN946_n_2248), .o(g65850_sb) );
na02s02 TIMEBOOST_cell_37243 ( .a(TIMEBOOST_net_10233), .b(g65745_sb), .o(n_2195) );
na03f02 TIMEBOOST_cell_73173 ( .a(n_1872), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q), .c(FE_OFN712_n_8140), .o(TIMEBOOST_net_14911) );
in01f02 g65851_u0 ( .a(FE_OFN959_n_2299), .o(g65851_sb) );
na03f02 TIMEBOOST_cell_73741 ( .a(TIMEBOOST_net_13677), .b(n_11831), .c(n_12357), .o(n_12616) );
na02f04 g65851_u2 ( .a(TIMEBOOST_net_23388), .b(FE_OFN959_n_2299), .o(g65851_db) );
na04m06 TIMEBOOST_cell_67279 ( .a(n_3739), .b(g64822_sb), .c(g64822_db), .d(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q), .o(TIMEBOOST_net_20605) );
in01s01 g65852_u0 ( .a(FE_OFN946_n_2248), .o(g65852_sb) );
na02f01 TIMEBOOST_cell_27203 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q), .b(FE_OFN1125_g64577_p), .o(TIMEBOOST_net_7706) );
in01s01 g65853_u0 ( .a(FE_OFN945_n_2248), .o(g65853_sb) );
na02s01 TIMEBOOST_cell_29361 ( .a(parchk_pci_ad_out_in_1178), .b(configuration_wb_err_data_581), .o(TIMEBOOST_net_8785) );
na02s01 g65853_u2 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(FE_OFN945_n_2248), .o(g65853_db) );
in01m01 g65854_u0 ( .a(FE_OFN2111_n_2248), .o(g65854_sb) );
na02f02 TIMEBOOST_cell_50716 ( .a(TIMEBOOST_net_15575), .b(g54203_sb), .o(TIMEBOOST_net_13389) );
na02f01 g65854_u2 ( .a(pci_target_unit_fifos_pcir_data_in_159), .b(FE_OFN2111_n_2248), .o(g65854_db) );
na02s02 TIMEBOOST_cell_48882 ( .a(TIMEBOOST_net_14658), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_10889) );
in01m01 g65855_u0 ( .a(FE_OFN1017_n_2053), .o(g65855_sb) );
in01s01 TIMEBOOST_cell_63607 ( .a(TIMEBOOST_net_20787), .o(TIMEBOOST_net_20786) );
na02m10 TIMEBOOST_cell_45235 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q), .o(TIMEBOOST_net_13512) );
in01f01 g65856_u0 ( .a(FE_OFN948_n_2248), .o(g65856_sb) );
na04f04 TIMEBOOST_cell_24788 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q), .b(g58814_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q), .d(FE_OFN2157_n_16439), .o(n_8627) );
na02m02 TIMEBOOST_cell_50444 ( .a(TIMEBOOST_net_15439), .b(g62994_sb), .o(n_5894) );
na04f04 TIMEBOOST_cell_24789 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q), .b(g58813_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q), .d(FE_OFN2153_n_16439), .o(n_8628) );
in01f01 g65857_u0 ( .a(FE_OFN945_n_2248), .o(g65857_sb) );
na02s01 TIMEBOOST_cell_29363 ( .a(parchk_pci_ad_out_in_1175), .b(configuration_wb_err_data_578), .o(TIMEBOOST_net_8786) );
na02m02 TIMEBOOST_cell_50248 ( .a(TIMEBOOST_net_15341), .b(g62899_sb), .o(n_6079) );
in01m04 g65858_u0 ( .a(FE_OFN776_n_15366), .o(g65858_sb) );
na02s01 TIMEBOOST_cell_38776 ( .a(TIMEBOOST_net_7106), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_11000) );
in01s01 TIMEBOOST_cell_73861 ( .a(TIMEBOOST_net_23425), .o(TIMEBOOST_net_23426) );
in01m02 g65859_u0 ( .a(FE_OFN948_n_2248), .o(g65859_sb) );
na02m02 TIMEBOOST_cell_68727 ( .a(TIMEBOOST_net_21571), .b(g65073_sb), .o(TIMEBOOST_net_9704) );
in01s01 g65860_u0 ( .a(FE_OFN945_n_2248), .o(g65860_sb) );
na02s01 g65860_u2 ( .a(pci_target_unit_fifos_pcir_data_in_161), .b(FE_OFN945_n_2248), .o(g65860_db) );
na03f06 TIMEBOOST_cell_66001 ( .a(g62861_sb), .b(FE_OFN2105_g64577_p), .c(TIMEBOOST_net_16972), .o(n_5244) );
in01s01 g65861_u0 ( .a(n_2299), .o(g65861_sb) );
na02m02 TIMEBOOST_cell_71869 ( .a(TIMEBOOST_net_23142), .b(g65805_sb), .o(n_1668) );
na02s01 TIMEBOOST_cell_43447 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q), .o(TIMEBOOST_net_12618) );
in01f02 g65862_u0 ( .a(FE_OFN948_n_2248), .o(g65862_sb) );
na02f02 g65862_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q), .b(g65862_sb), .o(g65862_da) );
na02f01 g65862_u2 ( .a(pci_target_unit_fifos_pcir_data_in_164), .b(FE_OFN948_n_2248), .o(g65862_db) );
na02f01 g65862_u3 ( .a(g65862_da), .b(g65862_db), .o(n_1707) );
in01m01 g65863_u0 ( .a(FE_OFN945_n_2248), .o(g65863_sb) );
na02s01 TIMEBOOST_cell_29365 ( .a(configuration_wb_err_cs_bit_567), .b(parchk_pci_cbe_out_in), .o(TIMEBOOST_net_8787) );
na02f02 TIMEBOOST_cell_39834 ( .a(n_3168), .b(FE_OFN1699_n_5751), .o(TIMEBOOST_net_11529) );
na03f02 TIMEBOOST_cell_65923 ( .a(TIMEBOOST_net_16408), .b(FE_OFN1174_n_5592), .c(g62076_sb), .o(n_5635) );
na02s02 TIMEBOOST_cell_49300 ( .a(TIMEBOOST_net_14867), .b(TIMEBOOST_net_10841), .o(TIMEBOOST_net_9411) );
na04f06 TIMEBOOST_cell_73582 ( .a(TIMEBOOST_net_15678), .b(FE_OFN1084_n_13221), .c(wishbone_slave_unit_del_sync_addr_out_reg_16__Q), .d(g54179_sb), .o(n_13432) );
in01s01 g65865_u0 ( .a(FE_OFN945_n_2248), .o(g65865_sb) );
na02s01 TIMEBOOST_cell_29367 ( .a(parchk_pci_ad_out_in_1186), .b(configuration_wb_err_data_589), .o(TIMEBOOST_net_8788) );
na02s01 g65865_u2 ( .a(pci_target_unit_fifos_pcir_data_in_169), .b(FE_OFN945_n_2248), .o(g65865_db) );
in01s01 g65866_u0 ( .a(FE_OFN946_n_2248), .o(g65866_sb) );
na02m01 g65866_u2 ( .a(pci_target_unit_fifos_pcir_data_in_168), .b(FE_OFN946_n_2248), .o(g65866_db) );
in01s01 g65867_u0 ( .a(FE_OFN945_n_2248), .o(g65867_sb) );
na02f02 TIMEBOOST_cell_53896 ( .a(TIMEBOOST_net_17165), .b(g62781_sb), .o(n_5429) );
na02s01 g65867_u2 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(FE_OFN945_n_2248), .o(g65867_db) );
na02s01 TIMEBOOST_cell_51571 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q), .o(TIMEBOOST_net_16003) );
in01s01 g65868_u0 ( .a(FE_OFN1016_n_2053), .o(g65868_sb) );
na02m02 TIMEBOOST_cell_69078 ( .a(g65054_sb), .b(n_3616), .o(TIMEBOOST_net_21747) );
na02m01 g65868_u2 ( .a(pci_target_unit_fifos_pcir_data_in_167), .b(FE_OFN1016_n_2053), .o(g65868_db) );
na02s02 TIMEBOOST_cell_64163 ( .a(TIMEBOOST_net_21067), .b(g57977_sb), .o(TIMEBOOST_net_9336) );
in01m01 g65869_u0 ( .a(FE_OFN1041_n_2037), .o(g65869_sb) );
na03m02 TIMEBOOST_cell_72611 ( .a(TIMEBOOST_net_21475), .b(FE_OFN651_n_4508), .c(TIMEBOOST_net_21715), .o(TIMEBOOST_net_17138) );
na03f02 TIMEBOOST_cell_73828 ( .a(TIMEBOOST_net_13797), .b(n_13873), .c(FE_OFN1593_n_13741), .o(n_14416) );
in01s01 g65870_u0 ( .a(n_2299), .o(g65870_sb) );
na02f01 TIMEBOOST_cell_45420 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13604), .o(TIMEBOOST_net_12034) );
na02s01 g65870_u2 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(n_2299), .o(g65870_db) );
na04f02 TIMEBOOST_cell_42553 ( .a(g52604_sb), .b(TIMEBOOST_net_11893), .c(n_3139), .d(n_10256), .o(n_11867) );
in01m02 g65871_u0 ( .a(FE_OFN644_n_4677), .o(g65871_sb) );
na03m02 TIMEBOOST_cell_73000 ( .a(TIMEBOOST_net_23181), .b(n_4482), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q), .o(TIMEBOOST_net_17122) );
na03m02 TIMEBOOST_cell_72588 ( .a(TIMEBOOST_net_21432), .b(g64755_sb), .c(TIMEBOOST_net_21635), .o(TIMEBOOST_net_20950) );
in01s01 g65872_u0 ( .a(FE_OFN1042_n_2037), .o(g65872_sb) );
na03s02 TIMEBOOST_cell_64446 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q), .b(g65849_sb), .c(g65885_db), .o(n_1657) );
na03m02 TIMEBOOST_cell_72586 ( .a(TIMEBOOST_net_21430), .b(g64761_sb), .c(TIMEBOOST_net_21623), .o(TIMEBOOST_net_20956) );
in01m01 g65873_u0 ( .a(n_4490), .o(g65873_sb) );
na03f06 TIMEBOOST_cell_73648 ( .a(FE_OFN1712_n_13563), .b(FE_OFN1946_n_13784), .c(TIMEBOOST_net_13545), .o(n_13731) );
na02m01 g65873_u2 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q), .b(n_4490), .o(g65873_db) );
in01s02 g65874_u0 ( .a(FE_OFN1042_n_2037), .o(g65874_sb) );
na02s02 g65874_u2 ( .a(pci_target_unit_fifos_pcir_data_in_166), .b(FE_OFN1042_n_2037), .o(g65874_db) );
na04f04 TIMEBOOST_cell_24315 ( .a(n_9651), .b(g57282_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q), .d(FE_OFN1405_n_8567), .o(n_11473) );
in01m01 g65875_u0 ( .a(n_2299), .o(g65875_sb) );
in01s01 TIMEBOOST_cell_73990 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .o(TIMEBOOST_net_23555) );
na02f01 g65875_u2 ( .a(pci_target_unit_fifos_pcir_data_in_158), .b(n_2299), .o(g65875_db) );
in01m02 g65876_u0 ( .a(FE_OFN1015_n_2053), .o(g65876_sb) );
na02s01 TIMEBOOST_cell_48815 ( .a(FE_OFN1666_n_9477), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q), .o(TIMEBOOST_net_14625) );
in01m01 g65877_u0 ( .a(FE_OFN1016_n_2053), .o(g65877_sb) );
na02m01 g64980_u2 ( .a(FE_OFN685_n_4417), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q), .o(g64980_db) );
na03f02 TIMEBOOST_cell_66678 ( .a(TIMEBOOST_net_17133), .b(FE_OFN1322_n_6436), .c(g62636_sb), .o(n_6278) );
na02s01 TIMEBOOST_cell_53067 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q), .b(g58283_sb), .o(TIMEBOOST_net_16751) );
in01m01 g65878_u0 ( .a(FE_OFN959_n_2299), .o(g65878_sb) );
na02m01 g65878_u2 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(FE_OFN959_n_2299), .o(g65878_db) );
na04m02 TIMEBOOST_cell_46565 ( .a(FE_OFN231_n_9839), .b(FE_OFN572_n_9502), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q), .d(g58324_sb), .o(n_9490) );
in01m01 g65879_u0 ( .a(n_4669), .o(g65879_sb) );
in01s01 TIMEBOOST_cell_45896 ( .a(TIMEBOOST_net_13857), .o(TIMEBOOST_net_13856) );
na03m02 TIMEBOOST_cell_72495 ( .a(n_3747), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q), .c(TIMEBOOST_net_21732), .o(TIMEBOOST_net_17027) );
in01m01 g65880_u0 ( .a(FE_OFN1017_n_2053), .o(g65880_sb) );
na02s01 g65880_u2 ( .a(TIMEBOOST_net_21183), .b(FE_OFN1017_n_2053), .o(g65880_db) );
in01m01 g65881_u0 ( .a(FE_OFN1016_n_2053), .o(g65881_sb) );
na03f08 TIMEBOOST_cell_64445 ( .a(wishbone_slave_unit_pcim_if_wbw_addr_data_in_390), .b(FE_OFN2059_n_13447), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q), .o(TIMEBOOST_net_20402) );
na03f04 TIMEBOOST_cell_66681 ( .a(TIMEBOOST_net_17016), .b(FE_OFN1248_n_4093), .c(g62917_sb), .o(n_6045) );
in01s02 g65882_u0 ( .a(FE_OFN2113_n_2053), .o(g65882_sb) );
na02f01 TIMEBOOST_cell_63863 ( .a(TIMEBOOST_net_20917), .b(FE_OFN1128_g64577_p), .o(TIMEBOOST_net_15162) );
na02m02 g65882_u2 ( .a(TIMEBOOST_net_21191), .b(FE_OFN2113_n_2053), .o(g65882_db) );
na03f02 TIMEBOOST_cell_65220 ( .a(FE_OFN1689_n_9528), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q), .c(g58303_sb), .o(TIMEBOOST_net_14646) );
in01m01 g65883_u0 ( .a(FE_OFN651_n_4508), .o(g65883_sb) );
na02m02 TIMEBOOST_cell_68946 ( .a(n_4476), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q), .o(TIMEBOOST_net_21681) );
in01m04 g65884_u0 ( .a(FE_OFN2113_n_2053), .o(g65884_sb) );
na02m10 TIMEBOOST_cell_45467 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q), .o(TIMEBOOST_net_13628) );
na02m06 g65884_u2 ( .a(TIMEBOOST_net_21211), .b(FE_OFN2113_n_2053), .o(g65884_db) );
na02s02 TIMEBOOST_cell_53069 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_16752) );
na02s01 TIMEBOOST_cell_29369 ( .a(parchk_pci_ad_out_in_1194), .b(configuration_wb_err_data_597), .o(TIMEBOOST_net_8789) );
na02s01 g65885_u2 ( .a(pci_target_unit_fifos_pcir_data_in_178), .b(FE_OFN945_n_2248), .o(g65885_db) );
na02m02 TIMEBOOST_cell_70337 ( .a(TIMEBOOST_net_22376), .b(g63609_sb), .o(n_7155) );
na02f02 TIMEBOOST_cell_72075 ( .a(TIMEBOOST_net_23245), .b(g60687_sb), .o(n_7218) );
in01m02 g65887_u0 ( .a(FE_OFN1041_n_2037), .o(g65887_sb) );
na03m02 TIMEBOOST_cell_72592 ( .a(TIMEBOOST_net_21434), .b(g64773_sb), .c(TIMEBOOST_net_21523), .o(TIMEBOOST_net_20544) );
na02m02 TIMEBOOST_cell_50332 ( .a(TIMEBOOST_net_15383), .b(g62932_sb), .o(n_6017) );
na02s02 TIMEBOOST_cell_54172 ( .a(TIMEBOOST_net_17303), .b(g58179_db), .o(TIMEBOOST_net_9540) );
in01m01 g65888_u0 ( .a(FE_OFN682_n_4460), .o(g65888_sb) );
na02s01 TIMEBOOST_cell_52430 ( .a(TIMEBOOST_net_16432), .b(g58454_sb), .o(TIMEBOOST_net_9476) );
in01m01 g65889_u0 ( .a(FE_OFN634_n_4454), .o(g65889_sb) );
na02m06 TIMEBOOST_cell_69720 ( .a(FE_OFN1677_n_4655), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q), .o(TIMEBOOST_net_22068) );
na02f01 TIMEBOOST_cell_44348 ( .a(TIMEBOOST_net_13068), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_11321) );
in01m01 g65890_u0 ( .a(FE_OFN1041_n_2037), .o(g65890_sb) );
na04m04 TIMEBOOST_cell_72965 ( .a(TIMEBOOST_net_13893), .b(g65768_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q), .d(TIMEBOOST_net_12828), .o(TIMEBOOST_net_22315) );
na03f02 TIMEBOOST_cell_66931 ( .a(FE_OFN1575_n_12028), .b(TIMEBOOST_net_13624), .c(FE_OFN1556_n_12042), .o(n_12499) );
in01s01 g65891_u0 ( .a(FE_OFN946_n_2248), .o(g65891_sb) );
na03f02 TIMEBOOST_cell_73274 ( .a(TIMEBOOST_net_23316), .b(FE_OFN1166_n_5615), .c(g62115_sb), .o(n_5581) );
in01s02 g65892_u0 ( .a(FE_OFN775_n_15366), .o(g65892_sb) );
na02s01 TIMEBOOST_cell_49399 ( .a(pci_target_unit_del_sync_addr_in_222), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_14917) );
na02f02 TIMEBOOST_cell_70530 ( .a(TIMEBOOST_net_13109), .b(FE_OFN1130_g64577_p), .o(TIMEBOOST_net_22473) );
in01s02 g65893_u0 ( .a(FE_OFN775_n_15366), .o(g65893_sb) );
na03s02 TIMEBOOST_cell_65796 ( .a(TIMEBOOST_net_17268), .b(g57937_sb), .c(TIMEBOOST_net_12917), .o(TIMEBOOST_net_9413) );
na02m02 TIMEBOOST_cell_47669 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q), .b(g65958_sb), .o(TIMEBOOST_net_14052) );
in01s01 g65894_u0 ( .a(FE_OFN1041_n_2037), .o(g65894_sb) );
na04m06 TIMEBOOST_cell_67425 ( .a(g58190_db), .b(FE_OFN239_n_9832), .c(g58190_sb), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q), .o(TIMEBOOST_net_16848) );
na03f02 TIMEBOOST_cell_72997 ( .a(TIMEBOOST_net_21619), .b(n_4470), .c(FE_OFN1278_n_4097), .o(TIMEBOOST_net_22772) );
na02f01 TIMEBOOST_cell_63955 ( .a(TIMEBOOST_net_20963), .b(FE_OFN1249_n_4093), .o(TIMEBOOST_net_15809) );
na02f01 TIMEBOOST_cell_18393 ( .a(n_8527), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .o(TIMEBOOST_net_5560) );
na03f08 TIMEBOOST_cell_64443 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q), .b(FE_OFN2059_n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_386), .o(TIMEBOOST_net_16983) );
na03f02 TIMEBOOST_cell_35065 ( .a(TIMEBOOST_net_9593), .b(FE_OFN1439_n_9372), .c(g58459_sb), .o(n_9396) );
in01s01 g65896_u0 ( .a(FE_OFN1015_n_2053), .o(g65896_sb) );
na02s01 TIMEBOOST_cell_68183 ( .a(TIMEBOOST_net_21299), .b(g65964_sb), .o(n_2159) );
na02m01 g65896_u2 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(FE_OFN1015_n_2053), .o(g65896_db) );
in01m01 g65897_u0 ( .a(FE_OFN1678_n_4655), .o(g65897_sb) );
na02m02 TIMEBOOST_cell_71972 ( .a(g65931_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q), .o(TIMEBOOST_net_23194) );
na03m02 TIMEBOOST_cell_69048 ( .a(FE_OFN615_n_4501), .b(g64976_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q), .o(TIMEBOOST_net_21732) );
in01s01 g65899_u0 ( .a(FE_OFN1042_n_2037), .o(g65899_sb) );
na02s02 g65899_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q), .b(g65899_sb), .o(g65899_da) );
na02s02 g65899_u2 ( .a(TIMEBOOST_net_21195), .b(FE_OFN1042_n_2037), .o(g65899_db) );
na02s02 g65899_u3 ( .a(g65899_db), .b(g65899_da), .o(n_1719) );
in01m02 g65900_u0 ( .a(FE_OFN948_n_2248), .o(g65900_sb) );
na04f04 TIMEBOOST_cell_24790 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q), .b(g58812_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q), .d(FE_OFN2153_n_16439), .o(n_8629) );
na04f04 TIMEBOOST_cell_24791 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q), .b(g58811_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q), .d(FE_OFN2158_n_16439), .o(n_8630) );
in01m01 g65901_u0 ( .a(FE_OFN1044_n_2037), .o(g65901_sb) );
na04f04 TIMEBOOST_cell_24316 ( .a(n_9653), .b(g57280_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q), .d(FE_OFN1415_n_8567), .o(n_11474) );
na02s02 TIMEBOOST_cell_71426 ( .a(FE_OFN266_n_9884), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q), .o(TIMEBOOST_net_22921) );
na03f02 TIMEBOOST_cell_73789 ( .a(TIMEBOOST_net_16528), .b(FE_OFN1602_n_13995), .c(FE_OCPN2218_n_13997), .o(g53298_p) );
in01s01 g65902_u0 ( .a(FE_OFN946_n_2248), .o(g65902_sb) );
na02s01 g65902_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q), .b(g65902_sb), .o(g65902_da) );
na02s01 g65902_u2 ( .a(pci_target_unit_fifos_pcir_data_in_165), .b(FE_OFN946_n_2248), .o(g65902_db) );
in01f01 g65903_u0 ( .a(FE_OFN959_n_2299), .o(g65903_sb) );
na02s02 TIMEBOOST_cell_44439 ( .a(g58427_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q), .o(TIMEBOOST_net_13114) );
na04s02 TIMEBOOST_cell_46563 ( .a(TIMEBOOST_net_10781), .b(g65829_sb), .c(g61894_sb), .d(g61894_db), .o(n_8039) );
in01f02 g65904_u0 ( .a(FE_OFN959_n_2299), .o(g65904_sb) );
na02f04 g65904_u2 ( .a(TIMEBOOST_net_23384), .b(FE_OFN959_n_2299), .o(g65904_db) );
na02s02 TIMEBOOST_cell_71367 ( .a(TIMEBOOST_net_22891), .b(g58049_sb), .o(TIMEBOOST_net_14936) );
in01f01 g65905_u0 ( .a(FE_OFN912_n_4727), .o(g65905_sb) );
na02f02 g65905_u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q), .b(g65905_sb), .o(g65905_da) );
na03m02 TIMEBOOST_cell_69948 ( .a(TIMEBOOST_net_12719), .b(FE_OFN1033_n_4732), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_22182) );
na02s01 TIMEBOOST_cell_47636 ( .a(TIMEBOOST_net_14035), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_385), .o(n_13168) );
in01s01 g65906_u0 ( .a(FE_OFN2113_n_2053), .o(g65906_sb) );
na02s01 g65906_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q), .b(g65906_sb), .o(g65906_da) );
no03f04 TIMEBOOST_cell_72437 ( .a(TIMEBOOST_net_101), .b(n_2430), .c(TIMEBOOST_net_12318), .o(g63943_p) );
in01s01 g65907_u0 ( .a(n_2299), .o(g65907_sb) );
na02m04 TIMEBOOST_cell_69614 ( .a(pci_target_unit_fifos_pciw_addr_data_in_137), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q), .o(TIMEBOOST_net_22015) );
na02m01 g65907_u2 ( .a(pci_target_unit_fifos_pcir_data_in_172), .b(n_2299), .o(g65907_db) );
na03f02 TIMEBOOST_cell_73141 ( .a(TIMEBOOST_net_14726), .b(g63549_sb), .c(g63549_db), .o(TIMEBOOST_net_9310) );
in01m01 g65908_u0 ( .a(FE_OFN1016_n_2053), .o(g65908_sb) );
na02m01 TIMEBOOST_cell_68313 ( .a(TIMEBOOST_net_21364), .b(n_3752), .o(TIMEBOOST_net_17113) );
na03f02 TIMEBOOST_cell_73763 ( .a(TIMEBOOST_net_13703), .b(FE_OFN1774_n_13800), .c(FE_OFN1771_n_14054), .o(g53175_p) );
in01f01 g65909_u0 ( .a(FE_OFN1797_n_2299), .o(g65909_sb) );
na03f02 TIMEBOOST_cell_66942 ( .a(FE_OFN1752_n_12086), .b(TIMEBOOST_net_16018), .c(FE_OFN2209_n_11027), .o(n_12596) );
in01s01 g65910_u0 ( .a(FE_OFN1016_n_2053), .o(g65910_sb) );
no03f10 TIMEBOOST_cell_23671 ( .a(g63430_p), .b(FE_RN_151_0), .c(FE_RN_150_0), .o(n_2939) );
na02s01 g65910_u2 ( .a(pci_target_unit_fifos_pcir_data_in_183), .b(FE_OFN1016_n_2053), .o(g65910_db) );
na03f02 TIMEBOOST_cell_73443 ( .a(TIMEBOOST_net_20965), .b(FE_OFN1250_n_4093), .c(g62530_sb), .o(n_6514) );
na03m04 TIMEBOOST_cell_72668 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(FE_OFN644_n_4677), .c(TIMEBOOST_net_23214), .o(n_1871) );
na04m06 TIMEBOOST_cell_67372 ( .a(g65407_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q), .c(n_4452), .d(FE_OFN642_n_4677), .o(n_4232) );
na02m01 TIMEBOOST_cell_71828 ( .a(FE_OFN1817_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q), .o(TIMEBOOST_net_23122) );
na02m02 TIMEBOOST_cell_52775 ( .a(FE_OFN619_n_4490), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q), .o(TIMEBOOST_net_16605) );
na02s01 g65912_u2 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(FE_OFN945_n_2248), .o(g65912_db) );
in01m01 g65913_u0 ( .a(FE_OFN1015_n_2053), .o(g65913_sb) );
na03f02 TIMEBOOST_cell_68838 ( .a(n_4488), .b(g64995_db), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q), .o(TIMEBOOST_net_21627) );
no03f02 TIMEBOOST_cell_66933 ( .a(FE_OCP_RBN2291_FE_OFN1575_n_12028), .b(FE_RN_726_0), .c(TIMEBOOST_net_13634), .o(n_12647) );
na03f02 TIMEBOOST_cell_34933 ( .a(TIMEBOOST_net_9522), .b(FE_OFN1391_n_8567), .c(g57587_sb), .o(n_10290) );
in01f01 g65914_u0 ( .a(FE_OFN948_n_2248), .o(g65914_sb) );
na02s02 TIMEBOOST_cell_25335 ( .a(wishbone_slave_unit_delayed_write_data_comp_wdata_out_84), .b(FE_OFN2118_wishbone_slave_unit_pci_initiator_if_data_source), .o(TIMEBOOST_net_6772) );
in01m01 g65915_u0 ( .a(FE_OFN1035_n_4732), .o(g65915_sb) );
na02m01 g65915_u2 ( .a(pci_target_unit_fifos_pciw_control_in_157), .b(FE_OFN1035_n_4732), .o(g65915_db) );
na02m02 TIMEBOOST_cell_69670 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q), .b(FE_OFN2257_n_8060), .o(TIMEBOOST_net_22043) );
in01m01 g65916_u0 ( .a(FE_OFN1640_n_4671), .o(g65916_sb) );
na02f02 TIMEBOOST_cell_69207 ( .a(TIMEBOOST_net_21811), .b(n_2022), .o(TIMEBOOST_net_17176) );
na02s01 TIMEBOOST_cell_53694 ( .a(TIMEBOOST_net_17064), .b(TIMEBOOST_net_11117), .o(TIMEBOOST_net_9514) );
na03f02 TIMEBOOST_cell_73583 ( .a(TIMEBOOST_net_22827), .b(FE_OFN1083_n_13221), .c(TIMEBOOST_net_22872), .o(n_13499) );
na04f04 TIMEBOOST_cell_73491 ( .a(n_3290), .b(pciu_bar0_in_376), .c(n_3040), .d(n_2826), .o(n_4652) );
na03s01 TIMEBOOST_cell_64742 ( .a(pci_target_unit_del_sync_addr_in_231), .b(g66415_sb), .c(g66415_db), .o(n_2518) );
in01m02 g65919_u0 ( .a(FE_OFN1017_n_2053), .o(g65919_sb) );
na02m04 TIMEBOOST_cell_45347 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q), .o(TIMEBOOST_net_13568) );
na02s04 g65919_u2 ( .a(TIMEBOOST_net_21201), .b(FE_OFN1015_n_2053), .o(g65919_db) );
na02f01 TIMEBOOST_cell_54676 ( .a(TIMEBOOST_net_17555), .b(FE_OFN1283_n_4097), .o(TIMEBOOST_net_15391) );
in01f01 g65920_u0 ( .a(FE_OFN948_n_2248), .o(g65920_sb) );
na04f04 TIMEBOOST_cell_24792 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q), .b(g58810_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q), .d(FE_OFN2153_n_16439), .o(n_8631) );
na02m08 TIMEBOOST_cell_69452 ( .a(g65075_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q), .o(TIMEBOOST_net_21934) );
na04f04 TIMEBOOST_cell_24793 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q), .b(g58809_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q), .d(FE_OFN2158_n_16439), .o(n_8632) );
in01m06 g65921_u0 ( .a(FE_OFN661_n_4392), .o(g65921_sb) );
na02m02 TIMEBOOST_cell_69054 ( .a(g64960_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q), .o(TIMEBOOST_net_21735) );
na02m08 g65921_u2 ( .a(FE_OFN661_n_4392), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q), .o(g65921_db) );
in01s01 TIMEBOOST_cell_73973 ( .a(TIMEBOOST_net_23537), .o(TIMEBOOST_net_23538) );
na03f02 TIMEBOOST_cell_47176 ( .a(TIMEBOOST_net_13450), .b(g53904_sb), .c(FE_OFN1327_n_13547), .o(n_13537) );
na02f04 TIMEBOOST_cell_42824 ( .a(TIMEBOOST_net_12306), .b(g58797_sb), .o(n_9868) );
na03f02 TIMEBOOST_cell_49643 ( .a(n_1748), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q), .c(FE_OFN720_n_8060), .o(TIMEBOOST_net_15039) );
in01s01 g65923_u0 ( .a(FE_OFN946_n_2248), .o(g65923_sb) );
na02f02 TIMEBOOST_cell_39679 ( .a(TIMEBOOST_net_11451), .b(g62791_sb), .o(n_5406) );
na02s02 g65923_u2 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(FE_OFN946_n_2248), .o(g65923_db) );
na02f02 TIMEBOOST_cell_54433 ( .a(n_4349), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q), .o(TIMEBOOST_net_17434) );
in01m02 g65924_u0 ( .a(FE_OFN1043_n_2037), .o(g65924_sb) );
na03f02 TIMEBOOST_cell_72571 ( .a(TIMEBOOST_net_23135), .b(g60688_sb), .c(FE_OFN1132_g64577_p), .o(TIMEBOOST_net_22482) );
na03s02 TIMEBOOST_cell_64440 ( .a(TIMEBOOST_net_12832), .b(g61969_db), .c(g63612_sb), .o(TIMEBOOST_net_16382) );
na03f02 TIMEBOOST_cell_73764 ( .a(TIMEBOOST_net_16057), .b(FE_OFN1774_n_13800), .c(FE_OFN1770_n_14054), .o(n_16226) );
in01s01 TIMEBOOST_cell_73924 ( .a(wbm_dat_i_13_), .o(TIMEBOOST_net_23489) );
na02m02 TIMEBOOST_cell_49644 ( .a(TIMEBOOST_net_15039), .b(g61782_sb), .o(n_8241) );
na03f02 TIMEBOOST_cell_65681 ( .a(TIMEBOOST_net_20388), .b(FE_OFN2128_n_16497), .c(g54309_sb), .o(n_13022) );
na02s01 TIMEBOOST_cell_68428 ( .a(g58161_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q), .o(TIMEBOOST_net_21422) );
na02s01 TIMEBOOST_cell_42772 ( .a(TIMEBOOST_net_12280), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_387), .o(n_13166) );
na02s01 TIMEBOOST_cell_39771 ( .a(TIMEBOOST_net_11497), .b(g58133_db), .o(n_9072) );
na02f02 TIMEBOOST_cell_42816 ( .a(TIMEBOOST_net_12302), .b(g67040_sb), .o(n_1502) );
na02m02 TIMEBOOST_cell_39665 ( .a(TIMEBOOST_net_11444), .b(g63132_sb), .o(n_4986) );
na02m02 TIMEBOOST_cell_38796 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q), .b(g63566_sb), .o(TIMEBOOST_net_11010) );
in01s01 TIMEBOOST_cell_67793 ( .a(pci_target_unit_fifos_pcir_data_in_160), .o(TIMEBOOST_net_21220) );
na02s01 TIMEBOOST_cell_62944 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q), .b(FE_OFN258_n_9862), .o(TIMEBOOST_net_20419) );
na02f02 TIMEBOOST_cell_38798 ( .a(g58407_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q), .o(TIMEBOOST_net_11011) );
na03s02 TIMEBOOST_cell_64439 ( .a(TIMEBOOST_net_12833), .b(g61964_db), .c(g63597_sb), .o(TIMEBOOST_net_16381) );
na02s01 TIMEBOOST_cell_38800 ( .a(TIMEBOOST_net_7108), .b(FE_OFN776_n_15366), .o(TIMEBOOST_net_11012) );
na02s02 TIMEBOOST_cell_42776 ( .a(TIMEBOOST_net_12282), .b(g65268_db), .o(TIMEBOOST_net_10171) );
na03f02 TIMEBOOST_cell_72914 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q), .b(g64304_sb), .c(TIMEBOOST_net_22102), .o(TIMEBOOST_net_20924) );
na02m02 TIMEBOOST_cell_68769 ( .a(TIMEBOOST_net_21592), .b(TIMEBOOST_net_16201), .o(TIMEBOOST_net_17017) );
in01m01 g65931_u0 ( .a(FE_OFN614_n_4501), .o(g65931_sb) );
na02s02 TIMEBOOST_cell_68627 ( .a(TIMEBOOST_net_21521), .b(FE_OFN1015_n_2053), .o(TIMEBOOST_net_20378) );
na03f02 TIMEBOOST_cell_34794 ( .a(TIMEBOOST_net_9545), .b(FE_OFN1380_n_8567), .c(g57512_sb), .o(n_10319) );
no02f01 g65932_u0 ( .a(n_2171), .b(n_2044), .o(g65932_p) );
ao12f01 g65932_u1 ( .a(g65932_p), .b(n_2171), .c(n_2044), .o(n_2172) );
na02f02 TIMEBOOST_cell_50446 ( .a(TIMEBOOST_net_15440), .b(g62344_sb), .o(n_6911) );
na02s02 TIMEBOOST_cell_70466 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q), .b(FE_OFN603_n_9687), .o(TIMEBOOST_net_22441) );
na03m04 TIMEBOOST_cell_73142 ( .a(FE_OFN1077_n_4740), .b(TIMEBOOST_net_17276), .c(g64080_sb), .o(n_4075) );
in01f01 g65934_u0 ( .a(FE_OFN959_n_2299), .o(g65934_sb) );
na02f01 TIMEBOOST_cell_63877 ( .a(TIMEBOOST_net_20924), .b(FE_OFN1134_g64577_p), .o(TIMEBOOST_net_15194) );
na02f02 g65934_u2 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(FE_OFN959_n_2299), .o(g65934_db) );
in01m01 g65935_u0 ( .a(FE_OFN959_n_2299), .o(g65935_sb) );
na03f02 TIMEBOOST_cell_68031 ( .a(TIMEBOOST_net_17387), .b(FE_OFN1212_n_4151), .c(g63184_sb), .o(n_5784) );
na02m10 TIMEBOOST_cell_45263 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q), .o(TIMEBOOST_net_13526) );
na02m02 TIMEBOOST_cell_44427 ( .a(n_4726), .b(n_271), .o(TIMEBOOST_net_13108) );
in01f02 g65936_u0 ( .a(FE_OFN948_n_2248), .o(g65936_sb) );
na02f02 g65936_u1 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q), .b(g65936_sb), .o(g65936_da) );
na02m02 g65936_u2 ( .a(pci_target_unit_fifos_pcir_data_in_162), .b(FE_OFN948_n_2248), .o(g65936_db) );
na02f04 g65936_u3 ( .a(g65936_da), .b(g65936_db), .o(n_1564) );
no02f01 g65937_u0 ( .a(n_2376), .b(FE_OCPN1854_n_2071), .o(g65937_p) );
ao12f01 g65937_u1 ( .a(g65937_p), .b(n_2376), .c(FE_OCPN1854_n_2071), .o(n_2377) );
no02f01 g65938_u0 ( .a(n_1847), .b(n_1698), .o(g65938_p) );
ao12f01 g65938_u1 ( .a(g65938_p), .b(n_1847), .c(n_1698), .o(n_1848) );
no02f01 g65939_u0 ( .a(n_2566), .b(n_1061), .o(g65939_p) );
ao12f01 g65939_u1 ( .a(g65939_p), .b(n_2566), .c(n_1061), .o(n_2580) );
in01m01 g65940_u0 ( .a(n_2301), .o(g65940_sb) );
na03f02 TIMEBOOST_cell_72987 ( .a(configuration_wb_err_addr_547), .b(n_5633), .c(TIMEBOOST_net_20441), .o(n_5580) );
na02s01 g65940_u2 ( .a(n_8511), .b(n_2301), .o(g65940_db) );
na03m08 TIMEBOOST_cell_72988 ( .a(FE_OFN1050_n_16657), .b(TIMEBOOST_net_16314), .c(g64215_sb), .o(n_3954) );
na04m20 TIMEBOOST_cell_67120 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q), .b(pci_target_unit_fifos_pcir_flush_in), .c(g57780_sb), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q), .o(TIMEBOOST_net_15866) );
na03f02 TIMEBOOST_cell_73431 ( .a(TIMEBOOST_net_20578), .b(FE_OFN1197_n_4090), .c(g62613_sb), .o(n_6331) );
na03f02 TIMEBOOST_cell_34993 ( .a(TIMEBOOST_net_9569), .b(g57291_sb), .c(FE_OFN2191_n_8567), .o(n_11462) );
in01m01 g65942_u0 ( .a(FE_OFN2111_n_2248), .o(g65942_sb) );
na04f04 TIMEBOOST_cell_73332 ( .a(n_3858), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q), .c(FE_OFN1131_g64577_p), .d(g63111_sb), .o(n_5033) );
na02m01 g65942_u2 ( .a(pci_target_unit_fifos_pcir_data_in_181), .b(FE_OFN2111_n_2248), .o(g65942_db) );
in01s01 g65943_u0 ( .a(FE_OFN1044_n_2037), .o(g65943_sb) );
na02m02 TIMEBOOST_cell_68123 ( .a(TIMEBOOST_net_21269), .b(g61943_sb), .o(TIMEBOOST_net_17286) );
na03f02 TIMEBOOST_cell_72672 ( .a(TIMEBOOST_net_6912), .b(g52647_sb), .c(FE_OCPUNCON1952_FE_OFN697_n_16760), .o(n_14741) );
na03m01 TIMEBOOST_cell_73065 ( .a(TIMEBOOST_net_14596), .b(FE_OFN2258_n_8060), .c(g61809_sb), .o(n_8175) );
na03f02 TIMEBOOST_cell_73649 ( .a(TIMEBOOST_net_9955), .b(FE_OFN1236_n_6391), .c(g62627_sb), .o(n_6301) );
na02s02 TIMEBOOST_cell_49250 ( .a(TIMEBOOST_net_14842), .b(TIMEBOOST_net_10860), .o(TIMEBOOST_net_9409) );
na02m02 TIMEBOOST_cell_69117 ( .a(TIMEBOOST_net_21766), .b(g65379_sb), .o(TIMEBOOST_net_16255) );
na03f01 TIMEBOOST_cell_68114 ( .a(TIMEBOOST_net_13996), .b(FE_OFN1818_i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q), .o(TIMEBOOST_net_21265) );
na02s01 g65946_u2 ( .a(n_2648), .b(n_2301), .o(g65946_db) );
na02m02 TIMEBOOST_cell_49636 ( .a(TIMEBOOST_net_15035), .b(g62024_sb), .o(n_7849) );
na02f06 TIMEBOOST_cell_68205 ( .a(TIMEBOOST_net_21310), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q), .o(TIMEBOOST_net_16143) );
na02s01 TIMEBOOST_cell_42778 ( .a(TIMEBOOST_net_12283), .b(g58774_da), .o(n_9889) );
no03f06 TIMEBOOST_cell_67022 ( .a(FE_RN_827_0), .b(FE_RN_828_0), .c(FE_RN_829_0), .o(n_14402) );
na02m01 TIMEBOOST_cell_62508 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q), .b(pci_target_unit_fifos_pcir_control_in_192), .o(TIMEBOOST_net_20201) );
na03f02 TIMEBOOST_cell_66164 ( .a(TIMEBOOST_net_17001), .b(FE_OFN1182_n_3476), .c(g60637_sb), .o(n_5696) );
in01m01 g65949_u0 ( .a(FE_OFN948_n_2248), .o(g65949_sb) );
na04f04 TIMEBOOST_cell_24794 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q), .b(g58808_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q), .d(FE_OFN2153_n_16439), .o(n_8633) );
na03m04 TIMEBOOST_cell_72989 ( .a(TIMEBOOST_net_21995), .b(FE_OFN1051_n_16657), .c(TIMEBOOST_net_23260), .o(TIMEBOOST_net_21062) );
na04f04 TIMEBOOST_cell_24795 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q), .b(g58807_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q), .d(FE_OFN2153_n_16439), .o(n_8634) );
na03m02 TIMEBOOST_cell_295 ( .a(n_2174), .b(g61735_sb), .c(g61996_db), .o(n_7903) );
na02m01 TIMEBOOST_cell_71880 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q), .b(FE_OFN670_n_4505), .o(TIMEBOOST_net_23148) );
in01s01 g65951_u0 ( .a(n_2299), .o(g65951_sb) );
na02s01 TIMEBOOST_cell_45421 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q), .o(TIMEBOOST_net_13605) );
na02s01 g65951_u2 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(n_2299), .o(g65951_db) );
na02f02 TIMEBOOST_cell_45422 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13605), .o(TIMEBOOST_net_12035) );
in01s01 g65952_u0 ( .a(FE_OFN1015_n_2053), .o(g65952_sb) );
na02s06 TIMEBOOST_cell_47555 ( .a(wbs_dat_i_25_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q), .o(TIMEBOOST_net_13995) );
na02s01 g65952_u2 ( .a(pci_target_unit_fifos_pcir_data_in_177), .b(FE_OFN1015_n_2053), .o(g65952_db) );
na02m04 TIMEBOOST_cell_70764 ( .a(wbm_adr_o_25_), .b(g59231_sb), .o(TIMEBOOST_net_22590) );
in01f02 g65953_u0 ( .a(FE_OFN1797_n_2299), .o(g65953_sb) );
na03f02 TIMEBOOST_cell_66502 ( .a(TIMEBOOST_net_17107), .b(FE_OFN1312_n_6624), .c(g62961_sb), .o(n_5960) );
na03f02 TIMEBOOST_cell_73742 ( .a(TIMEBOOST_net_13676), .b(n_11831), .c(FE_OCP_RBN1973_n_12381), .o(n_12665) );
na02m02 TIMEBOOST_cell_54632 ( .a(TIMEBOOST_net_17533), .b(FE_OFN1295_n_4098), .o(TIMEBOOST_net_15446) );
in01s01 g65954_u0 ( .a(FE_OFN1015_n_2053), .o(g65954_sb) );
na02f01 TIMEBOOST_cell_70570 ( .a(TIMEBOOST_net_15103), .b(FE_OFN882_g64577_p), .o(TIMEBOOST_net_22493) );
na02s01 TIMEBOOST_cell_42784 ( .a(TIMEBOOST_net_12286), .b(n_8832), .o(n_9228) );
na02m02 TIMEBOOST_cell_68125 ( .a(TIMEBOOST_net_21270), .b(g54171_sb), .o(TIMEBOOST_net_12276) );
na03s02 TIMEBOOST_cell_64934 ( .a(g65741_db), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q), .c(TIMEBOOST_net_8236), .o(TIMEBOOST_net_12830) );
in01m01 g65957_u0 ( .a(n_2299), .o(g65957_sb) );
na02f01 g65957_u2 ( .a(pci_target_unit_fifos_pcir_data_in_170), .b(n_2299), .o(g65957_db) );
na02s01 TIMEBOOST_cell_45423 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q), .o(TIMEBOOST_net_13606) );
in01m01 g65958_u0 ( .a(n_2299), .o(g65958_sb) );
na03s01 TIMEBOOST_cell_46503 ( .a(TIMEBOOST_net_12574), .b(FE_OFN227_n_9841), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q), .o(TIMEBOOST_net_9390) );
na02m01 g65958_u2 ( .a(pci_target_unit_fifos_pcir_data_in_171), .b(n_2299), .o(g65958_db) );
na03f02 TIMEBOOST_cell_66626 ( .a(TIMEBOOST_net_9193), .b(FE_OCPN1847_n_14981), .c(g59090_sb), .o(n_8714) );
na02m01 g65959_u2 ( .a(pci_target_unit_fifos_pcir_data_in_173), .b(n_2299), .o(g65959_db) );
na02m02 TIMEBOOST_cell_68994 ( .a(g64858_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q), .o(TIMEBOOST_net_21705) );
in01s01 g65960_u0 ( .a(n_2299), .o(g65960_sb) );
na04f02 TIMEBOOST_cell_73432 ( .a(n_4914), .b(FE_OFN1222_n_6391), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q), .d(g62479_sb), .o(n_7383) );
na02m01 g65960_u2 ( .a(pci_target_unit_fifos_pcir_data_in_174), .b(n_2299), .o(g65960_db) );
no03f02 TIMEBOOST_cell_67024 ( .a(n_12816), .b(n_12920), .c(n_12707), .o(FE_RN_23_0) );
na04f04 TIMEBOOST_cell_24205 ( .a(n_9513), .b(g57428_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q), .d(FE_OFN1384_n_8567), .o(n_11306) );
na02s01 g65961_u2 ( .a(pci_target_unit_fifos_pcir_data_in_175), .b(n_2299), .o(g65961_db) );
in01m01 g65962_u0 ( .a(FE_OFN959_n_2299), .o(g65962_sb) );
na02m01 g65962_u2 ( .a(pci_target_unit_fifos_pcir_data_in_176), .b(FE_OFN959_n_2299), .o(g65962_db) );
na03f02 TIMEBOOST_cell_73765 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q), .b(FE_OFN1774_n_13800), .c(TIMEBOOST_net_12228), .o(n_16233) );
na02s01 TIMEBOOST_cell_42786 ( .a(TIMEBOOST_net_12287), .b(FE_OFN945_n_2248), .o(TIMEBOOST_net_10228) );
in01s01 g65964_u0 ( .a(n_2299), .o(g65964_sb) );
na03m06 TIMEBOOST_cell_69868 ( .a(FE_OFN1056_n_4727), .b(TIMEBOOST_net_16609), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q), .o(TIMEBOOST_net_22142) );
in01f02 g65965_u0 ( .a(FE_OFN1797_n_2299), .o(g65965_sb) );
in01f02 g65966_u0 ( .a(FE_OFN1797_n_2299), .o(g65966_sb) );
na03s01 TIMEBOOST_cell_64406 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q), .b(FE_OFN603_n_9687), .c(FE_OFN229_n_9120), .o(TIMEBOOST_net_16673) );
na03f02 TIMEBOOST_cell_47375 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_13686), .c(FE_OFN1581_n_12306), .o(n_12498) );
in01f01 g65967_u0 ( .a(FE_OFN1797_n_2299), .o(g65967_sb) );
na02m02 g65967_u2 ( .a(TIMEBOOST_net_21129), .b(FE_OFN1797_n_2299), .o(g65967_db) );
in01s01 TIMEBOOST_cell_63557 ( .a(TIMEBOOST_net_20737), .o(TIMEBOOST_net_20736) );
na02s01 TIMEBOOST_cell_42788 ( .a(TIMEBOOST_net_12288), .b(FE_OFN945_n_2248), .o(TIMEBOOST_net_140) );
na02m02 g65968_u2 ( .a(pci_target_unit_del_sync_addr_in_220), .b(FE_OFN776_n_15366), .o(g65968_db) );
na02m02 TIMEBOOST_cell_68714 ( .a(n_3783), .b(n_119), .o(TIMEBOOST_net_21565) );
in01f02 g65969_u0 ( .a(FE_OFN1797_n_2299), .o(g65969_sb) );
na02m02 TIMEBOOST_cell_53376 ( .a(TIMEBOOST_net_16905), .b(FE_OFN789_n_2678), .o(TIMEBOOST_net_14536) );
in01f01 g65970_u0 ( .a(FE_OFN1797_n_2299), .o(g65970_sb) );
na03f04 TIMEBOOST_cell_73478 ( .a(wbm_adr_o_19_), .b(g61856_sb), .c(g52395_sb), .o(TIMEBOOST_net_22956) );
na03s04 TIMEBOOST_cell_72604 ( .a(FE_OFN1650_n_9428), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q), .c(FE_OFN241_n_9830), .o(TIMEBOOST_net_12811) );
in01f04 g65971_u0 ( .a(FE_OFN1797_n_2299), .o(g65971_sb) );
na03f02 TIMEBOOST_cell_66625 ( .a(TIMEBOOST_net_17053), .b(n_6232), .c(g62630_sb), .o(n_6295) );
na02s02 TIMEBOOST_cell_70413 ( .a(TIMEBOOST_net_22414), .b(g58429_sb), .o(n_9418) );
na03f02 TIMEBOOST_cell_47377 ( .a(FE_OFN1759_n_10780), .b(TIMEBOOST_net_13682), .c(FE_OFN1581_n_12306), .o(n_12493) );
in01f01 g65972_u0 ( .a(FE_OFN1797_n_2299), .o(g65972_sb) );
na02m02 TIMEBOOST_cell_49116 ( .a(TIMEBOOST_net_14775), .b(g61862_sb), .o(n_8114) );
na02f02 TIMEBOOST_cell_70351 ( .a(TIMEBOOST_net_22383), .b(g63016_sb), .o(n_5216) );
na02s02 TIMEBOOST_cell_68262 ( .a(g65775_sb), .b(TIMEBOOST_net_21141), .o(TIMEBOOST_net_21339) );
na04m04 TIMEBOOST_cell_73275 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q), .b(FE_OFN1812_n_7845), .c(n_1608), .d(g61817_sb), .o(n_8157) );
na03f02 TIMEBOOST_cell_69460 ( .a(TIMEBOOST_net_21157), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q), .c(g65969_sb), .o(TIMEBOOST_net_21938) );
na03f02 TIMEBOOST_cell_72228 ( .a(TIMEBOOST_net_20890), .b(FE_OFN1670_n_9477), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q), .o(TIMEBOOST_net_23322) );
in01s01 g65976_u0 ( .a(FE_OFN1017_n_2053), .o(g65976_sb) );
na02m06 TIMEBOOST_cell_45343 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q), .o(TIMEBOOST_net_13566) );
na03f02 TIMEBOOST_cell_72535 ( .a(TIMEBOOST_net_14194), .b(FE_OFN918_n_4725), .c(TIMEBOOST_net_23172), .o(TIMEBOOST_net_17320) );
in01s01 g65977_u0 ( .a(FE_OFN1015_n_2053), .o(g65977_sb) );
in01s01 TIMEBOOST_cell_67739 ( .a(pci_target_unit_fifos_pcir_data_in_173), .o(TIMEBOOST_net_21166) );
in01s01 g65978_u0 ( .a(FE_OFN1015_n_2053), .o(g65978_sb) );
na03f02 TIMEBOOST_cell_66935 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_16503), .c(FE_OFN2210_n_11027), .o(n_12729) );
in01s01 TIMEBOOST_cell_63600 ( .a(TIMEBOOST_net_20780), .o(TIMEBOOST_net_20715) );
ao12f40 g65981_u0 ( .a(n_313), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_), .o(n_938) );
no02m06 g65983_u0 ( .a(pci_target_unit_fifos_wb_clk_inGreyCount_1_), .b(pci_target_unit_fifos_outGreyCount_reg_1__Q), .o(g65983_p) );
ao12m08 g65983_u1 ( .a(g65983_p), .b(pci_target_unit_fifos_wb_clk_inGreyCount_1_), .c(pci_target_unit_fifos_outGreyCount_reg_1__Q), .o(n_1834) );
no02f10 g65984_u0 ( .a(n_202), .b(pci_target_unit_fifos_wb_clk_inGreyCount_0_), .o(g65984_p) );
ao12f06 g65984_u1 ( .a(g65984_p), .b(pci_target_unit_fifos_wb_clk_inGreyCount_0_), .c(n_202), .o(n_1832) );
na03f02 TIMEBOOST_cell_73529 ( .a(TIMEBOOST_net_17481), .b(FE_OFN1244_n_4092), .c(g62710_sb), .o(n_6150) );
no02s01 g65992_u0 ( .a(n_1847), .b(n_2376), .o(g65992_p) );
ao12s01 g65992_u1 ( .a(g65992_p), .b(n_1847), .c(n_2376), .o(n_1407) );
no02f01 g65993_u0 ( .a(n_2566), .b(n_2171), .o(g65993_p) );
ao12f01 g65993_u1 ( .a(g65993_p), .b(n_2566), .c(n_2171), .o(n_1406) );
in01f04 g65994_u0 ( .a(FE_OFN992_n_2373), .o(g65994_sb) );
na03f02 TIMEBOOST_cell_34841 ( .a(TIMEBOOST_net_9469), .b(FE_OFN1401_n_8567), .c(g57127_sb), .o(n_11618) );
na02f02 TIMEBOOST_cell_45424 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13606), .o(TIMEBOOST_net_12037) );
na02f01 g65995_u1 ( .a(g65994_sb), .b(wbu_pciif_devsel_reg_in), .o(g65995_da) );
na03s01 TIMEBOOST_cell_64325 ( .a(TIMEBOOST_net_13984), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_409), .c(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q), .o(TIMEBOOST_net_17568) );
na02s01 TIMEBOOST_cell_45425 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q), .o(TIMEBOOST_net_13607) );
na02f01 g65996_u1 ( .a(n_15302), .b(g65994_sb), .o(g65996_da) );
na02s01 g65996_u2 ( .a(n_1551), .b(FE_OFN992_n_2373), .o(g65996_db) );
na02f01 g65996_u3 ( .a(g65996_da), .b(g65996_db), .o(n_2372) );
na03s02 TIMEBOOST_cell_41805 ( .a(TIMEBOOST_net_10566), .b(g58451_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q), .o(TIMEBOOST_net_9566) );
na04f04 TIMEBOOST_cell_42525 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_774), .c(FE_OFN2135_n_13124), .d(g54369_sb), .o(n_13074) );
na02s01 TIMEBOOST_cell_48892 ( .a(TIMEBOOST_net_14663), .b(g57947_sb), .o(TIMEBOOST_net_10827) );
na03m08 TIMEBOOST_cell_64324 ( .a(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q), .b(n_13447), .c(wishbone_slave_unit_pcim_if_wbw_addr_data_in_398), .o(TIMEBOOST_net_16950) );
na03f02 TIMEBOOST_cell_73276 ( .a(TIMEBOOST_net_23319), .b(FE_OFN1174_n_5592), .c(g62113_sb), .o(n_5583) );
na02f01 TIMEBOOST_cell_47958 ( .a(TIMEBOOST_net_14196), .b(FE_OFN918_n_4725), .o(TIMEBOOST_net_12496) );
na02s01 TIMEBOOST_cell_53596 ( .a(TIMEBOOST_net_17015), .b(g58347_sb), .o(n_9474) );
na02f01 TIMEBOOST_cell_44248 ( .a(TIMEBOOST_net_13018), .b(FE_OFN1100_g64577_p), .o(TIMEBOOST_net_11170) );
na03m02 TIMEBOOST_cell_72812 ( .a(TIMEBOOST_net_21546), .b(g64935_sb), .c(TIMEBOOST_net_21839), .o(TIMEBOOST_net_17414) );
na04f04 TIMEBOOST_cell_42513 ( .a(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q), .b(pci_target_unit_pcit_if_pcir_fifo_data_in_773), .c(FE_OFN2135_n_13124), .d(g54368_sb), .o(n_13075) );
na03f02 TIMEBOOST_cell_34777 ( .a(TIMEBOOST_net_9366), .b(FE_OFN1409_n_8567), .c(g57132_sb), .o(n_11616) );
na02f01 g66001_u2 ( .a(n_1450), .b(FE_OFN992_n_2373), .o(g66001_db) );
na02m02 TIMEBOOST_cell_68925 ( .a(TIMEBOOST_net_21670), .b(g65072_db), .o(TIMEBOOST_net_17461) );
no02f20 g66002_u0 ( .a(n_595), .b(n_585), .o(g66002_p) );
ao12f10 g66002_u1 ( .a(g66002_p), .b(n_595), .c(n_585), .o(n_1405) );
no02f20 g66003_u0 ( .a(n_674), .b(n_598), .o(g66003_p) );
ao12f10 g66003_u1 ( .a(g66003_p), .b(n_674), .c(n_598), .o(n_1404) );
no02f20 g66004_u0 ( .a(n_672), .b(n_592), .o(g66004_p) );
ao12f20 g66004_u1 ( .a(g66004_p), .b(n_672), .c(n_592), .o(n_1403) );
no02f20 g66005_u0 ( .a(n_597), .b(n_663), .o(g66005_p) );
ao12f10 g66005_u1 ( .a(g66005_p), .b(n_597), .c(n_663), .o(n_1402) );
no02f20 g66006_u0 ( .a(n_678), .b(n_664), .o(g66006_p) );
ao12f10 g66006_u1 ( .a(g66006_p), .b(n_678), .c(n_664), .o(n_1401) );
no02f20 g66007_u0 ( .a(n_586), .b(n_584), .o(g66007_p) );
ao12f10 g66007_u1 ( .a(g66007_p), .b(n_586), .c(n_584), .o(n_1449) );
no02f20 g66008_u0 ( .a(n_603), .b(n_666), .o(g66008_p) );
ao12f10 g66008_u1 ( .a(g66008_p), .b(n_603), .c(n_666), .o(n_1400) );
no02f10 g66009_u0 ( .a(n_593), .b(n_656), .o(g66009_p) );
ao12f10 g66009_u1 ( .a(g66009_p), .b(n_593), .c(n_656), .o(n_1399) );
no02f20 g66010_u0 ( .a(n_667), .b(n_605), .o(g66010_p) );
ao12f10 g66010_u1 ( .a(g66010_p), .b(n_667), .c(n_605), .o(n_1398) );
no02f10 g66011_u0 ( .a(n_670), .b(n_652), .o(g66011_p) );
ao12f10 g66011_u1 ( .a(g66011_p), .b(n_670), .c(n_652), .o(n_1397) );
no02f20 g66012_u0 ( .a(n_650), .b(n_581), .o(g66012_p) );
ao12f10 g66012_u1 ( .a(g66012_p), .b(n_650), .c(n_581), .o(n_1396) );
no02f20 g66013_u0 ( .a(n_583), .b(n_606), .o(g66013_p) );
ao12f10 g66013_u1 ( .a(g66013_p), .b(n_606), .c(n_583), .o(n_1395) );
no02f20 g66014_u0 ( .a(n_673), .b(n_600), .o(g66014_p) );
ao12f10 g66014_u1 ( .a(g66014_p), .b(n_673), .c(n_600), .o(n_1439) );
no02f08 g66015_u0 ( .a(n_594), .b(n_677), .o(g66015_p) );
ao12f08 g66015_u1 ( .a(g66015_p), .b(n_677), .c(n_594), .o(n_1394) );
no02f20 g66016_u0 ( .a(n_675), .b(n_607), .o(g66016_p) );
ao12f10 g66016_u1 ( .a(g66016_p), .b(n_675), .c(n_607), .o(n_1393) );
na02m02 TIMEBOOST_cell_51853 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q), .b(TIMEBOOST_net_12368), .o(TIMEBOOST_net_16144) );
no02f40 g66065_u0 ( .a(n_1477), .b(n_208), .o(n_1985) );
na02f10 g66066_u0 ( .a(n_1361), .b(wbu_addr_in_251), .o(g66066_p) );
in01f10 g66066_u1 ( .a(g66066_p), .o(n_2225) );
in01f02 g66067_u0 ( .a(n_1965), .o(n_1561) );
na02f10 g66068_u0 ( .a(n_1357), .b(conf_wb_err_addr_in_943), .o(g66068_p) );
in01f10 g66068_u1 ( .a(g66068_p), .o(n_1965) );
na02m02 TIMEBOOST_cell_69022 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q), .b(FE_OFN614_n_4501), .o(TIMEBOOST_net_21719) );
na02m01 g66070_u0 ( .a(n_3030), .b(n_2301), .o(n_3217) );
na02m01 g66071_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1213), .o(n_2612) );
no02m04 g66072_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1208), .o(g66072_p) );
in01m08 g66072_u1 ( .a(g66072_p), .o(n_4498) );
na02f01 g66073_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1212), .o(n_2610) );
no02m04 g66074_u0 ( .a(parchk_pci_ad_reg_in_1206), .b(n_2493), .o(g66074_p) );
in01m08 g66074_u1 ( .a(g66074_p), .o(n_4672) );
no02f04 g66075_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1233), .o(g66075_p) );
in01f08 g66075_u1 ( .a(g66075_p), .o(n_4479) );
no02f02 g66076_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in), .o(g66076_p) );
in01f06 g66076_u1 ( .a(g66076_p), .o(n_4488) );
no02m02 g66077_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1214), .o(g66077_p) );
in01m06 g66077_u1 ( .a(g66077_p), .o(n_3747) );
no02m04 g66078_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1212), .o(g66078_p) );
in01m08 g66078_u1 ( .a(g66078_p), .o(n_4465) );
no02f01 g66079_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1211), .o(g66079_p) );
in01f04 g66079_u1 ( .a(g66079_p), .o(n_3764) );
no02m06 g66080_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1228), .o(g66080_p) );
in01m08 g66080_u1 ( .a(g66080_p), .o(n_4444) );
no02f01 g66081_u0 ( .a(n_2509), .b(n_2344), .o(g66081_p) );
in01f10 g66081_u1 ( .a(FE_OFN335_g66081_p), .o(n_3770) );
no02f01 g66082_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1213), .o(g66082_p) );
in01f04 g66082_u1 ( .a(g66082_p), .o(n_3783) );
na02f08 g66083_u0 ( .a(n_15922), .b(n_2308), .o(g66083_p) );
in01f06 g66083_u1 ( .a(g66083_p), .o(n_2562) );
no02f02 g66084_u0 ( .a(n_1122), .b(wishbone_slave_unit_del_sync_comp_cycle_count_10_), .o(g66084_p) );
in01f02 g66084_u1 ( .a(g66084_p), .o(n_1392) );
no02m01 g66085_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1229), .o(g66085_p) );
in01f10 g66085_u1 ( .a(FE_OFN1938_g66085_p), .o(n_3785) );
no02m04 g66086_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1235), .o(g66086_p) );
in01m08 g66086_u1 ( .a(g66086_p), .o(n_4645) );
no02m02 g66087_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1216), .o(g66087_p) );
in01m10 g66087_u1 ( .a(FE_OFN2061_g66087_p), .o(n_3777) );
na02f01 g66088_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1209), .o(n_2604) );
no02m02 g66089_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1205), .o(g66089_p) );
in01m10 g66089_u1 ( .a(FE_OFN337_g66089_p), .o(n_3774) );
no02f06 g66090_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1223), .o(g66090_p) );
in01f08 g66090_u1 ( .a(g66090_p), .o(n_4447) );
na02f01 g66092_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1207), .o(n_2788) );
no02m04 g66093_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1225), .o(g66093_p) );
in01m08 g66093_u1 ( .a(g66093_p), .o(n_4470) );
no02m04 g66094_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1217), .o(g66094_p) );
in01m08 g66094_u1 ( .a(g66094_p), .o(n_4452) );
no02m02 g66095_u0 ( .a(FE_OFN1781_parchk_pci_ad_reg_in_1221), .b(n_2493), .o(g66095_p) );
in01f08 g66095_u1 ( .a(FE_OFN1940_g66095_p), .o(n_4450) );
na02f02 g66096_u0 ( .a(n_1478), .b(n_1479), .o(g66096_p) );
in01f04 g66096_u1 ( .a(g66096_p), .o(n_2244) );
na02f10 g66097_u0 ( .a(n_2967), .b(n_1390), .o(g66097_p) );
in01f08 g66097_u1 ( .a(g66097_p), .o(n_1391) );
no02m02 g66098_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1220), .o(g66098_p) );
in01m06 g66098_u1 ( .a(g66098_p), .o(n_3744) );
na02f06 g66099_u0 ( .a(n_1378), .b(n_1480), .o(g66099_p) );
in01f04 g66099_u1 ( .a(g66099_p), .o(n_2243) );
no02f04 g66100_u0 ( .a(parchk_pci_ad_reg_in_1232), .b(n_2493), .o(g66100_p) );
in01f08 g66100_u1 ( .a(g66100_p), .o(n_4442) );
in01s01 g66105_u0 ( .a(n_3123), .o(n_2140) );
na02f40 g66106_u0 ( .a(n_1196), .b(pci_target_unit_pci_target_sm_backoff), .o(n_3123) );
no02m02 g66107_u0 ( .a(parchk_pci_ad_reg_in_1210), .b(n_2344), .o(g66107_p) );
in01f06 g66107_u1 ( .a(g66107_p), .o(n_3780) );
no02m04 g66108_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1218), .o(g66108_p) );
in01m08 g66108_u1 ( .a(g66108_p), .o(n_4476) );
na02m01 g66109_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1206), .o(n_2790) );
no02m02 g66110_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1207), .o(g66110_p) );
in01m06 g66110_u1 ( .a(g66110_p), .o(n_3739) );
na02f01 g66111_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1208), .o(n_2732) );
na02s01 g66112_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1210), .o(n_2783) );
na02f20 g66113_u0 ( .a(n_1482), .b(n_1481), .o(g66113_p) );
in01f10 g66113_u1 ( .a(g66113_p), .o(n_2397) );
no02f04 g66114_u0 ( .a(n_639), .b(n_1057), .o(n_2675) );
na02m01 g66117_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1211), .o(n_2606) );
no02f04 g66118_u0 ( .a(n_207), .b(n_1124), .o(g66118_p) );
in01f02 g66118_u1 ( .a(g66118_p), .o(n_1389) );
na02m01 g66119_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in_1205), .o(n_2779) );
no02f20 g66120_u0 ( .a(n_1435), .b(n_978), .o(n_2415) );
na02f10 g66121_u0 ( .a(n_1388), .b(n_2435), .o(g66121_p) );
in01f08 g66121_u1 ( .a(g66121_p), .o(n_2229) );
no02s01 g66122_u0 ( .a(n_1824), .b(pci_target_unit_pcit_if_req_req_pending_in), .o(g66122_p) );
in01f01 g66122_u1 ( .a(g66122_p), .o(n_1825) );
na02m01 g66123_u0 ( .a(n_2301), .b(parchk_pci_ad_reg_in), .o(n_2601) );
no02m04 g66124_u0 ( .a(n_2493), .b(parchk_pci_ad_reg_in_1231), .o(g66124_p) );
in01m08 g66124_u1 ( .a(g66124_p), .o(n_4482) );
no02m02 g66125_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1215), .o(g66125_p) );
in01m06 g66125_u1 ( .a(g66125_p), .o(n_3761) );
no02m02 g66127_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1227), .o(g66127_p) );
in01m06 g66127_u1 ( .a(g66127_p), .o(n_3741) );
no02m02 g66128_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1226), .o(g66128_p) );
in01m06 g66128_u1 ( .a(g66128_p), .o(n_3749) );
no02m02 g66129_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1224), .o(g66129_p) );
in01m06 g66129_u1 ( .a(g66129_p), .o(n_3752) );
no02m02 g66130_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1219), .o(g66130_p) );
in01m06 g66130_u1 ( .a(g66130_p), .o(n_3792) );
na02f04 g66131_u0 ( .a(n_1125), .b(pci_target_unit_del_sync_comp_cycle_count_6_), .o(n_1484) );
no02f06 g66132_u0 ( .a(n_2215), .b(pci_target_unit_wishbone_master_first_wb_data_access), .o(g66132_p) );
in01f04 g66132_u1 ( .a(g66132_p), .o(n_2390) );
no02m02 g66133_u0 ( .a(n_2344), .b(parchk_pci_ad_reg_in_1209), .o(g66133_p) );
in01m06 g66133_u1 ( .a(g66133_p), .o(n_3755) );
no02f04 g66134_u0 ( .a(n_2493), .b(FE_OFN1777_parchk_pci_ad_reg_in_1222), .o(g66134_p) );
in01f08 g66134_u1 ( .a(g66134_p), .o(n_4473) );
na02m08 g66135_u0 ( .a(n_1123), .b(wishbone_slave_unit_del_sync_comp_cycle_count_6_), .o(n_1485) );
no02m04 g66136_u0 ( .a(parchk_pci_ad_reg_in_1230), .b(n_2493), .o(g66136_p) );
in01m08 g66136_u1 ( .a(g66136_p), .o(n_4493) );
no02f01 g66137_u0 ( .a(n_1192), .b(n_5757), .o(n_2303) );
na02f10 g66138_u0 ( .a(n_2411), .b(n_1227), .o(g66138_p) );
in01f08 g66138_u1 ( .a(g66138_p), .o(n_1986) );
no02f08 g66139_u0 ( .a(n_869), .b(n_1019), .o(n_1387) );
no02f06 g66140_u0 ( .a(n_642), .b(n_626), .o(n_1170) );
na02s02 TIMEBOOST_cell_71969 ( .a(TIMEBOOST_net_23192), .b(g58402_sb), .o(TIMEBOOST_net_10882) );
na02m01 g66142_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q), .b(FE_OFN614_n_4501), .o(n_1559) );
no02f04 g66143_u0 ( .a(n_15291), .b(n_2127), .o(g66143_p) );
in01f06 g66143_u1 ( .a(g66143_p), .o(n_3019) );
na02f10 g66145_u0 ( .a(n_1229), .b(n_1228), .o(g66145_p) );
in01f08 g66145_u1 ( .a(g66145_p), .o(n_2753) );
na02s01 g66146_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pci_target_sm_rd_progress), .o(n_1823) );
no02f20 g66147_u0 ( .a(n_604), .b(n_601), .o(g66147_p) );
in01f20 g66147_u1 ( .a(g66147_p), .o(n_1036) );
na02s01 g66148_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q), .b(FE_OFN1795_n_9904), .o(n_1230) );
na02s01 g66150_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pci_target_if_same_read_reg), .o(n_2371) );
no02f04 g66151_u0 ( .a(n_1091), .b(n_851), .o(n_1486) );
na02s01 g66152_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q), .b(FE_OFN1800_n_9690), .o(n_1822) );
no02s01 g66153_u0 ( .a(configuration_rst_inactive), .b(n_2373), .o(g66153_p) );
in01s01 g66153_u1 ( .a(g66153_p), .o(n_1385) );
na02s01 g66154_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q), .b(FE_OFN519_n_9697), .o(n_1821) );
na02f04 g66155_u0 ( .a(n_2331), .b(n_16541), .o(g66155_p) );
in01f04 g66155_u1 ( .a(g66155_p), .o(n_3371) );
na03f02 TIMEBOOST_cell_66322 ( .a(TIMEBOOST_net_17139), .b(n_6319), .c(g62475_sb), .o(n_6639) );
na02m01 g66158_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q), .b(FE_OFN672_n_4505), .o(n_1488) );
na02m01 g66159_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q), .b(FE_OFN665_n_4495), .o(n_2138) );
na02f02 g66160_u0 ( .a(n_2560), .b(n_2129), .o(g66160_p) );
in01f02 g66160_u1 ( .a(g66160_p), .o(n_3246) );
na02s01 g66161_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q), .b(FE_OFN529_n_9899), .o(n_1820) );
in01f02 g66162_u0 ( .a(FE_OFN780_n_2746), .o(n_2747) );
na03f02 TIMEBOOST_cell_66503 ( .a(TIMEBOOST_net_17142), .b(FE_OFN1323_n_6436), .c(g62960_sb), .o(n_5962) );
no02f08 g66164_u0 ( .a(n_620), .b(n_622), .o(n_1169) );
no02s02 g66165_u0 ( .a(n_15276), .b(n_16291), .o(g66165_p) );
in01f02 g66165_u1 ( .a(g66165_p), .o(n_1819) );
no02f06 g66166_u0 ( .a(n_729), .b(n_734), .o(n_1037) );
no02m02 g66167_u0 ( .a(n_1192), .b(FE_OFN999_n_15978), .o(n_2370) );
na03f02 TIMEBOOST_cell_66163 ( .a(TIMEBOOST_net_16439), .b(FE_OFN1186_n_3476), .c(g60668_sb), .o(n_5650) );
na02m06 g66169_u0 ( .a(FE_OFN923_n_4740), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q), .o(n_1815) );
na02s01 g66170_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pci_target_sm_rd_from_fifo), .o(n_2369) );
na02s01 g66171_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN595_n_9694), .o(n_1814) );
no02f40 g66172_u0 ( .a(n_1033), .b(n_863), .o(n_1231) );
no02m04 g66173_u0 ( .a(n_1551), .b(output_backup_trdy_out_reg_Q), .o(n_2137) );
na02s01 g66174_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pci_target_sm_wr_progress), .o(n_2367) );
no02f03 g66175_u0 ( .a(n_737), .b(n_640), .o(n_1168) );
no02f02 g66176_u0 ( .a(n_3480), .b(n_691), .o(g66176_p) );
in01f02 g66176_u1 ( .a(g66176_p), .o(n_1557) );
no02f06 g66177_u0 ( .a(n_708), .b(n_649), .o(n_1167) );
na02f40 g66178_u0 ( .a(n_1813), .b(n_1812), .o(g66178_p) );
in01f40 g66178_u1 ( .a(g66178_p), .o(n_2447) );
na02m01 g66179_u0 ( .a(n_424), .b(FE_OFN622_n_4409), .o(n_1555) );
na02s01 g66180_u0 ( .a(n_1023), .b(FE_OFN2214_n_15366), .o(n_2366) );
in01s01 g66182_u0 ( .a(n_1554), .o(n_13817) );
no02f20 g66184_u0 ( .a(n_1366), .b(pci_target_unit_pci_target_sm_backoff), .o(g66184_p) );
in01f10 g66184_u1 ( .a(g66184_p), .o(n_1554) );
na02s01 g66185_u0 ( .a(FE_OFN2214_n_15366), .b(n_2078), .o(n_2364) );
na02s01 g66187_u0 ( .a(n_922), .b(n_1383), .o(n_1384) );
na02f02 TIMEBOOST_cell_18608 ( .a(TIMEBOOST_net_5667), .b(n_8757), .o(g52403_db) );
na02s01 g66189_u0 ( .a(FE_OFN2214_n_15366), .b(n_15998), .o(n_2363) );
na02f02 g66190_u0 ( .a(n_3194), .b(n_1381), .o(g66190_p) );
in01f02 g66190_u1 ( .a(g66190_p), .o(n_2754) );
na02s01 g66191_u0 ( .a(FE_OFN2214_n_15366), .b(n_16690), .o(n_2362) );
no02f40 g66193_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_), .o(n_313) );
na02f02 g66194_u0 ( .a(wbu_wb_init_complete_in), .b(n_779), .o(g66194_p) );
in01f02 g66194_u1 ( .a(g66194_p), .o(n_2558) );
na02f06 g66195_u0 ( .a(n_1241), .b(n_2433), .o(g66195_p) );
in01f06 g66195_u1 ( .a(g66195_p), .o(n_2236) );
na02f04 g66197_u0 ( .a(n_1479), .b(n_1378), .o(g66197_p) );
in01f04 g66197_u1 ( .a(g66197_p), .o(n_1379) );
no02f04 g66200_u0 ( .a(n_1504), .b(n_695), .o(n_2136) );
na02m01 g66201_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q), .b(FE_OFN1660_n_4490), .o(n_1377) );
na02f20 g66202_u0 ( .a(n_1812), .b(n_2795), .o(g66202_p) );
in01f10 g66202_u1 ( .a(g66202_p), .o(n_3107) );
no02f08 g66203_u0 ( .a(n_1008), .b(n_864), .o(n_1252) );
na02s01 g66204_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q), .b(FE_OFN562_n_9895), .o(n_1493) );
na02s01 g66205_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_del_sync_bc_in), .o(n_2361) );
no02f08 g66206_u0 ( .a(n_951), .b(n_1035), .o(n_1253) );
no02f06 g66207_u0 ( .a(n_624), .b(n_613), .o(n_1166) );
na02m01 g66208_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q), .b(FE_OFN648_n_4497), .o(n_1553) );
na02s01 g66209_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(n_2359) );
na02s01 g66212_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q), .b(FE_OFN577_n_9902), .o(n_1810) );
na02s01 TIMEBOOST_cell_63255 ( .a(TIMEBOOST_net_20574), .b(TIMEBOOST_net_12788), .o(TIMEBOOST_net_9364) );
no02f08 g66214_u0 ( .a(n_625), .b(n_610), .o(n_1073) );
no02m02 g66215_u0 ( .a(n_2493), .b(n_3480), .o(g66215_p) );
in01m02 g66215_u1 ( .a(g66215_p), .o(n_3481) );
in01f08 g66216_u0 ( .a(n_1548), .o(n_1549) );
na02f10 g66217_u0 ( .a(n_1270), .b(n_1269), .o(n_1548) );
na02f08 g66219_u0 ( .a(n_1808), .b(n_16159), .o(n_1809) );
na02f10 g66221_u0 ( .a(n_16160), .b(n_16151), .o(n_2966) );
na02f08 g66223_u0 ( .a(wbs_cyc_i), .b(wbu_wb_init_complete_in), .o(g66223_p) );
in01f06 g66223_u1 ( .a(g66223_p), .o(n_2557) );
no02f06 g66224_u0 ( .a(n_616), .b(n_643), .o(n_1080) );
na02f10 g66225_u0 ( .a(n_1373), .b(n_1374), .o(n_1974) );
no02f04 g66226_u0 ( .a(n_615), .b(n_612), .o(n_1207) );
na02f02 g66227_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q), .b(FE_OFN1623_n_4438), .o(n_1547) );
no02s01 g66228_u0 ( .a(n_15371), .b(n_2134), .o(n_2135) );
in01m01 TIMEBOOST_cell_45957 ( .a(pci_target_unit_fifos_pcir_data_in_178), .o(TIMEBOOST_net_13918) );
na02f20 g66230_u0 ( .a(n_1445), .b(n_16160), .o(n_3341) );
no02f02 g66231_u0 ( .a(n_2036), .b(n_2297), .o(n_2556) );
no02f10 g66232_u0 ( .a(n_849), .b(n_850), .o(g66232_p) );
in01f08 g66232_u1 ( .a(g66232_p), .o(n_1371) );
na02m01 g66233_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q), .b(FE_OFN659_n_4392), .o(n_1546) );
na02f04 g66234_u0 ( .a(n_1282), .b(n_2431), .o(g66234_p) );
in01f04 g66234_u1 ( .a(g66234_p), .o(n_2238) );
no02f20 g66236_u0 ( .a(n_847), .b(n_858), .o(n_1369) );
na02f01 g66237_u0 ( .a(n_15065), .b(wbu_am1_in), .o(g66237_p) );
in01f02 g66237_u1 ( .a(g66237_p), .o(n_2358) );
na02f20 g66239_u0 ( .a(n_2463), .b(n_2596), .o(g66239_p) );
in01f10 g66239_u1 ( .a(g66239_p), .o(n_1969) );
na02s01 g66240_u0 ( .a(n_535), .b(n_1120), .o(n_1545) );
no02f08 g66241_u0 ( .a(n_1012), .b(n_867), .o(n_1365) );
na02s01 g66242_u0 ( .a(n_497), .b(FE_OFN2214_n_15366), .o(n_2356) );
na02s01 g66245_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q), .b(FE_OFN601_n_9687), .o(n_1806) );
no02f20 g66246_u0 ( .a(n_1031), .b(n_870), .o(n_1363) );
no02f08 g66247_u0 ( .a(n_645), .b(n_617), .o(n_1208) );
na02f04 g66248_u0 ( .a(n_1361), .b(n_1378), .o(g66248_p) );
in01f02 g66248_u1 ( .a(g66248_p), .o(n_1362) );
in01f02 g66250_u0 ( .a(n_1805), .o(n_2132) );
na04f04 TIMEBOOST_cell_24216 ( .a(n_9525), .b(g57414_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q), .d(FE_OFN1384_n_8567), .o(n_11328) );
no02s01 g66252_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pcit_if_req_req_pending_in), .o(n_2353) );
na02m02 g66253_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q), .b(FE_OFN903_n_4736), .o(n_1804) );
na02s01 g66254_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q), .b(FE_OFN531_n_9823), .o(n_1542) );
na02f01 g66255_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q), .b(FE_OFN1012_n_4734), .o(n_1803) );
na02m01 g66256_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q), .b(FE_OFN634_n_4454), .o(n_1642) );
na02f01 TIMEBOOST_cell_53545 ( .a(TIMEBOOST_net_13098), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_16990) );
na02s01 g66258_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pci_target_sm_wr_to_fifo), .o(n_2352) );
no02f06 g66259_u0 ( .a(n_722), .b(n_658), .o(n_1164) );
na02s01 g66260_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q), .b(n_4417), .o(n_2131) );
no02m02 g66261_u0 ( .a(FE_OFN996_n_15366), .b(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q), .o(n_1802) );
na02s01 g66262_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q), .b(FE_OFN554_n_9864), .o(n_1800) );
no02f04 g66264_u0 ( .a(n_641), .b(n_614), .o(n_1209) );
na02s01 g66265_u0 ( .a(FE_OFN996_n_15366), .b(n_2314), .o(n_2351) );
na02f01 g66266_u0 ( .a(FE_OFN996_n_15366), .b(pci_target_unit_pci_target_if_norm_prf_en), .o(n_2350) );
na02f06 g66267_u0 ( .a(n_965), .b(n_2228), .o(g66267_p) );
in01f04 g66267_u1 ( .a(g66267_p), .o(n_1359) );
no02s01 g66268_u0 ( .a(n_2214), .b(n_1808), .o(n_3223) );
na02f04 g66269_u0 ( .a(n_1357), .b(n_1966), .o(g66269_p) );
in01f02 g66269_u1 ( .a(g66269_p), .o(n_1358) );
na02f02 g66270_u0 ( .a(n_1355), .b(n_1228), .o(n_1356) );
na02s01 g66271_u0 ( .a(FE_OFN2214_n_15366), .b(n_1519), .o(n_2349) );
no02f08 g66272_u0 ( .a(n_844), .b(n_838), .o(n_1354) );
na03f02 TIMEBOOST_cell_24999 ( .a(n_10656), .b(FE_RN_221_0), .c(n_12772), .o(n_12951) );
no02f08 g66274_u0 ( .a(n_1467), .b(n_1034), .o(n_1799) );
no02f02 g66275_u0 ( .a(n_721), .b(n_611), .o(n_1162) );
no02f04 g66276_u0 ( .a(n_711), .b(n_609), .o(n_1161) );
na02f10 g66277_u0 ( .a(n_329), .b(n_1211), .o(n_2430) );
na02f02 g66278_u0 ( .a(n_16541), .b(n_15755), .o(g66278_p) );
in01f02 g66278_u1 ( .a(g66278_p), .o(n_2555) );
in01f08 g66281_u0 ( .a(n_3023), .o(n_3386) );
in01f10 g66282_u0 ( .a(n_2804), .o(n_3023) );
no02f20 g66285_u0 ( .a(n_1306), .b(n_16860), .o(n_2804) );
no02f01 g66286_u0 ( .a(n_1217), .b(n_840), .o(g66286_p) );
in01f02 g66286_u1 ( .a(g66286_p), .o(n_1541) );
na02f10 g66287_u0 ( .a(n_1248), .b(n_15922), .o(g66287_p) );
in01f10 g66287_u1 ( .a(g66287_p), .o(n_2777) );
no02f04 g66288_u0 ( .a(n_742), .b(n_871), .o(n_1352) );
no02f10 g66289_u0 ( .a(n_866), .b(n_960), .o(n_1351) );
na02f10 g66290_dup_u0 ( .a(n_15065), .b(n_2129), .o(g66290_dup_p) );
in01f10 g66290_dup_u1 ( .a(g66290_dup_p), .o(n_15445) );
no02f02 g66291_u0 ( .a(n_1448), .b(pci_target_unit_wbm_sm_pci_tar_read_request), .o(g66291_p) );
in01f02 g66291_u1 ( .a(g66291_p), .o(n_1798) );
in01f02 g66292_u0 ( .a(n_3004), .o(n_3504) );
in01f02 g66293_u0 ( .a(n_3248), .o(n_3004) );
no02f10 g66294_u0 ( .a(n_2553), .b(n_15291), .o(n_3248) );
no02f02 g66295_u0 ( .a(n_2042), .b(n_1754), .o(n_2347) );
no02f04 g66297_u0 ( .a(n_999), .b(n_959), .o(n_1350) );
na02s01 g66298_u0 ( .a(n_16964), .b(n_1347), .o(g66298_p) );
in01s01 g66298_u1 ( .a(g66298_p), .o(n_1349) );
no02f06 g66299_u0 ( .a(n_952), .b(n_587), .o(g66299_p) );
in01f04 g66299_u1 ( .a(g66299_p), .o(n_1346) );
no02f06 g66301_u0 ( .a(n_950), .b(n_855), .o(n_1433) );
no02f06 g66302_u0 ( .a(n_2127), .b(n_2126), .o(g66302_p) );
in01f06 g66302_u1 ( .a(g66302_p), .o(n_4806) );
no02f10 g66303_u0 ( .a(n_2553), .b(n_2552), .o(g66303_p) );
in01f10 g66303_u1 ( .a(g66303_p), .o(n_3018) );
no02f06 g66305_u0 ( .a(n_2126), .b(n_1777), .o(n_3368) );
no02f10 g66309_u0 ( .a(n_2552), .b(n_2453), .o(n_3295) );
no02f10 g66310_u0 ( .a(n_841), .b(n_843), .o(g66310_p) );
in01f08 g66310_u1 ( .a(g66310_p), .o(n_1345) );
na02s01 g66311_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q), .b(FE_OFN587_n_9692), .o(n_1540) );
no02f08 g66312_u0 ( .a(n_865), .b(n_744), .o(n_1344) );
no02f40 g66313_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_), .o(n_1539) );
no02f08 g66315_u0 ( .a(n_2344), .b(n_2685), .o(g66315_p) );
in01f08 g66315_u1 ( .a(g66315_p), .o(n_2345) );
no02f08 g66316_u0 ( .a(n_839), .b(n_743), .o(n_1343) );
no02f06 g66317_u0 ( .a(n_836), .b(n_747), .o(n_1342) );
no02m01 g66319_u0 ( .a(n_7622), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_2343) );
no02f06 g66320_u0 ( .a(n_627), .b(n_623), .o(n_1160) );
no02f08 g66321_u0 ( .a(n_837), .b(n_1007), .o(n_1341) );
no02f04 g66322_u0 ( .a(n_559), .b(wishbone_slave_unit_del_sync_comp_done_reg_main), .o(g66322_p) );
in01f02 g66322_u1 ( .a(g66322_p), .o(n_1696) );
na02f06 g66323_u0 ( .a(n_2125), .b(n_2795), .o(g66323_p) );
in01f04 g66323_u1 ( .a(g66323_p), .o(n_3221) );
no02f04 g66324_u0 ( .a(n_725), .b(n_621), .o(n_1159) );
no02f06 g66325_u0 ( .a(n_1004), .b(n_833), .o(n_1340) );
na02f10 g66327_u0 ( .a(n_2094), .b(n_16424), .o(g66327_p) );
in01f10 g66327_u1 ( .a(g66327_p), .o(n_3231) );
in01f08 g66328_u0 ( .a(n_2768), .o(n_7031) );
in01f08 g66332_u0 ( .a(n_3026), .o(n_2768) );
na02f08 g66336_u0 ( .a(n_2341), .b(n_16036), .o(g66336_p) );
in01f08 g66336_u1 ( .a(g66336_p), .o(n_3026) );
no02f08 g66337_u0 ( .a(n_700), .b(n_648), .o(n_1189) );
na02f01 g66338_u0 ( .a(n_15755), .b(n_16424), .o(g66338_p) );
in01f02 g66338_u1 ( .a(g66338_p), .o(n_2339) );
na02s01 g66339_u0 ( .a(n_2316), .b(FE_OFN2214_n_15366), .o(n_2767) );
na02m02 TIMEBOOST_cell_63995 ( .a(TIMEBOOST_net_20983), .b(FE_OFN1274_n_4096), .o(TIMEBOOST_net_15881) );
in01s01 TIMEBOOST_cell_45944 ( .a(TIMEBOOST_net_13904), .o(TIMEBOOST_net_13905) );
in01f08 g66346_u0 ( .a(n_1999), .o(n_3250) );
no02f10 g66347_u0 ( .a(n_1808), .b(n_1998), .o(n_1999) );
na02f01 g66348_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q), .b(FE_OFN1046_n_16657), .o(n_1795) );
na02m01 g66349_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q), .b(FE_OFN682_n_4460), .o(n_1537) );
ao12m02 g66350_u0 ( .a(n_2494), .b(n_716), .c(conf_wb_err_bc_in_846), .o(n_3001) );
ao12s01 g66352_u0 ( .a(configuration_set_pci_err_cs_bit8), .b(configuration_sync_pci_err_cs_8_delayed_del_bit), .c(configuration_sync_pci_err_cs_8_sync_del_bit), .o(n_1191) );
na02f20 g66353_u0 ( .a(pci_target_unit_pci_target_sm_read_completed_reg), .b(n_2337), .o(n_2883) );
ao12s01 g66354_u0 ( .a(n_2031), .b(n_1512), .c(n_15295), .o(n_2547) );
oa12f10 g66356_u0 ( .a(n_1507), .b(n_1220), .c(n_730), .o(n_2000) );
na02f02 g66357_u0 ( .a(n_16001), .b(n_16541), .o(g66357_p) );
in01f02 g66357_u1 ( .a(g66357_p), .o(n_3372) );
na02f06 g66358_u0 ( .a(n_1446), .b(n_15125), .o(g66358_p) );
in01f06 g66358_u1 ( .a(g66358_p), .o(TIMEBOOST_net_3) );
no02f02 g66359_u0 ( .a(n_930), .b(n_1334), .o(n_1469) );
na02f02 TIMEBOOST_cell_49248 ( .a(TIMEBOOST_net_14841), .b(g58406_db), .o(n_9001) );
ao22m04 g66361_u0 ( .a(n_713), .b(n_345), .c(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_), .d(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(n_1338) );
ao22s02 g66362_u0 ( .a(n_567), .b(n_362), .c(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_), .d(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .o(n_1337) );
ao22s01 g66363_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_956), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_649), .o(n_1794) );
ao22f04 g66365_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_969), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_662), .o(n_1793) );
ao22f02 g66366_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_946), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_639), .o(n_2121) );
na04f04 TIMEBOOST_cell_24587 ( .a(n_9901), .b(g57154_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q), .d(FE_OFN2189_n_8567), .o(n_11597) );
ao22f04 g66369_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_943), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_636), .o(n_2120) );
ao22f02 g66370_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_951), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_644), .o(n_2119) );
ao22f02 g66371_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_959), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_652), .o(n_2117) );
ao22f06 g66372_u0 ( .a(n_2115), .b(conf_wb_err_addr_in_963), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_656), .o(n_2116) );
ao22f02 g66373_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_971), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_664), .o(n_1790) );
ao22f08 g66374_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_957), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_650), .o(n_2114) );
ao22f02 g66375_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_961), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_654), .o(n_2113) );
ao22f01 g66376_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_953), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_646), .o(n_2111) );
ao22f02 g66377_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_944), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_637), .o(n_2110) );
na03f02 TIMEBOOST_cell_67088 ( .a(FE_OFN1596_n_13741), .b(n_13903), .c(TIMEBOOST_net_13805), .o(n_14277) );
ao22s01 g66379_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_966), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_659), .o(n_2108) );
ao22s01 g66381_u0 ( .a(n_1787), .b(conf_wb_err_addr_in_967), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_660), .o(n_2106) );
ao22s01 g66382_u0 ( .a(FE_OFN1617_n_1787), .b(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_665), .o(n_1789) );
ao22s01 g66383_u0 ( .a(n_2046), .b(pci_target_unit_pci_target_if_target_rd_completed), .c(pciu_pciif_bckp_stop_in), .d(output_backup_devsel_out_reg_Q), .o(n_2765) );
ao22f02 g66384_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_968), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_661), .o(n_2105) );
ao22f02 g66385_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_962), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_655), .o(n_2104) );
ao22s01 g66386_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_948), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_641), .o(n_1788) );
ao22f02 g66387_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_958), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_651), .o(n_1786) );
ao22s01 g66388_u0 ( .a(FE_OFN1620_n_1787), .b(conf_wb_err_addr_in_945), .c(FE_OFN1611_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_638), .o(n_1785) );
ao22f02 g66389_u0 ( .a(n_2115), .b(conf_wb_err_addr_in_947), .c(FE_OFN1612_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_640), .o(n_2103) );
ao22f04 g66390_u0 ( .a(n_2115), .b(conf_wb_err_addr_in_970), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_663), .o(n_2102) );
ao22f02 g66391_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_950), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_643), .o(n_1784) );
ao22f08 g66393_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_964), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_657), .o(n_1782) );
ao22f02 g66394_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_952), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_645), .o(n_2101) );
ao22f04 g66395_u0 ( .a(FE_OFN1621_n_1787), .b(conf_wb_err_addr_in_954), .c(FE_OFN1609_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_647), .o(n_2100) );
ao22f02 g66396_u0 ( .a(FE_OFN1617_n_1787), .b(conf_wb_err_addr_in_955), .c(FE_OFN1610_n_2122), .d(wishbone_slave_unit_pcim_sm_data_in_648), .o(n_1781) );
in01m02 g66397_u0 ( .a(FE_OFN2095_n_2520), .o(g66397_sb) );
na02m02 TIMEBOOST_cell_44244 ( .a(TIMEBOOST_net_13016), .b(g63601_sb), .o(n_7197) );
na02f01 TIMEBOOST_cell_70892 ( .a(TIMEBOOST_net_16740), .b(FE_OFN1184_n_3476), .o(TIMEBOOST_net_22654) );
na02f02 TIMEBOOST_cell_49898 ( .a(TIMEBOOST_net_15166), .b(g63088_sb), .o(n_5078) );
in01s04 g66398_u0 ( .a(FE_OFN795_n_2520), .o(g66398_sb) );
na03f02 TIMEBOOST_cell_73584 ( .a(TIMEBOOST_net_17463), .b(FE_OFN1196_n_4090), .c(g63006_sb), .o(n_5870) );
na02s01 g66398_u2 ( .a(parchk_pci_ad_reg_in_1209), .b(FE_OFN795_n_2520), .o(g66398_db) );
na03f02 TIMEBOOST_cell_73433 ( .a(TIMEBOOST_net_20538), .b(FE_OFN1258_n_4143), .c(g62485_sb), .o(n_6617) );
in01s01 g66399_u0 ( .a(n_2520), .o(g66399_sb) );
na03m02 TIMEBOOST_cell_70172 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q), .b(FE_OFN923_n_4740), .c(pci_target_unit_fifos_pciw_control_in_155), .o(TIMEBOOST_net_22294) );
na02m02 TIMEBOOST_cell_72071 ( .a(TIMEBOOST_net_23243), .b(TIMEBOOST_net_9781), .o(n_1598) );
na03f02 TIMEBOOST_cell_73650 ( .a(TIMEBOOST_net_17420), .b(FE_OFN1285_n_4097), .c(g62976_sb), .o(n_5930) );
na02s01 g66400_u2 ( .a(parchk_pci_ad_reg_in_1211), .b(FE_OFN795_n_2520), .o(g66400_db) );
na03m02 TIMEBOOST_cell_322 ( .a(n_1956), .b(g61735_sb), .c(g61735_db), .o(n_8349) );
in01s02 g66402_u0 ( .a(FE_OFN2096_n_2520), .o(g66402_sb) );
na02s01 g66402_u2 ( .a(parchk_pci_ad_reg_in_1227), .b(FE_OFN2096_n_2520), .o(g66402_db) );
na04s08 TIMEBOOST_cell_64962 ( .a(n_3752), .b(g64805_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q), .d(FE_OFN649_n_4497), .o(n_3754) );
in01s04 g66403_u0 ( .a(FE_OFN2096_n_2520), .o(g66403_sb) );
na03m10 TIMEBOOST_cell_70270 ( .a(FE_OFN262_n_9851), .b(FE_OFN1666_n_9477), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q), .o(TIMEBOOST_net_22343) );
na02s01 g66403_u2 ( .a(parchk_pci_ad_reg_in_1220), .b(FE_OFN2096_n_2520), .o(g66403_db) );
na02s01 g66404_u2 ( .a(FE_OFN1780_parchk_pci_ad_reg_in_1221), .b(FE_OFN2096_n_2520), .o(g66404_db) );
na02f01 TIMEBOOST_cell_63361 ( .a(TIMEBOOST_net_20627), .b(FE_OFN1131_g64577_p), .o(TIMEBOOST_net_15138) );
na02m02 TIMEBOOST_cell_69055 ( .a(TIMEBOOST_net_21735), .b(TIMEBOOST_net_16240), .o(TIMEBOOST_net_17021) );
na02s01 g66405_u2 ( .a(parchk_pci_ad_reg_in_1217), .b(FE_OFN2096_n_2520), .o(g66405_db) );
na03s02 TIMEBOOST_cell_330 ( .a(n_1944), .b(g61764_sb), .c(g61764_db), .o(n_8283) );
in01s01 g66406_u0 ( .a(FE_OFN2095_n_2520), .o(g66406_sb) );
na02s01 g66406_u2 ( .a(parchk_pci_ad_reg_in_1230), .b(FE_OFN2095_n_2520), .o(g66406_db) );
na03f02 TIMEBOOST_cell_33493 ( .a(TIMEBOOST_net_8790), .b(FE_OFN1168_n_5592), .c(g62097_sb), .o(n_5607) );
na02s01 g66407_u2 ( .a(FE_OFN2096_n_2520), .b(parchk_pci_ad_reg_in_1225), .o(g66407_db) );
na02m06 TIMEBOOST_cell_72092 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q), .b(pci_target_unit_fifos_pciw_addr_data_in_144), .o(TIMEBOOST_net_23254) );
na02f01 TIMEBOOST_cell_71810 ( .a(TIMEBOOST_net_13707), .b(FE_OFN1774_n_13800), .o(TIMEBOOST_net_23113) );
na02s01 g66408_u2 ( .a(FE_OFN1778_parchk_pci_ad_reg_in_1222), .b(FE_OFN2096_n_2520), .o(g66408_db) );
na03f02 TIMEBOOST_cell_73743 ( .a(TIMEBOOST_net_13678), .b(FE_OFN1757_n_12681), .c(FE_OCPN1866_n_12377), .o(n_12742) );
na02s01 g66409_u2 ( .a(parchk_pci_ad_reg_in_1223), .b(FE_OFN2096_n_2520), .o(g66409_db) );
na02s01 TIMEBOOST_cell_63126 ( .a(FE_OFN1789_n_9823), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q), .o(TIMEBOOST_net_20510) );
na02f02 TIMEBOOST_cell_53546 ( .a(TIMEBOOST_net_16990), .b(g62775_sb), .o(n_5444) );
na02s01 g66410_u2 ( .a(parchk_pci_ad_reg_in_1208), .b(FE_OFN795_n_2520), .o(g66410_db) );
na03f02 TIMEBOOST_cell_66423 ( .a(TIMEBOOST_net_17544), .b(FE_OFN1320_n_6436), .c(g62618_sb), .o(n_7374) );
na02s01 g66411_u2 ( .a(n_2648), .b(n_2520), .o(g66411_db) );
na04f10 TIMEBOOST_cell_72405 ( .a(FE_RN_633_0), .b(n_15598), .c(n_360), .d(FE_RN_632_0), .o(FE_RN_636_0) );
na02s01 g66412_u2 ( .a(parchk_pci_ad_reg_in_1229), .b(n_2520), .o(g66412_db) );
na02s01 TIMEBOOST_cell_47966 ( .a(TIMEBOOST_net_14200), .b(FE_OFN950_n_2055), .o(TIMEBOOST_net_12493) );
na02m01 TIMEBOOST_cell_68185 ( .a(TIMEBOOST_net_21300), .b(FE_OFN937_n_2292), .o(TIMEBOOST_net_14091) );
na02s01 g66413_u2 ( .a(n_8511), .b(n_2520), .o(g66413_db) );
no03f04 TIMEBOOST_cell_66104 ( .a(FE_RN_396_0), .b(FE_OFN1707_n_4868), .c(FE_RN_124_0), .o(TIMEBOOST_net_771) );
na02s01 g66414_u2 ( .a(n_2520), .b(parchk_pci_ad_reg_in_1214), .o(g66414_db) );
na02m04 TIMEBOOST_cell_68578 ( .a(g64915_sb), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q), .o(TIMEBOOST_net_21497) );
in01s01 g66415_u0 ( .a(FE_OFN795_n_2520), .o(g66415_sb) );
na02s01 g66415_u2 ( .a(parchk_pci_ad_reg_in_1232), .b(FE_OFN795_n_2520), .o(g66415_db) );
na02s01 TIMEBOOST_cell_48725 ( .a(pci_target_unit_fifos_pciw_addr_data_in_132), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q), .o(TIMEBOOST_net_14580) );
na02s01 g66416_u2 ( .a(FE_OFN2095_n_2520), .b(parchk_pci_ad_reg_in_1215), .o(g66416_db) );
na02s04 TIMEBOOST_cell_63318 ( .a(FE_OFN264_n_9849), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q), .o(TIMEBOOST_net_20606) );
na02s01 g66417_u2 ( .a(parchk_pci_ad_reg_in_1206), .b(n_2520), .o(g66417_db) );
na02m10 TIMEBOOST_cell_42965 ( .a(pci_target_unit_fifos_pciw_addr_data_in_134), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q), .o(TIMEBOOST_net_12377) );
na02s01 g66418_u2 ( .a(parchk_pci_ad_reg_in_1226), .b(FE_OFN2095_n_2520), .o(g66418_db) );
na04f02 TIMEBOOST_cell_67939 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q), .b(FE_OFN1129_g64577_p), .c(n_4033), .d(g62851_sb), .o(n_5267) );
in01s01 TIMEBOOST_cell_45897 ( .a(TIMEBOOST_net_13963), .o(TIMEBOOST_net_13858) );
na02s01 g66419_u2 ( .a(parchk_pci_ad_reg_in_1210), .b(n_2520), .o(g66419_db) );
na03f08 TIMEBOOST_cell_21828 ( .a(FE_RN_360_0), .b(n_16474), .c(FE_RN_535_0), .o(n_16268) );
na02f01 TIMEBOOST_cell_18305 ( .a(configuration_pci_err_addr_481), .b(FE_OFN1185_n_3476), .o(TIMEBOOST_net_5516) );
na02s01 g66420_u2 ( .a(n_2509), .b(FE_OFN795_n_2520), .o(g66420_db) );
na02m06 TIMEBOOST_cell_52257 ( .a(g64337_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q), .o(TIMEBOOST_net_16346) );
na03f02 TIMEBOOST_cell_34827 ( .a(TIMEBOOST_net_9337), .b(FE_OFN1412_n_8567), .c(g57592_sb), .o(n_10286) );
na02s01 g66421_u2 ( .a(parchk_pci_ad_reg_in_1212), .b(FE_OFN795_n_2520), .o(g66421_db) );
na03f02 TIMEBOOST_cell_34829 ( .a(TIMEBOOST_net_9369), .b(FE_OFN1412_n_8567), .c(g57257_sb), .o(n_11496) );
na02f02 TIMEBOOST_cell_49828 ( .a(TIMEBOOST_net_15131), .b(g63175_sb), .o(n_4949) );
na02s01 g66422_u2 ( .a(parchk_pci_ad_reg_in_1233), .b(FE_OFN795_n_2520), .o(g66422_db) );
in01s01 TIMEBOOST_cell_67741 ( .a(pci_target_unit_fifos_pcir_data_in_164), .o(TIMEBOOST_net_21168) );
na02s01 TIMEBOOST_cell_45789 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q), .o(TIMEBOOST_net_13789) );
na02m02 TIMEBOOST_cell_69091 ( .a(TIMEBOOST_net_21753), .b(g65399_sb), .o(TIMEBOOST_net_12551) );
na03f02 TIMEBOOST_cell_34793 ( .a(TIMEBOOST_net_9557), .b(FE_OFN1381_n_8567), .c(g57425_sb), .o(n_10361) );
na02s01 g66424_u2 ( .a(parchk_pci_ad_reg_in_1228), .b(FE_OFN795_n_2520), .o(g66424_db) );
no03m08 TIMEBOOST_cell_67111 ( .a(n_16003), .b(n_15924), .c(n_16287), .o(TIMEBOOST_net_94) );
in01s01 TIMEBOOST_cell_45898 ( .a(TIMEBOOST_net_13858), .o(TIMEBOOST_net_13859) );
na02s01 g66425_u2 ( .a(n_2651), .b(n_2520), .o(g66425_db) );
in01s01 TIMEBOOST_cell_45899 ( .a(TIMEBOOST_net_13860), .o(wbs_dat_i_23_) );
na02s01 g66426_u2 ( .a(parchk_pci_ad_reg_in_1207), .b(n_2520), .o(g66426_db) );
in01s01 TIMEBOOST_cell_45900 ( .a(TIMEBOOST_net_13861), .o(TIMEBOOST_net_13860) );
na02s01 g66427_u2 ( .a(n_3030), .b(n_2520), .o(g66427_db) );
na02m01 TIMEBOOST_cell_52811 ( .a(n_3780), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q), .o(TIMEBOOST_net_16623) );
na02s01 g66428_u2 ( .a(parchk_pci_ad_reg_in_1219), .b(FE_OFN2096_n_2520), .o(g66428_db) );
na02s01 g66429_u2 ( .a(parchk_pci_ad_reg_in_1235), .b(FE_OFN795_n_2520), .o(g66429_db) );
na02f01 TIMEBOOST_cell_51623 ( .a(FE_OFN1736_n_16317), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q), .o(TIMEBOOST_net_16029) );
na04f04 TIMEBOOST_cell_73277 ( .a(configuration_wb_err_data_595), .b(FE_OFN1168_n_5592), .c(TIMEBOOST_net_13847), .d(g62096_sb), .o(n_5608) );
na02s01 g66430_u2 ( .a(parchk_pci_ad_reg_in_1218), .b(FE_OFN2095_n_2520), .o(g66430_db) );
in01s10 g66433_u0 ( .a(pci_target_unit_del_sync_req_done_reg), .o(g66433_sb) );
na03f02 TIMEBOOST_cell_66544 ( .a(TIMEBOOST_net_16792), .b(FE_OFN1331_n_13547), .c(g53906_sb), .o(n_13535) );
na02s01 g66433_u2 ( .a(pci_target_unit_del_sync_req_comp_pending), .b(pci_target_unit_del_sync_req_done_reg), .o(g66433_db) );
na02s02 TIMEBOOST_cell_51855 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q), .b(g65852_sb), .o(TIMEBOOST_net_16145) );
oa12s01 g66454_u0 ( .a(n_944), .b(n_1334), .c(n_1263), .o(n_1335) );
in01m02 g66456_u0 ( .a(n_325), .o(g66456_sb) );
na02m02 g66456_u3 ( .a(g66456_da), .b(g66456_db), .o(n_1532) );
na02m01 g66456_u2 ( .a(wishbone_slave_unit_del_sync_req_comp_pending), .b(n_325), .o(g66456_db) );
na02m02 g66456_u1 ( .a(wishbone_slave_unit_del_sync_sync_req_comp_pending), .b(g66456_sb), .o(g66456_da) );
in01m08 g66457_u0 ( .a(pci_target_unit_pci_target_sm_n_3), .o(g66457_sb) );
na02f02 TIMEBOOST_cell_45189 ( .a(n_14740), .b(n_14839), .o(TIMEBOOST_net_13489) );
na03m02 TIMEBOOST_cell_72414 ( .a(TIMEBOOST_net_23122), .b(TIMEBOOST_net_17193), .c(g61943_sb), .o(TIMEBOOST_net_16954) );
na03m01 TIMEBOOST_cell_72448 ( .a(TIMEBOOST_net_10206), .b(n_4730), .c(g60688_sb), .o(n_3872) );
no02m04 g66458_u0 ( .a(wbm_adr_o_3_), .b(wbm_adr_o_2_), .o(g66458_p0) );
ao12m02 g66458_u1 ( .a(g66458_p0), .b(wbm_adr_o_2_), .c(wbm_adr_o_3_), .o(n_740) );
na02f80 g66458_u2 ( .a(wbm_adr_o_2_), .b(wbm_adr_o_3_), .o(g66458_p) );
in01f40 g66458_u3 ( .a(g66458_p), .o(n_1674) );
no02s01 g66459_u0 ( .a(wbu_addr_in_252), .b(wbu_addr_in_251), .o(g66459_p0) );
ao12s01 g66459_u1 ( .a(g66459_p0), .b(wbu_addr_in_252), .c(wbu_addr_in_251), .o(n_739) );
in01s01 g66462_u0 ( .a(n_16030), .o(n_1133) );
no02s01 g66464_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(g66464_p0) );
ao12s01 g66464_u1 ( .a(g66464_p0), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_1225) );
na02s01 g66464_u2 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q), .o(g66464_p) );
in01s01 g66464_u3 ( .a(g66464_p), .o(n_1224) );
no02s01 g66465_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .o(g66465_p0) );
ao12s01 g66465_u1 ( .a(g66465_p0), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .o(n_741) );
na02f01 g66465_u2 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_), .o(g66465_p) );
in01f02 g66465_u3 ( .a(g66465_p), .o(n_1418) );
in01f40 g66467_u0 ( .a(n_568), .o(n_1413) );
in01f10 g66470_u0 ( .a(n_1011), .o(n_1175) );
in01s01 g66471_u0 ( .a(n_947), .o(n_566) );
in01s01 g66472_u0 ( .a(n_948), .o(n_733) );
no02f10 g66473_u0 ( .a(n_1332), .b(n_540), .o(g66473_p) );
ao12f08 g66473_u1 ( .a(g66473_p), .b(n_1332), .c(n_540), .o(n_1333) );
no02f10 g66475_u0 ( .a(n_1330), .b(n_558), .o(g66475_p) );
ao12f08 g66475_u1 ( .a(g66475_p), .b(n_1330), .c(n_558), .o(n_1331) );
ao22m01 g66476_u0 ( .a(n_76), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_), .d(n_816), .o(n_1329) );
na03m06 TIMEBOOST_cell_69192 ( .a(pci_target_unit_fifos_pciw_cbe_in_154), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q), .c(FE_OFN929_n_4730), .o(TIMEBOOST_net_21804) );
na02s01 TIMEBOOST_cell_52665 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q), .o(TIMEBOOST_net_16550) );
na04f02 TIMEBOOST_cell_35118 ( .a(wbs_dat_o_24_), .b(g52519_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_123), .d(FE_OFN1471_g52675_p), .o(n_13740) );
in01s01 g66479_u0 ( .a(wishbone_slave_unit_pci_initiator_if_write_req_int), .o(n_1780) );
in01s01 g66483_u0 ( .a(wishbone_slave_unit_del_sync_req_rty_exp_reg), .o(n_1327) );
in01s01 g66497_u0 ( .a(pci_target_unit_del_sync_req_rty_exp_reg), .o(n_249) );
in01s01 g66536_u0 ( .a(pci_target_unit_del_sync_comp_done_reg_main), .o(n_2146) );
in01f01 g66542_u0 ( .a(n_1325), .o(n_1326) );
no02f08 g66543_u0 ( .a(n_943), .b(n_288), .o(n_1325) );
na02f08 g66544_u0 ( .a(n_1107), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(g66544_p) );
in01f04 g66544_u1 ( .a(g66544_p), .o(n_908) );
no02f01 g66547_u0 ( .a(n_914), .b(n_1174), .o(g66547_p) );
in01f02 g66547_u1 ( .a(g66547_p), .o(n_1699) );
no02f02 g66548_u0 ( .a(n_1468), .b(output_backup_trdy_out_reg_Q), .o(n_1126) );
no02f40 g66549_u0 ( .a(n_412), .b(wishbone_slave_unit_wishbone_slave_img_hit_2_), .o(n_931) );
na02s01 g66550_u0 ( .a(n_1173), .b(wishbone_slave_unit_fifos_wbw_whole_waddr), .o(g66550_p) );
in01m01 g66550_u1 ( .a(g66550_p), .o(n_905) );
in01f02 g66551_u0 ( .a(n_1779), .o(n_7622) );
in01f04 g66552_u0 ( .a(n_15055), .o(n_1779) );
na02f02 g66554_u0 ( .a(n_929), .b(n_1263), .o(n_930) );
no02s01 g66555_u0 ( .a(n_2483), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(n_2999) );
no02f80 g66556_u0 ( .a(n_560), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_), .o(n_1715) );
no02s03 g66577_u0 ( .a(n_748), .b(wbs_adr_i_4_), .o(g66577_p) );
in01s02 g66577_u1 ( .a(g66577_p), .o(n_1666) );
na02f10 g66579_u0 ( .a(n_1317), .b(n_1293), .o(n_4736) );
no02f08 g66580_u0 ( .a(n_1334), .b(n_221), .o(n_1437) );
in01f02 g66581_u0 ( .a(n_1124), .o(n_1125) );
na02f08 g66582_u0 ( .a(n_937), .b(pci_target_unit_del_sync_comp_cycle_count_7_), .o(n_1124) );
na02f40 g66583_u0 ( .a(n_1294), .b(n_1316), .o(g66583_p) );
in01f20 g66583_u1 ( .a(g66583_p), .o(n_4727) );
na02f01 g66584_u0 ( .a(n_1318), .b(n_1174), .o(g66584_p) );
in01f04 g66584_u1 ( .a(g66584_p), .o(n_2299) );
in01m06 g66585_u0 ( .a(n_1122), .o(n_1123) );
na02m10 g66586_u0 ( .a(n_928), .b(wishbone_slave_unit_del_sync_comp_cycle_count_7_), .o(n_1122) );
in01f08 g66590_u0 ( .a(n_1808), .o(n_4874) );
na02f10 g66591_u0 ( .a(n_993), .b(n_1104), .o(n_1808) );
no02m08 g66592_u0 ( .a(n_915), .b(n_924), .o(n_2872) );
no02f10 g66593_u0 ( .a(n_900), .b(n_921), .o(n_1229) );
no02f02 g66594_u0 ( .a(n_927), .b(n_909), .o(n_1381) );
no02m10 g66595_u0 ( .a(n_901), .b(n_926), .o(n_2756) );
na02s01 g66596_u0 ( .a(configuration_sync_isr_2_delayed_del_bit), .b(configuration_sync_isr_2_sync_del_bit), .o(n_925) );
no02f20 g66597_u0 ( .a(n_877), .b(n_902), .o(n_1480) );
no02f02 g66598_u0 ( .a(n_16291), .b(n_16544), .o(n_2560) );
no02f80 g66599_u0 ( .a(wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_Q), .b(wishbone_slave_unit_del_sync_comp_flush_out), .o(n_9941) );
in01f04 g66600_u0 ( .a(n_2553), .o(n_2331) );
in01f10 g66602_u0 ( .a(n_2094), .o(n_2553) );
in01f10 g66603_u0 ( .a(n_1777), .o(n_2094) );
na02f20 g66604_u0 ( .a(n_15275), .b(n_15231), .o(n_1777) );
no02f10 g66605_u0 ( .a(n_904), .b(n_895), .o(n_2428) );
na02m10 g66607_u0 ( .a(n_257), .b(n_432), .o(g66607_p) );
in01m06 g66607_u1 ( .a(g66607_p), .o(n_1624) );
na02m01 g66608_u0 ( .a(n_15365), .b(parity_checker_frame_dec2), .o(n_3020) );
no02f20 g66612_u0 ( .a(n_924), .b(n_518), .o(n_2929) );
no02s01 g66613_u0 ( .a(n_2597), .b(n_1774), .o(n_2599) );
no02s01 g66614_u0 ( .a(n_1084), .b(configuration_isr_bit_2975), .o(n_1120) );
no02f20 g66615_u0 ( .a(n_923), .b(n_917), .o(n_2411) );
no02s01 g66616_u0 ( .a(n_976), .b(pci_target_unit_pci_target_sm_n_3), .o(n_922) );
no02f10 g66617_u0 ( .a(n_911), .b(n_921), .o(n_2235) );
no02f10 g66620_u0 ( .a(n_1005), .b(n_1009), .o(g66620_p) );
in01f10 g66620_u1 ( .a(g66620_p), .o(n_4501) );
no02m01 g66621_u0 ( .a(n_16867), .b(n_15680), .o(n_1322) );
no02f10 g66627_u0 ( .a(n_538), .b(n_1005), .o(g66627_p) );
in01f10 g66627_u1 ( .a(g66627_p), .o(n_4490) );
na02f01 g66628_u0 ( .a(n_1118), .b(n_1174), .o(g66628_p) );
in01f02 g66628_u1 ( .a(g66628_p), .o(n_2053) );
in01m01 g66630_u0 ( .a(n_1269), .o(n_1119) );
no02f20 g66631_u0 ( .a(n_886), .b(n_891), .o(n_1269) );
no02m40 g66632_u0 ( .a(n_919), .b(n_920), .o(n_2305) );
no02f20 g66633_u0 ( .a(n_894), .b(n_918), .o(n_1390) );
no02f08 g66634_u0 ( .a(n_927), .b(n_956), .o(n_2237) );
no02f20 g66636_u0 ( .a(n_910), .b(n_941), .o(n_2426) );
no02f08 g66637_u0 ( .a(n_917), .b(n_916), .o(n_1968) );
na02f01 g66638_u0 ( .a(n_1318), .b(n_1117), .o(n_2292) );
in01f01 g66639_u0 ( .a(n_1523), .o(n_1524) );
no02f06 g66640_u0 ( .a(n_790), .b(wishbone_slave_unit_wishbone_slave_c_state), .o(n_1523) );
no02f01 g66641_u0 ( .a(n_888), .b(n_939), .o(n_940) );
na02f01 g66642_u0 ( .a(n_1118), .b(n_1117), .o(n_2047) );
na04f04 TIMEBOOST_cell_24220 ( .a(n_9529), .b(g57409_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q), .d(FE_OFN1419_n_8567), .o(n_11334) );
no02f20 g66644_u0 ( .a(n_916), .b(n_915), .o(n_1227) );
no02f04 g66645_u0 ( .a(n_914), .b(n_1117), .o(n_2248) );
na02f20 g66646_u0 ( .a(n_913), .b(n_912), .o(g66646_p) );
in01f10 g66646_u1 ( .a(g66646_p), .o(n_1481) );
no02f20 g66647_u0 ( .a(n_911), .b(n_910), .o(n_1228) );
no02f10 g66648_u0 ( .a(n_563), .b(n_977), .o(n_1116) );
na02f02 g66649_u0 ( .a(n_1188), .b(n_1115), .o(g66649_p) );
in01f04 g66649_u1 ( .a(g66649_p), .o(n_9528) );
na02f40 g66650_u0 ( .a(n_1317), .b(n_1316), .o(g66650_p) );
in01f20 g66650_u1 ( .a(g66650_p), .o(n_4725) );
no02f10 g66651_u0 ( .a(n_892), .b(n_909), .o(n_2427) );
na02f02 g66652_u0 ( .a(n_1290), .b(n_1115), .o(g66652_p) );
in01f04 g66652_u1 ( .a(g66652_p), .o(n_9502) );
na02f08 g66653_u0 ( .a(n_1288), .b(n_1315), .o(n_9697) );
in01s01 g66655_u0 ( .a(FE_OCPN1875_n_14526), .o(n_1522) );
na02f20 g66658_u0 ( .a(n_1509), .b(n_1210), .o(g66658_p) );
in01f20 g66658_u1 ( .a(g66658_p), .o(n_4669) );
in01f04 g66660_u0 ( .a(n_2127), .o(n_2341) );
na02f08 g66661_u0 ( .a(n_15275), .b(n_15756), .o(n_2127) );
na02m01 g66662_u0 ( .a(n_2763), .b(n_653), .o(g66662_p) );
in01m02 g66662_u1 ( .a(g66662_p), .o(n_2764) );
no02f08 g66663_u0 ( .a(n_16033), .b(n_1291), .o(g66663_p) );
in01f06 g66663_u1 ( .a(g66663_p), .o(n_2126) );
no02f08 g66664_u0 ( .a(n_885), .b(n_881), .o(n_1270) );
in01f10 g66667_u0 ( .a(n_16151), .o(n_2215) );
no02f40 g66669_u0 ( .a(n_1316), .b(n_980), .o(g66669_p) );
in01f20 g66669_u1 ( .a(g66669_p), .o(n_16657) );
no02m04 g66670_u0 ( .a(n_1334), .b(n_906), .o(n_907) );
no02f02 g66671_u0 ( .a(n_946), .b(n_884), .o(n_2306) );
no02f40 g66672_u0 ( .a(n_1316), .b(n_813), .o(g66672_p) );
in01f40 g66672_u1 ( .a(g66672_p), .o(n_4740) );
in01f20 g66701_u0 ( .a(FE_OFN2214_n_15366), .o(n_2301) );
na02f10 g66710_u0 ( .a(n_1289), .b(n_1315), .o(n_9690) );
na02f02 g66711_u0 ( .a(n_1115), .b(n_1315), .o(n_9902) );
no02f20 g66712_u0 ( .a(n_904), .b(n_903), .o(n_1409) );
no02f02 g66713_u0 ( .a(n_902), .b(n_889), .o(n_2681) );
na02f20 g66714_u0 ( .a(n_1198), .b(n_1519), .o(g66714_p) );
in01f20 g66714_u1 ( .a(g66714_p), .o(n_2795) );
no02m20 g66715_u0 ( .a(n_901), .b(n_900), .o(n_2433) );
no02f20 g66716_u0 ( .a(n_899), .b(n_896), .o(n_1373) );
na02s01 g66717_u0 ( .a(n_1334), .b(n_1263), .o(n_944) );
na02f80 g66724_u0 ( .a(n_898), .b(wbm_ack_i), .o(n_1998) );
na02f10 g66726_u0 ( .a(n_791), .b(pci_target_unit_pci_target_sm_master_will_request_read), .o(g66726_p) );
in01f08 g66726_u1 ( .a(g66726_p), .o(n_1824) );
na02f20 g66727_u0 ( .a(n_16867), .b(n_15680), .o(n_1306) );
na02f40 g66728_u0 ( .a(n_1113), .b(n_1107), .o(g66728_p) );
in01f40 g66728_u1 ( .a(g66728_p), .o(n_4655) );
in01m08 g66732_u0 ( .a(n_1435), .o(n_9175) );
na03f80 g66733_u0 ( .a(n_61), .b(pci_target_unit_pci_target_sm_n_2), .c(n_278), .o(n_1435) );
in01s01 g66734_u0 ( .a(n_1304), .o(n_9178) );
na02s01 g66735_u0 ( .a(n_520), .b(n_1628), .o(n_1304) );
no02f40 g66736_u0 ( .a(n_897), .b(n_896), .o(n_2463) );
na02f04 g66737_u0 ( .a(n_2609), .b(n_2742), .o(g66737_p) );
in01f04 g66737_u1 ( .a(g66737_p), .o(n_3222) );
na02f20 g66738_u0 ( .a(n_534), .b(n_912), .o(g66738_p) );
in01f10 g66738_u1 ( .a(g66738_p), .o(n_2982) );
na02s01 g66739_u0 ( .a(FE_OFN1612_n_2122), .b(n_1111), .o(n_1112) );
na02f08 g66742_u0 ( .a(n_1173), .b(n_1288), .o(g66742_p) );
in01f10 g66742_u1 ( .a(g66742_p), .o(n_9428) );
no02f40 g66743_u0 ( .a(n_1197), .b(n_1519), .o(n_1813) );
no02f04 g66744_u0 ( .a(n_946), .b(n_945), .o(n_1282) );
oa12f08 g66745_u0 ( .a(n_1109), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .c(n_8953), .o(n_1110) );
na02s01 g66746_u0 ( .a(FE_OFN1612_n_2122), .b(wishbone_slave_unit_pcim_sm_be_in_558), .o(n_1108) );
no02f20 g66749_u0 ( .a(n_890), .b(n_895), .o(n_3007) );
in01s01 g66751_u0 ( .a(n_6943), .o(n_2134) );
na02f40 g66752_u0 ( .a(n_1432), .b(wishbone_slave_unit_wishbone_slave_c_state_2), .o(g66752_p) );
in01f40 g66752_u1 ( .a(g66752_p), .o(n_6943) );
na02f20 g66753_u0 ( .a(n_1107), .b(n_1195), .o(g66753_p) );
in01f20 g66753_u1 ( .a(g66753_p), .o(n_4671) );
no02f02 g66754_u0 ( .a(n_957), .b(n_956), .o(n_3194) );
no02f08 g66755_u0 ( .a(n_894), .b(n_893), .o(n_1478) );
na02f10 g66756_u0 ( .a(n_1188), .b(n_1440), .o(n_9692) );
no02m08 g66757_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .b(n_1014), .o(n_1299) );
na02f20 g66758_u0 ( .a(n_1195), .b(n_1194), .o(n_4392) );
na02f10 g66759_u0 ( .a(n_1017), .b(n_1316), .o(g66759_p) );
in01f10 g66759_u1 ( .a(g66759_p), .o(n_4730) );
no02f01 g66760_u0 ( .a(n_892), .b(n_512), .o(n_3192) );
na02f20 g66761_u0 ( .a(n_1106), .b(n_1107), .o(n_4409) );
in01f04 g66765_u0 ( .a(n_1514), .o(n_1515) );
no02f02 g66768_u0 ( .a(n_945), .b(n_887), .o(n_2755) );
na02s01 g66769_u0 ( .a(FE_OFN1612_n_2122), .b(wishbone_slave_unit_pcim_sm_be_in_557), .o(n_1105) );
na02f01 g66770_u0 ( .a(n_1290), .b(n_1440), .o(n_9694) );
na02f04 g66771_u0 ( .a(n_16307), .b(n_1774), .o(n_1513) );
no02f20 g66772_u0 ( .a(n_891), .b(n_890), .o(n_2228) );
na02f10 g66773_u0 ( .a(n_1210), .b(n_1201), .o(g66773_p) );
in01f20 g66773_u1 ( .a(g66773_p), .o(n_4677) );
no02f02 g66774_u0 ( .a(n_941), .b(n_549), .o(n_1355) );
no02f10 g66775_u0 ( .a(n_992), .b(n_1104), .o(n_3310) );
na02f01 g66776_u0 ( .a(n_1103), .b(n_1117), .o(n_2055) );
na02f08 g66777_u0 ( .a(n_1173), .b(n_1289), .o(g66777_p) );
in01f10 g66777_u1 ( .a(g66777_p), .o(n_9477) );
no02f08 g66778_u0 ( .a(n_874), .b(n_893), .o(n_964) );
no02f04 g66779_u0 ( .a(n_1739), .b(n_2078), .o(n_2329) );
na02f08 g66780_u0 ( .a(n_1294), .b(n_1293), .o(n_4734) );
no02f04 g66781_u0 ( .a(n_889), .b(n_888), .o(n_2705) );
in01f20 g66783_u0 ( .a(n_1366), .o(n_1196) );
na02f40 g66784_u0 ( .a(n_976), .b(pci_target_unit_pci_target_sm_n_3), .o(n_1366) );
na02m06 g66785_u0 ( .a(n_1440), .b(n_1315), .o(n_9687) );
no02f10 g66786_u0 ( .a(n_903), .b(n_530), .o(n_965) );
no02f20 g66787_u0 ( .a(n_746), .b(n_745), .o(n_2475) );
na02m20 g66788_u0 ( .a(n_1194), .b(n_1210), .o(n_4497) );
na02f01 g66789_u0 ( .a(n_1103), .b(n_1174), .o(g66789_p) );
in01f02 g66789_u1 ( .a(g66789_p), .o(n_2037) );
in01s04 g66794_u0 ( .a(n_1445), .o(n_2214) );
na02s01 g66796_u0 ( .a(FE_OFN1612_n_2122), .b(wishbone_slave_unit_pcim_sm_be_in_559), .o(n_1202) );
in01s01 g66797_u0 ( .a(n_1758), .o(n_1759) );
no02f01 g66798_u0 ( .a(n_1512), .b(n_1505), .o(n_1758) );
no02f40 g66799_u0 ( .a(n_899), .b(n_923), .o(n_2596) );
no02s01 g66800_u0 ( .a(n_2031), .b(output_backup_trdy_out_reg_Q), .o(n_2280) );
no02s01 g66801_u0 ( .a(n_2031), .b(n_15302), .o(n_2729) );
no02f20 g66802_u0 ( .a(n_533), .b(n_745), .o(n_2914) );
no02f02 g66803_u0 ( .a(n_887), .b(n_957), .o(n_2431) );
na02f40 g66805_u0 ( .a(n_812), .b(n_1316), .o(g66805_p) );
in01f20 g66805_u1 ( .a(g66805_p), .o(n_4732) );
in01f01 g66807_u0 ( .a(n_15065), .o(n_2449) );
in01f01 g66811_u0 ( .a(n_1447), .o(n_1448) );
no02f06 g66812_u0 ( .a(n_1200), .b(n_681), .o(n_1447) );
na02f10 g66813_u0 ( .a(n_1210), .b(n_1107), .o(g66813_p) );
in01f08 g66813_u1 ( .a(g66813_p), .o(n_4508) );
na02f10 g66814_u0 ( .a(n_1440), .b(n_1173), .o(n_9904) );
in01f01 g66820_u0 ( .a(n_15370), .o(n_1684) );
na02f40 g66822_u0 ( .a(n_1194), .b(n_1113), .o(n_4460) );
no02f06 g66823_u0 ( .a(n_16291), .b(FE_OCPN1868_n_16289), .o(n_1446) );
na04m04 TIMEBOOST_cell_73114 ( .a(TIMEBOOST_net_8272), .b(g65797_db), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q), .d(FE_OFN701_n_7845), .o(TIMEBOOST_net_14828) );
no02f02 g66825_u0 ( .a(wishbone_slave_unit_fifos_wbr_control_in), .b(n_2685), .o(g66825_p) );
in01f02 g66825_u1 ( .a(g66825_p), .o(n_3480) );
no02f40 g66826_u0 ( .a(n_977), .b(n_897), .o(n_1374) );
na02s01 g66827_u0 ( .a(n_1347), .b(n_16816), .o(g66827_p) );
in01s01 g66827_u1 ( .a(g66827_p), .o(n_1101) );
na02f20 g66829_u0 ( .a(n_1106), .b(n_1201), .o(n_4454) );
na02s01 g66830_u0 ( .a(n_1774), .b(n_5755), .o(n_1100) );
no02f40 g66831_u0 ( .a(n_886), .b(n_885), .o(n_2435) );
no02f10 g66832_u0 ( .a(n_920), .b(n_926), .o(n_1241) );
in01f10 g66852_u0 ( .a(n_2494), .o(n_2493) );
in01m06 g66853_u0 ( .a(n_2344), .o(n_2494) );
na02f40 g66854_u0 ( .a(n_1459), .b(wishbone_slave_unit_pci_initiator_sm_mabort1), .o(g66854_p) );
in01f20 g66854_u1 ( .a(g66854_p), .o(n_2344) );
no02f20 g66855_u0 ( .a(n_1221), .b(n_2742), .o(n_2028) );
na02f02 g66856_u0 ( .a(n_1173), .b(n_1115), .o(g66856_p) );
in01f04 g66856_u1 ( .a(g66856_p), .o(n_9531) );
no02f40 g66857_u0 ( .a(n_746), .b(n_528), .o(n_1442) );
na02f01 g66858_u0 ( .a(FE_OFN1612_n_2122), .b(wishbone_slave_unit_pcim_sm_data_in_635), .o(n_1099) );
na02f06 g66859_u0 ( .a(n_1290), .b(n_1289), .o(n_9864) );
in01f08 g66861_u0 ( .a(n_16001), .o(n_2453) );
na02f20 g66864_u0 ( .a(n_1509), .b(n_1113), .o(n_4417) );
no02f20 g66865_u0 ( .a(n_430), .b(n_884), .o(n_1415) );
no02s01 g66866_u0 ( .a(n_1201), .b(n_1509), .o(g66866_p) );
in01s01 g66866_u1 ( .a(g66866_p), .o(n_1510) );
no02f10 g66868_u0 ( .a(n_374), .b(n_956), .o(n_1378) );
na02f01 TIMEBOOST_cell_37332 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q), .b(n_4671), .o(TIMEBOOST_net_10278) );
ao12s01 g66870_u0 ( .a(n_1175), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_), .c(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_), .o(n_1098) );
na02f10 g66871_u0 ( .a(n_1290), .b(n_1288), .o(n_9899) );
ao12s02 g66872_u0 ( .a(n_987), .b(pci_target_unit_wishbone_master_read_count_1_), .c(pci_target_unit_wishbone_master_read_count_0_), .o(n_988) );
na03s03 TIMEBOOST_cell_72404 ( .a(g58794_sb), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__Q), .c(TIMEBOOST_net_12263), .o(n_9114) );
no02f40 g66874_u0 ( .a(n_232), .b(n_881), .o(n_1388) );
no02s01 g66875_u0 ( .a(n_1188), .b(n_1290), .o(g66875_p) );
in01s01 g66875_u1 ( .a(g66875_p), .o(n_1287) );
na02f20 g66876_u0 ( .a(n_411), .b(n_1165), .o(g66876_p) );
in01f10 g66876_u1 ( .a(g66876_p), .o(n_1966) );
in01s01 TIMEBOOST_cell_63578 ( .a(wishbone_slave_unit_del_sync_comp_done_reg_main), .o(TIMEBOOST_net_20758) );
na02m01 TIMEBOOST_cell_64112 ( .a(n_13548), .b(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q), .o(TIMEBOOST_net_21042) );
na02f20 g66879_u0 ( .a(n_1113), .b(n_1201), .o(n_4438) );
na02m10 g66880_u0 ( .a(n_1509), .b(n_1195), .o(n_4495) );
ao12m01 g66881_u0 ( .a(n_16860), .b(n_696), .c(n_2092), .o(n_1686) );
na02m20 g66882_u0 ( .a(n_1201), .b(n_1195), .o(n_4505) );
ao12s01 g66883_u0 ( .a(n_703), .b(wishbone_slave_unit_pci_initiator_if_read_count_0_), .c(wishbone_slave_unit_pci_initiator_if_read_count_1_), .o(n_990) );
in01s01 g66884_u0 ( .a(n_2088), .o(n_2328) );
ao12s01 g66885_u0 ( .a(n_2087), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q), .c(n_1041), .o(n_2088) );
no02f20 g66886_u0 ( .a(n_306), .b(n_885), .o(n_1482) );
no02f08 g66887_u0 ( .a(n_404), .b(n_918), .o(n_1479) );
na02f10 g66888_u0 ( .a(n_375), .b(n_994), .o(g66888_p) );
in01f08 g66888_u1 ( .a(g66888_p), .o(n_1357) );
na02f10 g66889_u0 ( .a(n_331), .b(n_994), .o(g66889_p) );
in01f08 g66889_u1 ( .a(g66889_p), .o(n_1414) );
ao12s01 g66891_u0 ( .a(n_546), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_0_), .c(wishbone_slave_unit_pci_initiator_sm_decode_count_1_), .o(n_1204) );
no02f02 g66892_u0 ( .a(n_524), .b(n_939), .o(n_1096) );
na02m02 TIMEBOOST_cell_18606 ( .a(TIMEBOOST_net_5666), .b(n_14839), .o(g52405_db) );
ao12m01 g66894_u0 ( .a(n_2046), .b(parchk_pci_trdy_reg_in), .c(pciu_pciif_stop_reg_in), .o(n_2086) );
na04m06 TIMEBOOST_cell_72839 ( .a(FE_OFN651_n_4508), .b(g65341_sb), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q), .d(TIMEBOOST_net_20249), .o(TIMEBOOST_net_17486) );
no02f06 g66896_u0 ( .a(n_304), .b(n_877), .o(n_1971) );
no02f20 g66897_u0 ( .a(n_191), .b(n_957), .o(n_2967) );
na03m02 TIMEBOOST_cell_72899 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q), .b(g64269_sb), .c(TIMEBOOST_net_12786), .o(n_3904) );
ao12f01 g66899_u0 ( .a(pci_target_unit_del_sync_bc_in_203), .b(pci_target_unit_pci_target_if_norm_prf_en), .c(pci_target_unit_del_sync_bc_in_202), .o(n_639) );
no02f10 g66900_u0 ( .a(n_350), .b(n_874), .o(n_1361) );
na02f08 g66901_u0 ( .a(n_1188), .b(n_1288), .o(n_9823) );
no02m08 g66902_u0 ( .a(n_1118), .b(n_1103), .o(g66902_p) );
in01m04 g66902_u1 ( .a(g66902_p), .o(n_7569) );
in01f08 g66903_u0 ( .a(n_1507), .o(n_1508) );
no02f08 g66905_u0 ( .a(n_1221), .b(n_1408), .o(n_2129) );
ao12f08 g66906_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_mabort2), .b(wishbone_slave_unit_pci_initiator_sm_mabort1), .c(wbu_pciif_frame_out_in), .o(n_2803) );
na02m06 g66908_u0 ( .a(n_1188), .b(n_1289), .o(n_9895) );
no02f20 g66909_u0 ( .a(n_405), .b(n_919), .o(n_1412) );
no02m08 g66911_u0 ( .a(n_996), .b(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q), .o(g66911_p) );
ao12m04 g66911_u1 ( .a(g66911_p), .b(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q), .c(n_996), .o(n_998) );
no02f04 g66912_u0 ( .a(parchk_pci_ad_reg_in_1214), .b(pci_target_unit_pcit_if_strd_addr_in_695), .o(g66912_p) );
ao12f02 g66912_u1 ( .a(g66912_p), .b(pci_target_unit_pcit_if_strd_addr_in_695), .c(parchk_pci_ad_reg_in_1214), .o(n_641) );
no02f20 g66913_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_22__Q), .b(wbu_addr_in_271), .o(g66913_p) );
ao12f08 g66913_u1 ( .a(g66913_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_22__Q), .c(wbu_addr_in_271), .o(n_999) );
no02f04 g66915_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_713), .b(parchk_pci_ad_reg_in_1232), .o(g66915_p) );
ao12f02 g66915_u1 ( .a(g66915_p), .b(pci_target_unit_pcit_if_strd_addr_in_713), .c(parchk_pci_ad_reg_in_1232), .o(n_640) );
ao12f80 g66916_u0 ( .a(n_341), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_), .o(n_872) );
no02f01 g66917_u0 ( .a(pci_target_unit_pcit_if_strd_bc_in_718), .b(n_2648), .o(g66917_p) );
ao12f01 g66917_u1 ( .a(g66917_p), .b(pci_target_unit_pcit_if_strd_bc_in_718), .c(n_2648), .o(n_2036) );
no02m10 g66918_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_712), .b(parchk_pci_ad_reg_in_1231), .o(g66918_p) );
ao12f06 g66918_u1 ( .a(g66918_p), .b(pci_target_unit_pcit_if_strd_addr_in_712), .c(parchk_pci_ad_reg_in_1231), .o(n_627) );
ao22f02 g66920_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_), .c(n_345), .d(n_425), .o(n_1095) );
no02f08 g66921_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_714), .b(parchk_pci_ad_reg_in_1233), .o(g66921_p) );
ao12f04 g66921_u1 ( .a(g66921_p), .b(pci_target_unit_pcit_if_strd_addr_in_714), .c(parchk_pci_ad_reg_in_1233), .o(n_695) );
no02m10 g66922_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_710), .b(parchk_pci_ad_reg_in_1229), .o(g66922_p) );
ao12f06 g66922_u1 ( .a(g66922_p), .b(pci_target_unit_pcit_if_strd_addr_in_710), .c(parchk_pci_ad_reg_in_1229), .o(n_626) );
no02f04 g66923_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_16__Q), .b(wbu_addr_in_265), .o(g66923_p) );
ao12f02 g66923_u1 ( .a(g66923_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_16__Q), .c(wbu_addr_in_265), .o(n_871) );
no02m40 g66924_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_706), .b(parchk_pci_ad_reg_in_1225), .o(g66924_p) );
ao12f10 g66924_u1 ( .a(g66924_p), .b(pci_target_unit_pcit_if_strd_addr_in_706), .c(parchk_pci_ad_reg_in_1225), .o(n_700) );
no02f20 g66925_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_6__Q), .b(wbu_addr_in_255), .o(g66925_p) );
ao12f08 g66925_u1 ( .a(g66925_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_6__Q), .c(wbu_addr_in_255), .o(n_1004) );
ao12f20 g66926_u0 ( .a(n_342), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .o(n_870) );
no02m06 g66927_u0 ( .a(parchk_pci_ad_reg_in_1206), .b(pci_target_unit_pcit_if_strd_addr_in_687), .o(g66927_p) );
ao12m04 g66927_u1 ( .a(g66927_p), .b(pci_target_unit_pcit_if_strd_addr_in_687), .c(parchk_pci_ad_reg_in_1206), .o(n_625) );
ao12s01 g66928_u0 ( .a(n_1266), .b(pci_target_unit_fifos_pcir_whole_waddr_94), .c(n_1174), .o(n_1755) );
no02f10 g66929_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_14__Q), .b(wbu_addr_in_263), .o(g66929_p) );
ao12f06 g66929_u1 ( .a(g66929_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_14__Q), .c(wbu_addr_in_263), .o(n_1007) );
no02f02 g66930_u0 ( .a(n_2651), .b(pci_target_unit_pcit_if_strd_bc_in_717), .o(g66930_p) );
ao12f02 g66930_u1 ( .a(g66930_p), .b(pci_target_unit_pcit_if_strd_bc_in_717), .c(n_2651), .o(n_1754) );
no02f40 g66931_u0 ( .a(wbu_addr_in), .b(wishbone_slave_unit_del_sync_addr_out_reg_0__Q), .o(g66931_p) );
ao12f10 g66931_u1 ( .a(g66931_p), .b(wbu_addr_in), .c(wishbone_slave_unit_del_sync_addr_out_reg_0__Q), .o(n_1008) );
no02f20 g66932_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_23__Q), .b(wbu_addr_in_272), .o(g66932_p) );
ao12f08 g66932_u1 ( .a(g66932_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_23__Q), .c(wbu_addr_in_272), .o(n_950) );
no02f40 g66933_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_27__Q), .b(wbu_addr_in_276), .o(g66933_p) );
ao12f10 g66933_u1 ( .a(g66933_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_27__Q), .c(wbu_addr_in_276), .o(n_869) );
no02f20 g66934_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_690), .b(parchk_pci_ad_reg_in_1209), .o(g66934_p) );
ao12f08 g66934_u1 ( .a(g66934_p), .b(pci_target_unit_pcit_if_strd_addr_in_690), .c(parchk_pci_ad_reg_in_1209), .o(n_708) );
no02f01 g66935_u0 ( .a(n_76), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_), .o(g66935_p) );
ao12f01 g66935_u1 ( .a(g66935_p), .b(n_76), .c(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_), .o(n_868) );
no02f01 g66936_u0 ( .a(pci_target_unit_pcit_if_strd_bc_in_719), .b(n_8511), .o(g66936_p) );
ao12f01 g66936_u1 ( .a(g66936_p), .b(pci_target_unit_pcit_if_strd_bc_in_719), .c(n_8511), .o(n_2042) );
no02f10 g66937_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_699), .b(parchk_pci_ad_reg_in_1218), .o(g66937_p) );
ao12f06 g66937_u1 ( .a(g66937_p), .b(pci_target_unit_pcit_if_strd_addr_in_699), .c(parchk_pci_ad_reg_in_1218), .o(n_624) );
in01f04 g66938_u0 ( .a(FE_OFN197_n_2683), .o(n_2043) );
oa12f06 g66939_u0 ( .a(n_1505), .b(parchk_pci_trdy_en_in), .c(n_34), .o(n_2683) );
no02f20 g66940_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_19__Q), .b(wbu_addr_in_268), .o(g66940_p) );
ao12f10 g66940_u1 ( .a(g66940_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_19__Q), .c(wbu_addr_in_268), .o(n_1012) );
no02f04 g66941_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_715), .b(n_2509), .o(g66941_p) );
ao12f02 g66941_u1 ( .a(g66941_p), .b(pci_target_unit_pcit_if_strd_addr_in_715), .c(n_2509), .o(n_1504) );
no02s06 g66942_u0 ( .a(FE_OCP_RBN2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q), .o(g66942_p) );
ao12m02 g66942_u1 ( .a(g66942_p), .b(FE_OCP_RBN2289_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q), .o(n_1217) );
ao12f06 g66943_u0 ( .a(n_433), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(n_952) );
no02f40 g66944_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_11__Q), .b(wbu_addr_in_260), .o(g66944_p) );
ao12f10 g66944_u1 ( .a(g66944_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_11__Q), .c(wbu_addr_in_260), .o(n_951) );
no02f02 g66945_u0 ( .a(wishbone_slave_unit_fifos_wbr_be_in), .b(wbu_sel_in), .o(g66945_p) );
ao12f02 g66945_u1 ( .a(g66945_p), .b(wishbone_slave_unit_fifos_wbr_be_in), .c(wbu_sel_in), .o(n_711) );
no02f20 g66946_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_17__Q), .b(wbu_addr_in_266), .o(g66946_p) );
ao12f10 g66946_u1 ( .a(g66946_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_17__Q), .c(wbu_addr_in_266), .o(n_867) );
no02f08 g66947_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_711), .b(parchk_pci_ad_reg_in_1230), .o(g66947_p) );
ao12f04 g66947_u1 ( .a(g66947_p), .b(pci_target_unit_pcit_if_strd_addr_in_711), .c(parchk_pci_ad_reg_in_1230), .o(n_623) );
no02f10 g66948_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_701), .b(parchk_pci_ad_reg_in_1220), .o(g66948_p) );
ao12f08 g66948_u1 ( .a(g66948_p), .b(pci_target_unit_pcit_if_strd_addr_in_701), .c(parchk_pci_ad_reg_in_1220), .o(n_622) );
no02f80 g66949_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_24__Q), .b(wbu_addr_in_273), .o(g66949_p) );
ao12f20 g66949_u1 ( .a(g66949_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_24__Q), .c(wbu_addr_in_273), .o(n_866) );
oa12m02 g66950_u0 ( .a(n_1093), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .c(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(n_1094) );
no02f08 g66951_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in), .b(parchk_pci_ad_reg_in), .o(g66951_p) );
ao12f04 g66951_u1 ( .a(g66951_p), .b(pci_target_unit_pcit_if_strd_addr_in), .c(parchk_pci_ad_reg_in), .o(n_621) );
no02f40 g66952_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_10__Q), .b(wbu_addr_in_259), .o(g66952_p) );
ao12f10 g66952_u1 ( .a(g66952_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_10__Q), .c(wbu_addr_in_259), .o(n_865) );
no02f10 g66953_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_698), .b(parchk_pci_ad_reg_in_1217), .o(g66953_p) );
ao12f08 g66953_u1 ( .a(g66953_p), .b(pci_target_unit_pcit_if_strd_addr_in_698), .c(parchk_pci_ad_reg_in_1217), .o(n_658) );
no02f40 g66954_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_29__Q), .b(n_261), .o(g66954_p) );
ao12f10 g66954_u1 ( .a(g66954_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_29__Q), .c(n_261), .o(n_1467) );
no02f40 g66955_u0 ( .a(wbu_addr_in_250), .b(wishbone_slave_unit_del_sync_addr_out_reg_1__Q), .o(g66955_p) );
ao12f10 g66955_u1 ( .a(g66955_p), .b(wbu_addr_in_250), .c(wishbone_slave_unit_del_sync_addr_out_reg_1__Q), .o(n_864) );
ao12f40 g66956_u0 ( .a(n_377), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_), .o(n_863) );
no02f02 g66957_u0 ( .a(wishbone_slave_unit_fifos_wbr_be_in_265), .b(wbu_sel_in_313), .o(g66957_p) );
ao12f02 g66957_u1 ( .a(g66957_p), .b(wishbone_slave_unit_fifos_wbr_be_in_265), .c(wbu_sel_in_313), .o(n_721) );
no02m04 g66959_u0 ( .a(parchk_pci_ad_reg_in_1216), .b(pci_target_unit_pcit_if_strd_addr_in_697), .o(g66959_p) );
ao12f04 g66959_u1 ( .a(g66959_p), .b(pci_target_unit_pcit_if_strd_addr_in_697), .c(parchk_pci_ad_reg_in_1216), .o(n_722) );
no02f06 g66960_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_31__Q), .b(n_539), .o(g66960_p) );
ao12f04 g66960_u1 ( .a(g66960_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_31__Q), .c(n_539), .o(n_1091) );
ao12f80 g66961_u0 ( .a(n_407), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_), .o(n_1016) );
oa12m02 g66962_u0 ( .a(n_1088), .b(n_961), .c(FE_OCP_RBN1930_parchk_pci_trdy_reg_in), .o(n_1089) );
no02f10 g66963_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_703), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(g66963_p) );
ao12f08 g66963_u1 ( .a(g66963_p), .b(pci_target_unit_pcit_if_strd_addr_in_703), .c(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(n_620) );
no02f06 g66964_u0 ( .a(n_3030), .b(pci_target_unit_pcit_if_strd_bc_in), .o(g66964_p) );
ao12f02 g66964_u1 ( .a(g66964_p), .b(pci_target_unit_pcit_if_strd_bc_in), .c(n_3030), .o(n_2297) );
no02f40 g66965_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_26__Q), .b(wbu_addr_in_275), .o(g66965_p) );
ao12f10 g66965_u1 ( .a(g66965_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_26__Q), .c(wbu_addr_in_275), .o(n_1019) );
no02m10 g66966_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_709), .b(parchk_pci_ad_reg_in_1228), .o(g66966_p) );
ao12f06 g66966_u1 ( .a(g66966_p), .b(pci_target_unit_pcit_if_strd_addr_in_709), .c(parchk_pci_ad_reg_in_1228), .o(n_642) );
no02f20 g66968_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_691), .b(parchk_pci_ad_reg_in_1210), .o(g66968_p) );
ao12f08 g66968_u1 ( .a(g66968_p), .b(pci_target_unit_pcit_if_strd_addr_in_691), .c(parchk_pci_ad_reg_in_1210), .o(n_643) );
ao12f80 g66970_u0 ( .a(n_335), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_), .o(n_861) );
no02f08 g66975_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_686), .b(parchk_pci_ad_reg_in_1205), .o(g66975_p) );
ao12f04 g66975_u1 ( .a(g66975_p), .b(pci_target_unit_pcit_if_strd_addr_in_686), .c(parchk_pci_ad_reg_in_1205), .o(n_725) );
ao12f20 g66976_u0 ( .a(n_364), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .o(n_858) );
no02f20 g66978_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_707), .b(parchk_pci_ad_reg_in_1226), .o(g66978_p) );
ao12f08 g66978_u1 ( .a(g66978_p), .b(pci_target_unit_pcit_if_strd_addr_in_707), .c(parchk_pci_ad_reg_in_1226), .o(n_617) );
oa12f01 g66982_u0 ( .a(n_1028), .b(n_1280), .c(pci_target_unit_wishbone_master_rty_counter_1_), .o(n_1281) );
no02f20 g66984_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_705), .b(parchk_pci_ad_reg_in_1224), .o(g66984_p) );
ao12f08 g66984_u1 ( .a(g66984_p), .b(pci_target_unit_pcit_if_strd_addr_in_705), .c(parchk_pci_ad_reg_in_1224), .o(n_645) );
no02f06 g66985_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_704), .b(parchk_pci_ad_reg_in_1223), .o(g66985_p) );
ao12f04 g66985_u1 ( .a(g66985_p), .b(pci_target_unit_pcit_if_strd_addr_in_704), .c(parchk_pci_ad_reg_in_1223), .o(n_729) );
no02f06 g66986_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_692), .b(parchk_pci_ad_reg_in_1211), .o(g66986_p) );
ao12f04 g66986_u1 ( .a(g66986_p), .b(pci_target_unit_pcit_if_strd_addr_in_692), .c(parchk_pci_ad_reg_in_1211), .o(n_616) );
no02m08 g66987_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_696), .b(parchk_pci_ad_reg_in_1215), .o(g66987_p) );
ao12f04 g66987_u1 ( .a(g66987_p), .b(pci_target_unit_pcit_if_strd_addr_in_696), .c(parchk_pci_ad_reg_in_1215), .o(n_615) );
no02f20 g66988_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_21__Q), .b(wbu_addr_in_270), .o(g66988_p) );
ao12f08 g66988_u1 ( .a(g66988_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_21__Q), .c(wbu_addr_in_270), .o(n_855) );
no02s01 g66989_u0 ( .a(pci_target_unit_fifos_pciw_inTransactionCount_0_), .b(n_852), .o(g66989_p) );
ao12s01 g66989_u1 ( .a(g66989_p), .b(pci_target_unit_fifos_pciw_inTransactionCount_0_), .c(n_852), .o(n_853) );
no02f02 g66990_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_28__Q), .b(wbu_addr_in_277), .o(g66990_p) );
ao12f02 g66990_u1 ( .a(g66990_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_28__Q), .c(wbu_addr_in_277), .o(n_851) );
ao12f20 g66991_u0 ( .a(n_408), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(n_850) );
ao12f20 g66993_u0 ( .a(n_230), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(n_849) );
ao12f20 g66995_u0 ( .a(n_340), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .o(n_847) );
no02f06 g66997_u0 ( .a(parchk_pci_ad_reg_in_1213), .b(pci_target_unit_pcit_if_strd_addr_in_694), .o(g66997_p) );
ao12f04 g66997_u1 ( .a(g66997_p), .b(pci_target_unit_pcit_if_strd_addr_in_694), .c(parchk_pci_ad_reg_in_1213), .o(n_614) );
ao12s01 g66999_u0 ( .a(n_1454), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .c(n_1316), .o(n_1752) );
ao12f20 g67000_u0 ( .a(n_409), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .o(n_1031) );
no02f10 g67001_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_702), .b(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(g67001_p) );
ao12f06 g67001_u1 ( .a(g67001_p), .b(pci_target_unit_pcit_if_strd_addr_in_702), .c(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(n_734) );
ao12f80 g67002_u0 ( .a(n_234), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_), .o(n_845) );
no02f20 g67003_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_5__Q), .b(wbu_addr_in_254), .o(g67003_p) );
ao12f08 g67003_u1 ( .a(g67003_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_5__Q), .c(wbu_addr_in_254), .o(n_844) );
ao12f40 g67004_u0 ( .a(n_268), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_), .o(n_1033) );
no02f02 g67005_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_716), .b(parchk_pci_ad_reg_in_1235), .o(g67005_p) );
ao12f02 g67005_u1 ( .a(g67005_p), .b(pci_target_unit_pcit_if_strd_addr_in_716), .c(parchk_pci_ad_reg_in_1235), .o(n_737) );
no02f10 g67006_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_700), .b(parchk_pci_ad_reg_in_1219), .o(g67006_p) );
ao12f06 g67006_u1 ( .a(g67006_p), .b(pci_target_unit_pcit_if_strd_addr_in_700), .c(parchk_pci_ad_reg_in_1219), .o(n_613) );
ao12f10 g67007_u0 ( .a(n_386), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .o(n_843) );
no02f10 g67008_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_708), .b(parchk_pci_ad_reg_in_1227), .o(g67008_p) );
ao12f08 g67008_u1 ( .a(g67008_p), .b(pci_target_unit_pcit_if_strd_addr_in_708), .c(parchk_pci_ad_reg_in_1227), .o(n_648) );
no02f06 g67010_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_689), .b(parchk_pci_ad_reg_in_1208), .o(g67010_p) );
ao12f04 g67010_u1 ( .a(g67010_p), .b(pci_target_unit_pcit_if_strd_addr_in_689), .c(parchk_pci_ad_reg_in_1208), .o(n_649) );
no02f01 g67011_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_693), .b(parchk_pci_ad_reg_in_1212), .o(g67011_p) );
ao12f02 g67011_u1 ( .a(g67011_p), .b(pci_target_unit_pcit_if_strd_addr_in_693), .c(parchk_pci_ad_reg_in_1212), .o(n_612) );
ao12f40 g67012_u0 ( .a(n_320), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_), .o(n_842) );
no02f80 g67014_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_25__Q), .b(wbu_addr_in_274), .o(g67014_p) );
ao12f20 g67014_u1 ( .a(g67014_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_25__Q), .c(wbu_addr_in_274), .o(n_960) );
no02f40 g67015_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_30__Q), .b(wbu_addr_in_279), .o(g67015_p) );
ao12f10 g67015_u1 ( .a(g67015_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_30__Q), .c(wbu_addr_in_279), .o(n_1034) );
ao12f10 g67016_u0 ( .a(n_420), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(n_841) );
no02s01 g67017_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_), .o(g67017_p) );
ao12m01 g67017_u1 ( .a(g67017_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q), .o(n_840) );
no02s01 g67018_u0 ( .a(n_358), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q), .o(g67018_p) );
ao12s01 g67018_u1 ( .a(g67018_p), .b(n_358), .c(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q), .o(n_1086) );
no02f20 g67019_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_9__Q), .b(wbu_addr_in_258), .o(g67019_p) );
ao12f08 g67019_u1 ( .a(g67019_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_9__Q), .c(wbu_addr_in_258), .o(n_1035) );
no02f40 g67020_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_15__Q), .b(wbu_addr_in_264), .o(g67020_p) );
ao12f10 g67020_u1 ( .a(g67020_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_15__Q), .c(wbu_addr_in_264), .o(n_839) );
no02f40 g67021_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_4__Q), .b(wbu_addr_in_253), .o(g67021_p) );
ao12f10 g67021_u1 ( .a(g67021_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_4__Q), .c(wbu_addr_in_253), .o(n_838) );
no02f40 g67022_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_13__Q), .b(wbu_addr_in_262), .o(g67022_p) );
ao12f10 g67022_u1 ( .a(g67022_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_13__Q), .c(wbu_addr_in_262), .o(n_837) );
no02f04 g67023_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_20__Q), .b(wbu_addr_in_269), .o(g67023_p) );
ao12f02 g67023_u1 ( .a(g67023_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_20__Q), .c(wbu_addr_in_269), .o(n_959) );
no02f02 g67024_u0 ( .a(wishbone_slave_unit_fifos_wbr_be_in_266), .b(wbu_sel_in_314), .o(g67024_p) );
ao12f02 g67024_u1 ( .a(g67024_p), .b(wishbone_slave_unit_fifos_wbr_be_in_266), .c(wbu_sel_in_314), .o(n_611) );
no02f20 g67025_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_2__Q), .b(wbu_addr_in_251), .o(g67025_p) );
ao12f08 g67025_u1 ( .a(g67025_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_2__Q), .c(wbu_addr_in_251), .o(n_836) );
no02f20 g67026_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_18__Q), .b(wbu_addr_in_267), .o(g67026_p) );
ao12f08 g67026_u1 ( .a(g67026_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_18__Q), .c(wbu_addr_in_267), .o(n_742) );
no02f40 g67029_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_688), .b(parchk_pci_ad_reg_in_1207), .o(g67029_p) );
ao12f10 g67029_u1 ( .a(g67029_p), .b(pci_target_unit_pcit_if_strd_addr_in_688), .c(parchk_pci_ad_reg_in_1207), .o(n_610) );
no02f40 g67030_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_8__Q), .b(wbu_addr_in_257), .o(g67030_p) );
ao12f10 g67030_u1 ( .a(g67030_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_8__Q), .c(wbu_addr_in_257), .o(n_744) );
no02f40 g67031_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_12__Q), .b(wbu_addr_in_261), .o(g67031_p) );
ao12f10 g67031_u1 ( .a(g67031_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_12__Q), .c(wbu_addr_in_261), .o(n_743) );
no02f20 g67032_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_7__Q), .b(wbu_addr_in_256), .o(g67032_p) );
ao12f08 g67032_u1 ( .a(g67032_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_7__Q), .c(wbu_addr_in_256), .o(n_833) );
no02f10 g67033_u0 ( .a(wbu_sel_in_312), .b(wishbone_slave_unit_fifos_wbr_be_in_264), .o(g67033_p) );
ao12f06 g67033_u1 ( .a(g67033_p), .b(wishbone_slave_unit_fifos_wbr_be_in_264), .c(wbu_sel_in_312), .o(n_609) );
ao22m06 g67034_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_), .c(n_362), .d(n_397), .o(n_1085) );
oa12s01 g67035_u0 ( .a(n_1038), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .c(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .o(n_1039) );
no02f20 g67036_u0 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_3__Q), .b(wbu_addr_in_252), .o(g67036_p) );
ao12f08 g67036_u1 ( .a(g67036_p), .b(wishbone_slave_unit_del_sync_addr_out_reg_3__Q), .c(wbu_addr_in_252), .o(n_747) );
na02f01 TIMEBOOST_cell_70612 ( .a(TIMEBOOST_net_17329), .b(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_22514) );
na02m02 TIMEBOOST_cell_68878 ( .a(n_4442), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q), .o(TIMEBOOST_net_21647) );
in01f02 g67040_u0 ( .a(FE_OFN989_n_574), .o(g67040_sb) );
na02m02 TIMEBOOST_cell_49222 ( .a(TIMEBOOST_net_14828), .b(g61818_sb), .o(n_8154) );
na03s01 TIMEBOOST_cell_31908 ( .a(configuration_sync_command_bit2), .b(wbu_wb_init_complete_in), .c(n_709), .o(TIMEBOOST_net_343) );
na02m02 TIMEBOOST_cell_30625 ( .a(n_9878), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q), .o(TIMEBOOST_net_9417) );
na02s01 TIMEBOOST_cell_49077 ( .a(TIMEBOOST_net_12726), .b(FE_OFN775_n_15366), .o(TIMEBOOST_net_14756) );
in01s01 g67042_u0 ( .a(conf_pci_init_complete_out), .o(g67042_sb) );
in01s01 TIMEBOOST_cell_63560 ( .a(TIMEBOOST_net_20740), .o(wbs_adr_i_25_) );
na02s01 g67042_u2 ( .a(pci_ad_i_6_), .b(conf_pci_init_complete_out), .o(g67042_db) );
na02s02 g58774_u1 ( .a(wbu_addr_in_265), .b(g58774_sb), .o(g58774_da) );
na02s01 g67043_u2 ( .a(pci_ad_i_8_), .b(conf_pci_init_complete_out), .o(g67043_db) );
na02m01 TIMEBOOST_cell_53409 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q), .b(FE_OFN636_n_4669), .o(TIMEBOOST_net_16922) );
in01f10 g67044_u0 ( .a(parchk_pci_cbe_en_in), .o(g67044_sb) );
na04f04 TIMEBOOST_cell_65710 ( .a(TIMEBOOST_net_7211), .b(FE_OFN1145_n_15261), .c(TIMEBOOST_net_649), .d(g54181_da), .o(TIMEBOOST_net_15817) );
in01s06 TIMEBOOST_cell_67743 ( .a(pci_target_unit_fifos_pcir_data_in_185), .o(TIMEBOOST_net_21170) );
na02f02 g67045_u1 ( .a(pci_cbe_i_1_), .b(g57790_sb), .o(g67045_da) );
na03f04 TIMEBOOST_cell_67000 ( .a(FE_OCP_RBN1998_n_13971), .b(TIMEBOOST_net_16522), .c(FE_OFN1587_n_13736), .o(g53267_p) );
in01f10 g67046_u0 ( .a(parchk_pci_cbe_en_in), .o(g67046_sb) );
in01s01 TIMEBOOST_cell_45959 ( .a(TIMEBOOST_net_13920), .o(TIMEBOOST_net_13871) );
in01s01 TIMEBOOST_cell_45958 ( .a(TIMEBOOST_net_13918), .o(TIMEBOOST_net_13919) );
in01f10 g67047_u0 ( .a(n_1211), .o(n_832) );
in01f10 g67048_u0 ( .a(conf_wb_err_bc_in), .o(g67048_sb) );
na02f02 TIMEBOOST_cell_69057 ( .a(TIMEBOOST_net_21736), .b(g65333_sb), .o(TIMEBOOST_net_10591) );
in01s01 g67049_u0 ( .a(conf_pci_init_complete_out), .o(g67049_sb) );
na02s01 g67049_u2 ( .a(pci_ad_i_19_), .b(conf_pci_init_complete_out), .o(g67049_db) );
na03m02 TIMEBOOST_cell_72673 ( .a(TIMEBOOST_net_14264), .b(FE_OFN955_n_1699), .c(g65791_sb), .o(n_1595) );
na02f04 TIMEBOOST_cell_70762 ( .a(g58261_sb), .b(wbm_adr_o_30_), .o(TIMEBOOST_net_22589) );
na02s01 g67050_u2 ( .a(pci_ad_i_31_), .b(conf_pci_init_complete_out), .o(g67050_db) );
in01f08 g67051_u0 ( .a(FE_OFN989_n_574), .o(g67051_sb) );
na03f10 TIMEBOOST_cell_159 ( .a(n_7044), .b(FE_RN_533_0), .c(n_2883), .o(n_15402) );
na02s01 TIMEBOOST_cell_63229 ( .a(TIMEBOOST_net_20561), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_9346) );
na02m04 TIMEBOOST_cell_53781 ( .a(n_3623), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q), .o(TIMEBOOST_net_17108) );
na02m02 TIMEBOOST_cell_68806 ( .a(TIMEBOOST_net_12389), .b(FE_OFN917_n_4725), .o(TIMEBOOST_net_21611) );
na02m02 TIMEBOOST_cell_70480 ( .a(pci_cbe_o_1_), .b(n_14389), .o(TIMEBOOST_net_22448) );
na02m01 TIMEBOOST_cell_54047 ( .a(n_3739), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q), .o(TIMEBOOST_net_17241) );
na02f02 TIMEBOOST_cell_71435 ( .a(TIMEBOOST_net_22925), .b(n_4871), .o(n_4872) );
na03f06 TIMEBOOST_cell_72515 ( .a(g63548_sb), .b(pci_target_unit_fifos_pciw_addr_data_in), .c(TIMEBOOST_net_23161), .o(TIMEBOOST_net_14834) );
na02m02 TIMEBOOST_cell_49092 ( .a(TIMEBOOST_net_14763), .b(g61900_sb), .o(n_8024) );
na02f02 TIMEBOOST_cell_71583 ( .a(TIMEBOOST_net_22999), .b(n_12362), .o(n_12676) );
in01s01 TIMEBOOST_cell_45901 ( .a(TIMEBOOST_net_13862), .o(TIMEBOOST_net_5281) );
in01f01 g67057_u0 ( .a(n_2373), .o(g67057_sb) );
na03f40 TIMEBOOST_cell_79 ( .a(n_15414), .b(n_16854), .c(n_15417), .o(n_16015) );
na02s01 TIMEBOOST_cell_53636 ( .a(TIMEBOOST_net_17035), .b(FE_OFN231_n_9839), .o(TIMEBOOST_net_9387) );
na02s01 TIMEBOOST_cell_39368 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q), .b(g58369_sb), .o(TIMEBOOST_net_11296) );
na03f02 TIMEBOOST_cell_73434 ( .a(TIMEBOOST_net_17525), .b(FE_OFN1282_n_4097), .c(g62527_sb), .o(n_6521) );
na02s01 TIMEBOOST_cell_30965 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_28__Q), .b(FE_OFN270_n_9836), .o(TIMEBOOST_net_9587) );
na03f02 TIMEBOOST_cell_70546 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q), .b(FE_OFN1127_g64577_p), .c(n_4528), .o(TIMEBOOST_net_22481) );
in01f20 g67064_u0 ( .a(n_1551), .o(n_12179) );
na04m02 TIMEBOOST_cell_73066 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q), .b(FE_OFN699_n_7845), .c(n_2151), .d(g62022_sb), .o(n_7853) );
in01s01 TIMEBOOST_cell_73974 ( .a(wbm_dat_i_7_), .o(TIMEBOOST_net_23539) );
na02f02 TIMEBOOST_cell_45426 ( .a(FE_OFN2202_n_12042), .b(TIMEBOOST_net_13607), .o(TIMEBOOST_net_12038) );
na02f02 TIMEBOOST_cell_70707 ( .a(TIMEBOOST_net_22561), .b(g61835_sb), .o(n_6977) );
na03f02 TIMEBOOST_cell_71146 ( .a(n_4915), .b(n_395), .c(FE_OFN1243_n_4092), .o(TIMEBOOST_net_22781) );
na02m02 TIMEBOOST_cell_64048 ( .a(n_1860), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q), .o(TIMEBOOST_net_21010) );
in01f10 g67070_u0 ( .a(parchk_pci_cbe_en_in), .o(g67070_sb) );
na02s01 TIMEBOOST_cell_48661 ( .a(n_2651), .b(g65235_sb), .o(TIMEBOOST_net_14548) );
na02s01 TIMEBOOST_cell_68509 ( .a(TIMEBOOST_net_21462), .b(g66410_db), .o(n_2527) );
na02m08 TIMEBOOST_cell_52859 ( .a(wbs_dat_i_19_), .b(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q), .o(TIMEBOOST_net_16647) );
na03m02 TIMEBOOST_cell_72416 ( .a(TIMEBOOST_net_23123), .b(TIMEBOOST_net_13993), .c(g61943_sb), .o(TIMEBOOST_net_17290) );
na04m02 TIMEBOOST_cell_73067 ( .a(n_2162), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q), .c(FE_OFN699_n_7845), .d(g61998_sb), .o(n_7899) );
na04f02 TIMEBOOST_cell_72990 ( .a(TIMEBOOST_net_21981), .b(g65953_sb), .c(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q), .d(FE_OFN706_n_8119), .o(TIMEBOOST_net_22274) );
na03f02 TIMEBOOST_cell_73651 ( .a(TIMEBOOST_net_17514), .b(FE_OFN1235_n_6391), .c(g62931_sb), .o(n_6019) );
na02m02 TIMEBOOST_cell_54486 ( .a(TIMEBOOST_net_17460), .b(FE_OFN1219_n_6886), .o(TIMEBOOST_net_15345) );
na02f02 TIMEBOOST_cell_44362 ( .a(TIMEBOOST_net_13075), .b(FE_OFN1133_g64577_p), .o(TIMEBOOST_net_11400) );
na02s01 g67074_u2 ( .a(pci_ad_i_18_), .b(conf_pci_init_complete_out), .o(g67074_db) );
na02s01 g67075_u2 ( .a(pci_ad_i_11_), .b(conf_pci_init_complete_out), .o(g67075_db) );
na02m03 TIMEBOOST_cell_52773 ( .a(pci_target_unit_fifos_pciw_addr_data_in_122), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q), .o(TIMEBOOST_net_16604) );
in01f10 g67080_u0 ( .a(n_1192), .o(n_1436) );
in01f40 g67082_u0 ( .a(parchk_pci_trdy_en_in), .o(g67082_sb) );
na03f02 TIMEBOOST_cell_34875 ( .a(TIMEBOOST_net_9355), .b(FE_OFN1382_n_8567), .c(g57483_sb), .o(n_10334) );
na02s01 g67083_u2 ( .a(pci_ad_i_1_), .b(conf_pci_init_complete_out), .o(g67083_db) );
na04f04 TIMEBOOST_cell_24226 ( .a(n_9041), .b(g57399_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q), .d(FE_OFN1405_n_8567), .o(n_10370) );
na02m02 TIMEBOOST_cell_54474 ( .a(TIMEBOOST_net_17454), .b(FE_OFN1241_n_4092), .o(TIMEBOOST_net_15663) );
na04f04 TIMEBOOST_cell_24229 ( .a(n_9542), .b(g57396_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q), .d(FE_OFN1417_n_8567), .o(n_11345) );
na02s01 g67085_u2 ( .a(pci_ad_i_21_), .b(conf_pci_init_complete_out), .o(g67085_db) );
na03s02 TIMEBOOST_cell_72656 ( .a(TIMEBOOST_net_21121), .b(FE_OFN1015_n_2053), .c(TIMEBOOST_net_14480), .o(TIMEBOOST_net_22352) );
na02f02 TIMEBOOST_cell_70997 ( .a(TIMEBOOST_net_22706), .b(g62995_sb), .o(n_5892) );
na02s02 TIMEBOOST_cell_48860 ( .a(TIMEBOOST_net_14647), .b(g58129_sb), .o(TIMEBOOST_net_10852) );
na03f02 TIMEBOOST_cell_73652 ( .a(TIMEBOOST_net_17457), .b(FE_OFN1213_n_4151), .c(g62974_sb), .o(n_5934) );
na02m02 TIMEBOOST_cell_69809 ( .a(TIMEBOOST_net_22112), .b(TIMEBOOST_net_14680), .o(TIMEBOOST_net_17125) );
in01s01 TIMEBOOST_cell_45902 ( .a(TIMEBOOST_net_13863), .o(TIMEBOOST_net_13862) );
in01m01 g67089_u0 ( .a(n_1536), .o(n_1450) );
ao22f20 g67090_u0 ( .a(pci_stop_i), .b(n_454), .c(n_205), .d(parchk_pci_trdy_en_in), .o(n_1536) );
na03f02 TIMEBOOST_cell_72688 ( .a(TIMEBOOST_net_21411), .b(TIMEBOOST_net_6961), .c(FE_OFN1122_g64577_p), .o(TIMEBOOST_net_22519) );
na04f02 TIMEBOOST_cell_35120 ( .a(wbs_dat_o_21_), .b(g52515_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_120), .d(FE_OFN1472_g52675_p), .o(n_13806) );
na03m06 TIMEBOOST_cell_68650 ( .a(g65070_sb), .b(FE_OFN665_n_4495), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q), .o(TIMEBOOST_net_21533) );
na02s03 TIMEBOOST_cell_43113 ( .a(pci_target_unit_fifos_pcir_data_in_182), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q), .o(TIMEBOOST_net_12451) );
na02f02 TIMEBOOST_cell_71101 ( .a(TIMEBOOST_net_22758), .b(g63145_sb), .o(n_5850) );
na02f02 TIMEBOOST_cell_70507 ( .a(TIMEBOOST_net_22461), .b(g63136_sb), .o(n_4978) );
na03f02 TIMEBOOST_cell_73530 ( .a(n_4205), .b(FE_OFN1697_n_5751), .c(TIMEBOOST_net_20663), .o(n_14817) );
na04m06 TIMEBOOST_cell_72991 ( .a(FE_OFN1046_n_16657), .b(TIMEBOOST_net_12709), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q), .d(g60676_sb), .o(TIMEBOOST_net_16973) );
na04f04 TIMEBOOST_cell_68035 ( .a(n_3233), .b(n_4880), .c(n_3440), .d(FE_OFN1942_n_3241), .o(n_4879) );
na02f01 TIMEBOOST_cell_70340 ( .a(TIMEBOOST_net_17287), .b(FE_OFN2_n_4778), .o(TIMEBOOST_net_22378) );
no02m01 g67095_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .o(g67095_p) );
ao12m01 g67095_u1 ( .a(g67095_p), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .c(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(n_4939) );
no02f40 g67096_u0 ( .a(parchk_pci_ad_out_in_1180), .b(parchk_pci_ad_out_in_1179), .o(g67096_p) );
ao12f20 g67096_u1 ( .a(g67096_p), .b(parchk_pci_ad_out_in_1180), .c(parchk_pci_ad_out_in_1179), .o(n_652) );
no02f40 g67097_u0 ( .a(parchk_pci_ad_reg_in_1231), .b(parchk_pci_ad_reg_in_1230), .o(g67097_p) );
ao12f20 g67097_u1 ( .a(g67097_p), .b(parchk_pci_ad_reg_in_1231), .c(parchk_pci_ad_reg_in_1230), .o(n_607) );
no02f01 g67098_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_), .o(g67098_p) );
ao12f01 g67098_u1 ( .a(g67098_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_), .o(n_1083) );
no02s01 g67099_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_1_), .b(n_321), .o(g67099_p) );
ao12s01 g67099_u1 ( .a(g67099_p), .b(pci_target_unit_del_sync_comp_cycle_count_1_), .c(n_321), .o(n_963) );
no02f80 g67100_u0 ( .a(parchk_pci_ad_out_in_1190), .b(parchk_pci_ad_out_in_1189), .o(g67100_p) );
ao12f40 g67100_u1 ( .a(g67100_p), .b(parchk_pci_ad_out_in_1190), .c(parchk_pci_ad_out_in_1189), .o(n_606) );
no02f80 g67102_u0 ( .a(parchk_pci_ad_out_in_1198), .b(parchk_pci_ad_out_in_1197), .o(g67102_p) );
ao12f40 g67102_u1 ( .a(g67102_p), .b(parchk_pci_ad_out_in_1198), .c(parchk_pci_ad_out_in_1197), .o(n_605) );
no02f80 g67103_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .o(g67103_p) );
ao12f20 g67103_u1 ( .a(g67103_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_), .o(n_604) );
no02f80 g67104_u0 ( .a(parchk_pci_ad_out_in_1194), .b(parchk_pci_ad_out_in_1193), .o(g67104_p) );
ao12f40 g67104_u1 ( .a(g67104_p), .b(parchk_pci_ad_out_in_1194), .c(parchk_pci_ad_out_in_1193), .o(n_603) );
no02f40 g67105_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .o(g67105_p) );
ao12f20 g67105_u1 ( .a(g67105_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .o(n_602) );
no02s01 g67106_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .o(g67106_p) );
ao12m01 g67106_u1 ( .a(g67106_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(n_655) );
no02s01 g67107_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(g67107_p) );
ao12s01 g67107_u1 ( .a(g67107_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(n_829) );
no02s01 g67108_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(g67108_p) );
ao12s01 g67108_u1 ( .a(g67108_p), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .c(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(n_1199) );
no02s01 g67109_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(g67109_p) );
ao12s01 g67109_u1 ( .a(g67109_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q), .c(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(n_971) );
no02f40 g67110_u0 ( .a(parchk_pci_ad_reg_in_1233), .b(parchk_pci_ad_reg_in_1232), .o(g67110_p) );
ao12f20 g67110_u1 ( .a(g67110_p), .b(parchk_pci_ad_reg_in_1233), .c(parchk_pci_ad_reg_in_1232), .o(n_656) );
no02m01 g67111_u0 ( .a(n_46), .b(n_16071), .o(g67111_p) );
ao12m01 g67111_u1 ( .a(g67111_p), .b(n_46), .c(n_16071), .o(n_969) );
no02m01 g67112_u0 ( .a(n_160), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q), .o(g67112_p) );
ao12m01 g67112_u1 ( .a(g67112_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q), .c(n_160), .o(n_973) );
no02f80 g67113_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .o(g67113_p) );
ao12f20 g67113_u1 ( .a(g67113_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_), .o(n_601) );
no02m40 g67114_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_), .o(g67114_p) );
ao12m20 g67114_u1 ( .a(g67114_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_), .o(n_659) );
no02f80 g67115_u0 ( .a(parchk_pci_ad_reg_in_1212), .b(parchk_pci_ad_reg_in_1213), .o(g67115_p) );
ao12f40 g67115_u1 ( .a(g67115_p), .b(parchk_pci_ad_reg_in_1213), .c(parchk_pci_ad_reg_in_1212), .o(n_678) );
no02f40 g67116_u0 ( .a(parchk_pci_ad_reg_in_1219), .b(parchk_pci_ad_reg_in_1218), .o(g67116_p) );
ao12f20 g67116_u1 ( .a(g67116_p), .b(parchk_pci_ad_reg_in_1219), .c(parchk_pci_ad_reg_in_1218), .o(n_600) );
no02s01 g67117_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(g67117_p) );
ao12s01 g67117_u1 ( .a(g67117_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_), .o(n_599) );
no02f40 g67118_u0 ( .a(parchk_pci_ad_reg_in_1227), .b(parchk_pci_ad_reg_in_1226), .o(g67118_p) );
ao12f20 g67118_u1 ( .a(g67118_p), .b(parchk_pci_ad_reg_in_1227), .c(parchk_pci_ad_reg_in_1226), .o(n_674) );
no02s01 g67119_u0 ( .a(conf_wb_err_addr_in_943), .b(conf_wb_err_addr_in_944), .o(g67119_p) );
ao12s01 g67119_u1 ( .a(g67119_p), .b(conf_wb_err_addr_in_943), .c(conf_wb_err_addr_in_944), .o(n_662) );
no02f40 g67120_u0 ( .a(parchk_pci_ad_reg_in_1225), .b(parchk_pci_ad_reg_in_1224), .o(g67120_p) );
ao12f20 g67120_u1 ( .a(g67120_p), .b(parchk_pci_ad_reg_in_1225), .c(parchk_pci_ad_reg_in_1224), .o(n_598) );
no02f80 g67122_u0 ( .a(parchk_pci_ad_reg_in_1211), .b(parchk_pci_ad_reg_in_1210), .o(g67122_p) );
ao12f40 g67122_u1 ( .a(g67122_p), .b(parchk_pci_ad_reg_in_1211), .c(parchk_pci_ad_reg_in_1210), .o(n_597) );
no02f80 g67123_u0 ( .a(parchk_pci_ad_reg_in_1209), .b(parchk_pci_ad_reg_in_1208), .o(g67123_p) );
ao12f40 g67123_u1 ( .a(g67123_p), .b(parchk_pci_ad_reg_in_1209), .c(parchk_pci_ad_reg_in_1208), .o(n_663) );
no02f03 g67125_u0 ( .a(n_1061), .b(n_15854), .o(g67125_p) );
ao12f06 g67125_u1 ( .a(g67125_p), .b(n_15854), .c(n_1061), .o(n_1081) );
no02f40 g67126_u0 ( .a(parchk_pci_ad_reg_in_1214), .b(parchk_pci_ad_reg_in_1215), .o(g67126_p) );
ao12f20 g67126_u1 ( .a(g67126_p), .b(parchk_pci_ad_reg_in_1215), .c(parchk_pci_ad_reg_in_1214), .o(n_664) );
no02f80 g67127_u0 ( .a(parchk_pci_ad_out_in_1192), .b(parchk_pci_ad_out_in_1191), .o(g67127_p) );
ao12f40 g67127_u1 ( .a(g67127_p), .b(parchk_pci_ad_out_in_1192), .c(parchk_pci_ad_out_in_1191), .o(n_666) );
no02f01 g67128_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .o(g67128_p) );
ao12f02 g67128_u1 ( .a(g67128_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_), .o(n_596) );
no02m04 g67129_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(g67129_p) );
ao12m02 g67129_u1 ( .a(g67129_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(n_1079) );
no02f80 g67130_u0 ( .a(parchk_pci_ad_out_in_1172), .b(parchk_pci_ad_out_in_1171), .o(g67130_p) );
ao12f40 g67130_u1 ( .a(g67130_p), .b(parchk_pci_ad_out_in_1172), .c(parchk_pci_ad_out_in_1171), .o(n_595) );
no02s01 g67131_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_), .o(g67131_p) );
ao12s01 g67131_u1 ( .a(g67131_p), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_), .c(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .o(n_669) );
no02f80 g67132_u0 ( .a(parchk_pci_ad_out_in_1196), .b(parchk_pci_ad_out_in_1195), .o(g67132_p) );
ao12f40 g67132_u1 ( .a(g67132_p), .b(parchk_pci_ad_out_in_1196), .c(parchk_pci_ad_out_in_1195), .o(n_667) );
no02f20 g67133_u0 ( .a(FE_OFN1781_parchk_pci_ad_reg_in_1221), .b(parchk_pci_ad_reg_in_1220), .o(g67133_p) );
ao12f10 g67133_u1 ( .a(g67133_p), .b(FE_OFN1781_parchk_pci_ad_reg_in_1221), .c(parchk_pci_ad_reg_in_1220), .o(n_594) );
no02f10 g67134_u0 ( .a(n_2509), .b(parchk_pci_ad_reg_in_1235), .o(g67134_p) );
ao12f10 g67134_u1 ( .a(g67134_p), .b(n_2509), .c(parchk_pci_ad_reg_in_1235), .o(n_593) );
no02f02 g67135_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .o(g67135_p) );
ao12f02 g67135_u1 ( .a(g67135_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_), .o(n_668) );
no02f80 g67136_u0 ( .a(parchk_pci_ad_out_in_1176), .b(parchk_pci_ad_out_in_1175), .o(g67136_p) );
ao12f40 g67136_u1 ( .a(g67136_p), .b(parchk_pci_ad_out_in_1176), .c(parchk_pci_ad_out_in_1175), .o(n_592) );
no02f10 g67138_u0 ( .a(parchk_pci_ad_reg_in_1205), .b(parchk_pci_ad_reg_in), .o(g67138_p) );
ao12f08 g67138_u1 ( .a(g67138_p), .b(parchk_pci_ad_reg_in_1205), .c(parchk_pci_ad_reg_in), .o(n_588) );
no02f40 g67139_u0 ( .a(parchk_pci_ad_out_in_1182), .b(parchk_pci_ad_out_in_1181), .o(g67139_p) );
ao12f20 g67139_u1 ( .a(g67139_p), .b(parchk_pci_ad_out_in_1182), .c(parchk_pci_ad_out_in_1181), .o(n_670) );
no02f10 g67140_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(g67140_p) );
ao12f06 g67140_u1 ( .a(g67140_p), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_), .c(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(n_587) );
no02m02 g67141_u0 ( .a(n_150), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q), .o(g67141_p) );
ao12s02 g67141_u1 ( .a(g67141_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q), .c(n_150), .o(n_826) );
no02s01 g67142_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(g67142_p) );
ao12s01 g67142_u1 ( .a(g67142_p), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .c(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(n_1465) );
no02f80 g67143_u0 ( .a(parchk_pci_ad_out_in_1170), .b(parchk_pci_ad_out_in_1169), .o(g67143_p) );
ao12f40 g67143_u1 ( .a(g67143_p), .b(parchk_pci_ad_out_in_1170), .c(parchk_pci_ad_out_in_1169), .o(n_586) );
na02f02 TIMEBOOST_cell_70509 ( .a(TIMEBOOST_net_22462), .b(g62830_sb), .o(n_5315) );
no02f80 g67145_u0 ( .a(parchk_pci_ad_out_in_1178), .b(parchk_pci_ad_out_in_1177), .o(g67145_p) );
ao12f40 g67145_u1 ( .a(g67145_p), .b(parchk_pci_ad_out_in_1178), .c(parchk_pci_ad_out_in_1177), .o(n_672) );
no02f40 g67146_u0 ( .a(parchk_pci_ad_reg_in_1217), .b(parchk_pci_ad_reg_in_1216), .o(g67146_p) );
ao12f20 g67146_u1 ( .a(g67146_p), .b(parchk_pci_ad_reg_in_1217), .c(parchk_pci_ad_reg_in_1216), .o(n_673) );
na02f02 TIMEBOOST_cell_70511 ( .a(TIMEBOOST_net_22463), .b(g62824_sb), .o(n_5330) );
no02f80 g67148_u0 ( .a(parchk_pci_ad_out_in_1188), .b(parchk_pci_ad_out_in_1187), .o(g67148_p) );
ao12f40 g67148_u1 ( .a(g67148_p), .b(parchk_pci_ad_out_in_1188), .c(parchk_pci_ad_out_in_1187), .o(n_583) );
no02f80 g67149_u0 ( .a(parchk_pci_ad_reg_in_1207), .b(parchk_pci_ad_reg_in_1206), .o(g67149_p) );
ao12f20 g67149_u1 ( .a(g67149_p), .b(parchk_pci_ad_reg_in_1207), .c(parchk_pci_ad_reg_in_1206), .o(n_582) );
no02m02 g67150_u0 ( .a(n_150), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q), .o(g67150_p) );
ao12s02 g67150_u1 ( .a(g67150_p), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q), .c(n_150), .o(n_982) );
no02f80 g67151_u0 ( .a(parchk_pci_ad_out_in_1186), .b(parchk_pci_ad_out_in_1185), .o(g67151_p) );
ao12f40 g67151_u1 ( .a(g67151_p), .b(parchk_pci_ad_out_in_1186), .c(parchk_pci_ad_out_in_1185), .o(n_581) );
no02f80 g67152_u0 ( .a(parchk_pci_ad_out_in_1184), .b(parchk_pci_ad_out_in_1183), .o(g67152_p) );
ao12f40 g67152_u1 ( .a(g67152_p), .b(parchk_pci_ad_out_in_1184), .c(parchk_pci_ad_out_in_1183), .o(n_650) );
no02s01 g67153_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_1_), .b(n_282), .o(g67153_p) );
ao12s01 g67153_u1 ( .a(g67153_p), .b(wishbone_slave_unit_del_sync_comp_cycle_count_1_), .c(n_282), .o(n_983) );
no02f40 g67154_u0 ( .a(parchk_pci_ad_reg_in_1229), .b(parchk_pci_ad_reg_in_1228), .o(g67154_p) );
ao12f20 g67154_u1 ( .a(g67154_p), .b(parchk_pci_ad_reg_in_1229), .c(parchk_pci_ad_reg_in_1228), .o(n_675) );
no02m01 g67155_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_), .o(g67155_p) );
ao12m01 g67155_u1 ( .a(g67155_p), .b(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_), .c(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_), .o(n_580) );
no02s01 g67156_u0 ( .a(parchk_pci_cbe_out_in_1203), .b(parchk_pci_cbe_out_in_1202), .o(g67156_p) );
ao12s01 g67156_u1 ( .a(g67156_p), .b(parchk_pci_cbe_out_in_1203), .c(parchk_pci_cbe_out_in_1202), .o(n_676) );
no02f40 g67157_u0 ( .a(parchk_pci_ad_reg_in_1223), .b(FE_OFN1777_parchk_pci_ad_reg_in_1222), .o(g67157_p) );
ao12f20 g67157_u1 ( .a(g67157_p), .b(parchk_pci_ad_reg_in_1223), .c(FE_OFN1777_parchk_pci_ad_reg_in_1222), .o(n_677) );
in01f03 g67176_u0 ( .a(n_2031), .o(n_2520) );
in01s20 g67185_u0 ( .a(n_2597), .o(n_2031) );
in01f40 g67231_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_mabort2), .o(n_1459) );
in01s01 g67246_u0 ( .a(wishbone_slave_unit_del_sync_sync_comp_req_pending), .o(n_1460) );
in01s01 g67261_u0 ( .a(pci_target_unit_wishbone_master_burst_chopped_delayed), .o(n_824) );
in01f20 g67306_u0 ( .a(n_1009), .o(n_1509) );
na02f40 g67307_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(n_143), .o(n_1009) );
no02f06 g67308_u0 ( .a(n_689), .b(pci_target_unit_fifos_pcir_whole_waddr_94), .o(n_1118) );
in01s01 g67310_u0 ( .a(n_7426), .o(n_2040) );
na02s01 g67311_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1216), .o(g67311_p) );
in01s02 g67311_u1 ( .a(g67311_p), .o(n_7426) );
in01s01 g67312_u0 ( .a(n_7279), .o(n_2041) );
na02s01 g67313_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1215), .o(g67313_p) );
in01s01 g67313_u1 ( .a(g67313_p), .o(n_7279) );
no02f40 g67314_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(n_242), .o(n_1195) );
in01f02 g67317_u0 ( .a(n_2464), .o(n_7802) );
na02m01 g67318_u0 ( .a(FE_OCPN1854_n_2071), .b(parchk_pci_ad_reg_in_1205), .o(TIMEBOOST_net_5261) );
no02f08 g67319_u0 ( .a(pciu_pciif_stop_reg_in), .b(n_707), .o(n_2685) );
in01f01 g67320_u0 ( .a(n_1014), .o(n_1826) );
na02f40 g67322_u0 ( .a(wishbone_slave_unit_del_sync_req_comp_pending), .b(n_709), .o(n_1014) );
in01m02 g67323_u0 ( .a(n_7269), .o(n_2084) );
na02f01 g67324_u0 ( .a(n_2044), .b(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(g67324_p) );
in01f02 g67324_u1 ( .a(g67324_p), .o(n_7269) );
na02f01 g67325_u0 ( .a(FE_OCPN1855_n_2071), .b(parchk_pci_ad_reg_in_1211), .o(n_3265) );
in01s01 g67326_u0 ( .a(n_7244), .o(n_2083) );
na02s01 g67327_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1229), .o(g67327_p) );
in01s01 g67327_u1 ( .a(g67327_p), .o(n_7244) );
in01s01 g67328_u0 ( .a(n_7285), .o(n_2286) );
na02s01 g67329_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1230), .o(g67329_p) );
in01s01 g67329_u1 ( .a(g67329_p), .o(n_7285) );
in01m01 g67331_u0 ( .a(n_2046), .o(n_2287) );
na02m08 g67332_u0 ( .a(n_15302), .b(n_565), .o(n_2046) );
in01s01 g67333_u0 ( .a(n_1290), .o(n_1218) );
no02f80 g67335_u0 ( .a(n_349), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(n_1290) );
no02f40 g67336_u0 ( .a(n_143), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .o(n_1201) );
na02f01 g67337_u0 ( .a(pciu_pciif_bckp_stop_in), .b(output_backup_trdy_out_reg_Q), .o(n_1512) );
in01m02 g67339_u0 ( .a(n_7287), .o(n_2082) );
na02f01 g67340_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1226), .o(g67340_p) );
in01f02 g67340_u1 ( .a(g67340_p), .o(n_7287) );
na02f40 g67341_u0 ( .a(n_1104), .b(n_16906), .o(n_819) );
na02f10 g67342_u0 ( .a(n_15998), .b(n_15924), .o(n_1408) );
in01s01 g67350_u0 ( .a(n_8540), .o(n_6996) );
na02s01 g67351_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1235), .o(TIMEBOOST_net_5259) );
in01s01 g67352_u0 ( .a(n_7424), .o(n_1746) );
na02s01 g67353_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1217), .o(g67353_p) );
in01s02 g67353_u1 ( .a(g67353_p), .o(n_7424) );
in01f04 g67354_u0 ( .a(n_7806), .o(n_8517) );
na02m01 g67355_u0 ( .a(FE_OCPN1854_n_2071), .b(parchk_pci_ad_reg_in), .o(g67355_p) );
in01f02 g67355_u1 ( .a(g67355_p), .o(n_7806) );
no02m10 g67356_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(n_713) );
in01s01 g67358_u0 ( .a(n_2080), .o(n_7239) );
na02s01 g67359_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1231), .o(n_2080) );
na02m20 g67360_u0 ( .a(n_715), .b(conf_wb_err_bc_in_848), .o(g67360_p) );
in01m06 g67360_u1 ( .a(g67360_p), .o(n_716) );
in01s02 g67362_u0 ( .a(n_2079), .o(n_7234) );
na02s01 g67363_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1232), .o(TIMEBOOST_net_21137) );
na02f10 g67364_u0 ( .a(n_763), .b(n_2078), .o(g67364_p) );
in01f08 g67364_u1 ( .a(g67364_p), .o(n_2609) );
in01m08 g67365_u0 ( .a(n_816), .o(n_817) );
no02m20 g67366_u0 ( .a(n_148), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .o(n_816) );
na02f01 g67367_u0 ( .a(FE_OCPN1855_n_2071), .b(parchk_pci_ad_reg_in_1207), .o(n_3277) );
na02m40 g67369_u0 ( .a(n_653), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(g67369_p) );
in01m20 g67369_u1 ( .a(g67369_p), .o(n_1615) );
in01s01 g67370_u0 ( .a(n_1265), .o(n_1266) );
no02m40 g67371_u0 ( .a(n_1174), .b(pci_target_unit_fifos_pcir_whole_waddr_94), .o(g67371_p) );
in01m10 g67371_u1 ( .a(g67371_p), .o(n_1265) );
na02m10 g67372_u0 ( .a(n_148), .b(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_), .o(n_1283) );
in01s01 g67375_u0 ( .a(n_3280), .o(n_7289) );
na02s01 g67376_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1212), .o(TIMEBOOST_net_5265) );
in01f10 g67377_u0 ( .a(n_1219), .o(n_1220) );
no02f40 g67378_u0 ( .a(n_815), .b(pci_target_unit_pcit_if_strd_bc_in), .o(n_1219) );
na02s01 g67379_u0 ( .a(n_1263), .b(n_705), .o(n_1264) );
in01f40 g67380_u0 ( .a(n_1017), .o(n_980) );
no02f80 g67382_u0 ( .a(n_573), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(n_1017) );
na02s01 g67383_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_7_), .b(n_705), .o(n_1261) );
in01m02 g67385_u0 ( .a(n_7265), .o(n_2077) );
na02f01 g67386_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1224), .o(g67386_p) );
in01f02 g67386_u1 ( .a(g67386_p), .o(n_7265) );
na02s01 g67387_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_6_), .b(n_705), .o(n_1260) );
in01m02 g67388_u0 ( .a(n_7254), .o(n_2076) );
na02f01 g67389_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1227), .o(g67389_p) );
in01f02 g67389_u1 ( .a(g67389_p), .o(n_7254) );
na02f80 g67390_u0 ( .a(n_242), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(g67390_p) );
in01f80 g67390_u1 ( .a(g67390_p), .o(n_1113) );
in01m02 g67391_u0 ( .a(n_7267), .o(n_2075) );
na02f01 g67392_u0 ( .a(n_2044), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(g67392_p) );
in01f02 g67392_u1 ( .a(g67392_p), .o(n_7267) );
in01m02 g67393_u0 ( .a(n_7272), .o(n_2074) );
na02f01 g67394_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1220), .o(g67394_p) );
in01f02 g67394_u1 ( .a(g67394_p), .o(n_7272) );
na02f40 g67396_u0 ( .a(n_349), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(g67396_p) );
in01f20 g67396_u1 ( .a(g67396_p), .o(n_1188) );
na02s01 g67397_u0 ( .a(FE_OCPN1854_n_2071), .b(parchk_pci_ad_reg_in_1210), .o(g67397_p) );
in01s01 g67397_u1 ( .a(g67397_p), .o(n_7792) );
no02m40 g67398_u0 ( .a(n_2), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(n_1288) );
in01s02 g67400_u0 ( .a(n_2072), .o(n_7295) );
na02s01 g67401_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1233), .o(n_2072) );
in01s01 g67402_u0 ( .a(n_7282), .o(n_1743) );
na02s01 g67403_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1214), .o(g67403_p) );
in01s02 g67403_u1 ( .a(g67403_p), .o(n_7282) );
in01f10 g67404_u0 ( .a(n_1197), .o(n_1198) );
no02f40 g67405_u0 ( .a(n_1023), .b(n_551), .o(g67405_p) );
in01f20 g67405_u1 ( .a(g67405_p), .o(n_1197) );
no02s01 g67406_u0 ( .a(n_85), .b(pci_target_unit_pcit_if_strd_bc_in_718), .o(n_661) );
na02s01 g67407_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_5_), .b(n_705), .o(n_1077) );
in01f01 g67409_u0 ( .a(n_2319), .o(n_7800) );
na02f01 g67410_u0 ( .a(FE_OCPN1854_n_2071), .b(parchk_pci_ad_reg_in_1206), .o(TIMEBOOST_net_5263) );
na02f02 g67411_u0 ( .a(n_16685), .b(n_15998), .o(g67411_p) );
in01f02 g67411_u1 ( .a(g67411_p), .o(n_1742) );
na02m02 g67412_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .b(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q), .o(n_1093) );
na02s01 g67413_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_3_), .b(n_705), .o(n_1259) );
in01s01 g67415_u0 ( .a(n_2070), .o(n_7291) );
na02s01 g67416_u0 ( .a(n_1061), .b(n_2509), .o(n_2070) );
in01f04 g67419_u0 ( .a(n_2337), .o(n_8498) );
na02f20 g67421_u0 ( .a(pci_target_unit_del_sync_req_comp_pending), .b(n_373), .o(g67421_p) );
in01s20 g67421_u1 ( .a(g67421_p), .o(n_2337) );
no02s01 g67422_u0 ( .a(n_181), .b(pci_target_unit_pcit_if_strd_bc_in_718), .o(n_671) );
in01f20 g67423_u0 ( .a(n_812), .o(n_813) );
na02f40 g67425_u0 ( .a(n_573), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(g67425_p) );
in01f40 g67425_u1 ( .a(g67425_p), .o(n_812) );
in01f10 g67426_u0 ( .a(n_16326), .o(n_1074) );
in01s01 g67429_u0 ( .a(n_7440), .o(n_1740) );
na02s01 g67430_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1219), .o(g67430_p) );
in01s02 g67430_u1 ( .a(g67430_p), .o(n_7440) );
in01m02 g67431_u0 ( .a(n_7259), .o(n_2069) );
na02f01 g67432_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1225), .o(g67432_p) );
in01f02 g67432_u1 ( .a(g67432_p), .o(n_7259) );
in01f01 g67433_u0 ( .a(n_1027), .o(n_1028) );
na02f40 g67434_u0 ( .a(n_1280), .b(pci_target_unit_wishbone_master_rty_counter_1_), .o(g67434_p) );
in01f20 g67434_u1 ( .a(g67434_p), .o(n_1027) );
in01f06 g67435_u0 ( .a(n_16033), .o(n_1072) );
na02m20 g67437_u0 ( .a(n_2), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(g67437_p) );
in01f10 g67437_u1 ( .a(g67437_p), .o(n_1289) );
na02f01 g67438_u0 ( .a(FE_OCPN1855_n_2071), .b(parchk_pci_ad_reg_in_1209), .o(n_3275) );
in01m01 g67442_u0 ( .a(n_2068), .o(n_7249) );
na02s01 g67443_u0 ( .a(n_1061), .b(parchk_pci_ad_reg_in_1228), .o(n_2068) );
na02s01 g67444_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_4_), .b(n_705), .o(n_1475) );
in01m02 g67445_u0 ( .a(n_7241), .o(n_2067) );
na02f01 g67446_u0 ( .a(n_2044), .b(parchk_pci_ad_reg_in_1223), .o(g67446_p) );
in01f02 g67446_u1 ( .a(g67446_p), .o(n_7241) );
no02f10 g67447_u0 ( .a(n_2316), .b(n_2742), .o(n_2778) );
in01f20 g67448_u0 ( .a(n_15757), .o(n_1221) );
no02s01 g67452_u0 ( .a(n_5755), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(n_1069) );
na02f20 g67453_u0 ( .a(n_689), .b(pci_target_unit_fifos_pcir_whole_waddr_94), .o(g67453_p) );
in01f10 g67453_u1 ( .a(g67453_p), .o(n_1103) );
no02s01 g67454_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_), .o(n_567) );
no02s01 g67456_u0 ( .a(configuration_set_isr_bit2), .b(configuration_sync_isr_2_del_bit_reg_Q), .o(n_1084) );
no02m02 g67457_u0 ( .a(n_16685), .b(n_15998), .o(g67457_p) );
in01f02 g67457_u1 ( .a(g67457_p), .o(n_1739) );
in01s01 g67458_u0 ( .a(n_1453), .o(n_1454) );
no02f20 g67459_u0 ( .a(n_1316), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(g67459_p) );
in01f08 g67459_u1 ( .a(g67459_p), .o(n_1453) );
in01f08 g67460_u0 ( .a(n_992), .o(n_993) );
na02f20 g67461_u0 ( .a(n_16904), .b(n_681), .o(n_992) );
in01s01 g67462_u0 ( .a(n_7231), .o(n_1737) );
na02s01 g67463_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1213), .o(g67463_p) );
in01s02 g67463_u1 ( .a(g67463_p), .o(n_7231) );
no02s01 g67464_u0 ( .a(configuration_set_pci_err_cs_bit8), .b(configuration_sync_pci_err_cs_8_del_bit_reg_Q), .o(n_736) );
no02f01 g67466_u0 ( .a(n_1724), .b(n_2314), .o(n_2315) );
in01s01 g67467_u0 ( .a(n_7422), .o(n_2052) );
na02s01 g67468_u0 ( .a(n_1698), .b(parchk_pci_ad_reg_in_1218), .o(g67468_p) );
in01s02 g67468_u1 ( .a(g67468_p), .o(n_7422) );
na02f20 g67469_u0 ( .a(wishbone_slave_unit_pcim_sm_be_in_558), .b(n_57), .o(n_564) );
in01f10 g67479_u0 ( .a(n_1258), .o(n_2115) );
in01f10 g67480_u0 ( .a(FE_OFN1619_n_1787), .o(n_1258) );
no02f40 g67481_u0 ( .a(n_541), .b(n_504), .o(n_1787) );
na02s01 g67483_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q), .b(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .o(n_1038) );
no02m08 g67484_u0 ( .a(n_763), .b(n_2078), .o(n_3108) );
na02f01 g67485_u0 ( .a(FE_OCPN1855_n_2071), .b(parchk_pci_ad_reg_in_1208), .o(n_3273) );
na02s01 g67486_u0 ( .a(n_123), .b(pci_rst_i), .o(wb_rst_o) );
na02f40 g67487_u0 ( .a(wbu_addr_in_265), .b(wbu_addr_in_262), .o(n_191) );
in01f01 g67488_u0 ( .a(n_560), .o(n_561) );
no02f80 g67489_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_), .o(g67489_p) );
in01f40 g67489_u1 ( .a(g67489_p), .o(n_560) );
no02f80 g67490_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_), .o(n_335) );
na02f02 g67491_u0 ( .a(wbu_addr_in_274), .b(wbu_addr_in_275), .o(n_888) );
in01f20 g67492_u0 ( .a(n_1005), .o(n_1106) );
no02f40 g67493_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(g67493_p) );
in01f20 g67493_u1 ( .a(g67493_p), .o(n_1005) );
na02f10 g67494_u0 ( .a(pciu_am1_in_535), .b(parchk_pci_ad_reg_in_1230), .o(n_336) );
na02f40 g67495_u0 ( .a(pciu_bar1_in_387), .b(pciu_am1_in_525), .o(g67495_p) );
in01f10 g67495_u1 ( .a(g67495_p), .o(n_3404) );
na02m06 TIMEBOOST_cell_52827 ( .a(pci_target_unit_fifos_pciw_addr_data_in_148), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q), .o(TIMEBOOST_net_16631) );
na02f80 g67497_u0 ( .a(wbm_adr_o_15_), .b(wbm_adr_o_16_), .o(n_923) );
no02f04 g67498_u0 ( .a(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q), .b(wishbone_slave_unit_del_sync_comp_rty_exp_reg), .o(g67498_p) );
in01f02 g67498_u1 ( .a(g67498_p), .o(n_559) );
na02f40 g67499_u0 ( .a(conf_wb_err_addr_in_961), .b(conf_wb_err_addr_in_962), .o(n_895) );
na02f02 g67500_u0 ( .a(pci_target_unit_fifos_pcir_whole_waddr_94), .b(pci_target_unit_fifos_pcir_whole_waddr), .o(n_914) );
na02f10 g67501_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_0_), .b(pci_target_unit_wishbone_master_rty_counter_1_), .o(n_1334) );
na02f80 g67502_u0 ( .a(conf_wb_err_addr_in_946), .b(conf_wb_err_addr_in_947), .o(g67502_p) );
in01f40 g67502_u1 ( .a(g67502_p), .o(n_994) );
na02f20 g67503_u0 ( .a(n_539), .b(wbu_am1_in), .o(n_558) );
na02f10 g67504_u0 ( .a(parchk_pci_ad_reg_in_1225), .b(pciu_am1_in_530), .o(n_204) );
na02f40 g67505_u0 ( .a(pciu_am1_in_532), .b(pciu_bar1_in_394), .o(g67505_p) );
in01f20 g67505_u1 ( .a(g67505_p), .o(n_3078) );
na02s06 g67506_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_11_), .b(pci_target_unit_del_sync_comp_cycle_count_12_), .o(g67506_p) );
in01s02 g67506_u1 ( .a(g67506_p), .o(n_1989) );
na02s01 g67507_u0 ( .a(pci_target_unit_pci_target_sm_rd_progress), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(g67507_p) );
in01f02 g67507_u1 ( .a(g67507_p), .o(n_7530) );
na02f02 g67510_u0 ( .a(pciu_am1_in_525), .b(parchk_pci_ad_reg_in_1220), .o(n_290) );
no02f20 g67511_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_), .o(n_340) );
na02f40 g67512_u0 ( .a(wbm_adr_o_21_), .b(wbm_adr_o_22_), .o(n_915) );
no02f80 g67514_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_), .o(g67514_p) );
in01f20 g67514_u1 ( .a(g67514_p), .o(n_1011) );
no02f80 g67515_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_), .o(n_341) );
in01f10 g67518_u0 ( .a(n_562), .o(n_563) );
na02f80 g67519_u0 ( .a(wbm_adr_o_5_), .b(wbm_adr_o_6_), .o(g67519_p) );
in01f40 g67519_u1 ( .a(g67519_p), .o(n_562) );
no02f80 g67520_u0 ( .a(n_16690), .b(n_15998), .o(n_1812) );
na02f02 g67521_u0 ( .a(wbu_addr_in_259), .b(wbu_addr_in_260), .o(n_945) );
na02f08 g67522_u0 ( .a(wbu_addr_in_253), .b(wbu_addr_in_254), .o(n_430) );
na02f01 g67523_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(g67523_p) );
in01f02 g67523_u1 ( .a(g67523_p), .o(n_1115) );
na02f10 g67526_u0 ( .a(pciu_am1_in_526), .b(FE_OFN1780_parchk_pci_ad_reg_in_1221), .o(n_287) );
na02m04 g67527_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q), .b(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_), .o(n_554) );
no02f80 g67528_u0 ( .a(parchk_pci_ad_reg_in), .b(parchk_pci_ad_reg_in_1205), .o(n_343) );
na02f10 g67530_u0 ( .a(wbu_addr_in_253), .b(wbu_addr_in_252), .o(n_350) );
na02m20 g67531_u0 ( .a(wbm_adr_o_27_), .b(wbm_adr_o_28_), .o(g67531_p) );
in01m08 g67531_u1 ( .a(g67531_p), .o(n_879) );
na02m03 g67532_u0 ( .a(pci_target_unit_pci_target_sm_n_2), .b(n_1628), .o(n_1383) );
na02f20 g67533_u0 ( .a(wbu_addr_in_254), .b(wbu_addr_in_255), .o(n_874) );
na02f40 g67534_u0 ( .a(pciu_am1_in_522), .b(pciu_bar1_in_384), .o(g67534_p) );
in01f20 g67534_u1 ( .a(g67534_p), .o(n_2812) );
na02s20 g67535_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_6_), .b(pci_target_unit_del_sync_comp_cycle_count_5_), .o(g67535_p) );
in01s08 g67535_u1 ( .a(g67535_p), .o(n_1690) );
na02f40 g67536_u0 ( .a(pciu_am1_in_520), .b(pciu_bar1_in_382), .o(g67536_p) );
in01f20 g67536_u1 ( .a(g67536_p), .o(n_2818) );
na02f40 g67537_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(g67537_p) );
in01f20 g67537_u1 ( .a(g67537_p), .o(n_1173) );
no02s01 g67538_u0 ( .a(configuration_cache_line_size_reg), .b(configuration_cache_line_size_reg_2996), .o(g67538_p) );
in01s01 g67538_u1 ( .a(g67538_p), .o(n_434) );
na02f08 g67539_u0 ( .a(n_551), .b(n_16695), .o(n_1291) );
na02f80 g67540_u0 ( .a(conf_wb_err_addr_in_962), .b(conf_wb_err_addr_in_963), .o(n_745) );
na02f10 g67542_u0 ( .a(pciu_am1_in_529), .b(parchk_pci_ad_reg_in_1224), .o(n_419) );
no02f40 g67543_u0 ( .a(n_1519), .b(n_15998), .o(n_2016) );
na02f40 g67544_u0 ( .a(pciu_bar1_in_388), .b(pciu_am1_in_526), .o(g67544_p) );
in01f10 g67544_u1 ( .a(g67544_p), .o(n_2869) );
na02f20 g67545_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .b(wishbone_slave_unit_fifos_wbr_whole_waddr), .o(g67545_p) );
in01f20 g67545_u1 ( .a(g67545_p), .o(n_1210) );
in01f04 g67546_u0 ( .a(n_549), .o(n_550) );
na02f06 g67547_u0 ( .a(wbm_adr_o_24_), .b(wbm_adr_o_25_), .o(n_549) );
no02m10 g67548_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .b(wishbone_slave_unit_fifos_wbr_be_in_264), .o(n_235) );
na02f40 g67549_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_1_), .b(pci_target_unit_del_sync_comp_cycle_count_0_), .o(g67549_p) );
in01f10 g67549_u1 ( .a(g67549_p), .o(n_948) );
na02f40 g67550_u0 ( .a(wbm_adr_o_23_), .b(wbm_adr_o_24_), .o(n_924) );
na02f20 g67551_u0 ( .a(parchk_pci_ad_reg_in_1227), .b(pciu_am1_in_532), .o(n_357) );
na02f20 g67553_u0 ( .a(pciu_am1_in_528), .b(parchk_pci_ad_reg_in_1223), .o(n_360) );
na02f40 g67554_u0 ( .a(wbu_addr_in_266), .b(wbu_addr_in_265), .o(n_956) );
na02f20 g67556_u0 ( .a(wbu_addr_in_271), .b(wbu_addr_in_272), .o(n_892) );
no02f01 g67557_u0 ( .a(n_2629), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(n_2313) );
na02m40 g67558_u0 ( .a(wbm_adr_o_14_), .b(wbm_adr_o_15_), .o(n_900) );
na02f40 g67559_u0 ( .a(pciu_bar1_in_402), .b(pciu_am1_in_540), .o(g67559_p) );
in01f20 g67559_u1 ( .a(g67559_p), .o(n_3592) );
no02f08 g67560_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_11_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_12_), .o(n_1993) );
no02m06 g67562_u0 ( .a(pci_target_unit_fifos_pcir_whole_waddr_94), .b(pci_target_unit_fifos_pcir_whole_waddr), .o(n_1318) );
na02f04 g67563_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_bound), .b(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_4869) );
na02f10 g67564_u0 ( .a(wbu_addr_in_267), .b(wbu_addr_in_268), .o(n_927) );
na02f40 g67565_u0 ( .a(wbm_adr_o_10_), .b(wbm_adr_o_11_), .o(n_926) );
in01s01 g67568_u0 ( .a(n_546), .o(n_547) );
no02s01 g67569_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_decode_count_0_), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_1_), .o(n_546) );
in01f01 g67570_u0 ( .a(n_544), .o(TIMEBOOST_net_12240) );
na02f40 g67571_u0 ( .a(conf_wb_err_bc_in_847), .b(conf_wb_err_bc_in_848), .o(n_544) );
in01m02 g67573_u0 ( .a(n_703), .o(n_660) );
no02f03 g67574_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_0_), .b(wishbone_slave_unit_pci_initiator_if_read_count_1_), .o(n_703) );
in01f20 g67576_u0 ( .a(n_15859), .o(n_2354) );
na02s01 g67579_u0 ( .a(configuration_wb_err_cs_bit0), .b(configuration_icr_bit_2961), .o(n_369) );
no02s01 g67580_u0 ( .a(wbu_cache_line_size_in_206), .b(wbu_cache_line_size_in_207), .o(n_802) );
na02f10 g67581_u0 ( .a(wbm_adr_o_26_), .b(wbm_adr_o_27_), .o(g67581_p) );
in01f08 g67581_u1 ( .a(g67581_p), .o(n_875) );
na02f20 g67582_u0 ( .a(conf_wb_err_addr_in_945), .b(conf_wb_err_addr_in_948), .o(g67582_p) );
in01f10 g67582_u1 ( .a(g67582_p), .o(n_331) );
na02f80 g67583_u0 ( .a(n_541), .b(n_324), .o(g67583_p) );
in01f40 g67583_u1 ( .a(g67583_p), .o(n_2122) );
no02s04 g67584_u0 ( .a(pci_target_unit_wishbone_master_read_count_0_), .b(pci_target_unit_wishbone_master_read_count_reg_2__Q), .o(n_3164) );
no02f40 g67585_u0 ( .a(wishbone_slave_unit_wishbone_slave_img_hit_4_), .b(wishbone_slave_unit_wishbone_slave_img_hit_3_), .o(n_370) );
no02f80 g67586_u0 ( .a(wbm_rty_i), .b(wbm_err_i), .o(n_898) );
no02f20 g67588_u0 ( .a(n_629), .b(n_2078), .o(n_3503) );
in01f10 g67589_u0 ( .a(n_730), .o(n_731) );
na02f40 g67590_u0 ( .a(pci_target_unit_pcit_if_strd_bc_in_718), .b(pci_target_unit_pcit_if_strd_bc_in_719), .o(n_730) );
na02f80 g67591_u0 ( .a(wbm_adr_o_9_), .b(wbm_adr_o_8_), .o(n_920) );
na02f20 g67592_u0 ( .a(conf_wb_err_addr_in_944), .b(conf_wb_err_addr_in_945), .o(g67592_p) );
in01f10 g67592_u1 ( .a(g67592_p), .o(n_375) );
na02f80 g67593_u0 ( .a(conf_wb_err_addr_in_955), .b(conf_wb_err_addr_in_956), .o(n_886) );
na02f20 g67594_u0 ( .a(wbu_am2_in), .b(n_539), .o(n_540) );
in01f40 g67595_u0 ( .a(n_538), .o(n_1194) );
no02f40 g67596_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .o(g67596_p) );
in01f40 g67596_u1 ( .a(g67596_p), .o(n_538) );
na02f04 g67598_u0 ( .a(wbu_addr_in_266), .b(wbu_addr_in_267), .o(n_304) );
no02f80 g67599_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_), .o(n_234) );
na02f08 g67600_u0 ( .a(pciu_am1_in_540), .b(parchk_pci_ad_reg_in_1235), .o(g67600_p) );
in01f06 g67600_u1 ( .a(g67600_p), .o(n_372) );
na02f10 g67601_u0 ( .a(wbu_addr_in_267), .b(wbu_addr_in_264), .o(n_374) );
na02f10 g67602_u0 ( .a(wbu_addr_in_269), .b(wbu_addr_in_270), .o(n_909) );
na02f40 g67603_u0 ( .a(conf_wb_err_addr_in_968), .b(conf_wb_err_addr_in_969), .o(g67603_p) );
in01f20 g67603_u1 ( .a(g67603_p), .o(n_1441) );
na02s03 g67604_u0 ( .a(wbs_bte_i_0_), .b(wbs_bte_i_1_), .o(n_382) );
na02f40 g67605_u0 ( .a(pciu_bar1_in_396), .b(pciu_am1_in_534), .o(g67605_p) );
in01f20 g67605_u1 ( .a(g67605_p), .o(n_2833) );
no02f40 g67606_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_), .o(n_268) );
no02s01 g67607_u0 ( .a(wbm_ack_i), .b(wbm_err_i), .o(TIMEBOOST_net_13941) );
na02f40 g67608_u0 ( .a(conf_wb_err_addr_in_957), .b(conf_wb_err_addr_in_958), .o(n_891) );
na02f40 g67610_u0 ( .a(pciu_bar1_in_399), .b(pciu_am1_in_537), .o(g67610_p) );
in01f20 g67610_u1 ( .a(g67610_p), .o(n_2825) );
na02f10 g67611_u0 ( .a(pciu_am1_in), .b(parchk_pci_ad_reg_in_1212), .o(n_376) );
na02f40 g67613_u0 ( .a(pciu_am1_in_519), .b(pciu_bar1_in_381), .o(g67613_p) );
in01f10 g67613_u1 ( .a(g67613_p), .o(n_2822) );
na02f10 g67614_u0 ( .a(wbu_addr_in_264), .b(wbu_addr_in_263), .o(n_957) );
in01s01 g67616_u0 ( .a(n_535), .o(n_536) );
na02s01 g67617_u0 ( .a(wb_int_i), .b(configuration_icr_bit2_0), .o(n_535) );
na02f80 g67618_u0 ( .a(conf_wb_err_addr_in_964), .b(conf_wb_err_addr_in_965), .o(n_746) );
na02f20 g67619_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_1), .b(wishbone_slave_unit_wishbone_slave_c_state), .o(n_943) );
na02m40 g67620_u0 ( .a(wbm_adr_o_13_), .b(wbm_adr_o_12_), .o(n_901) );
no02f40 g67621_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_), .o(n_377) );
na02f20 g67624_u0 ( .a(pci_target_unit_fifos_pciw_whole_waddr), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(g67624_p) );
in01f20 g67624_u1 ( .a(g67624_p), .o(n_1317) );
na02f08 g67625_u0 ( .a(pciu_am1_in_539), .b(n_2509), .o(g67625_p) );
in01f06 g67625_u1 ( .a(g67625_p), .o(n_233) );
na02f40 g67626_u0 ( .a(pciu_bar1_in_398), .b(pciu_am1_in_536), .o(g67626_p) );
in01f20 g67626_u1 ( .a(g67626_p), .o(n_2841) );
na02f10 g67627_u0 ( .a(parchk_pci_ad_reg_in_1214), .b(pciu_am1_in_519), .o(n_439) );
no02m04 g67628_u0 ( .a(n_2308), .b(n_2316), .o(n_2995) );
na02f80 g67629_u0 ( .a(wbm_adr_o_6_), .b(wbm_adr_o_7_), .o(n_919) );
na02f40 g67630_u0 ( .a(conf_wb_err_addr_in_949), .b(conf_wb_err_addr_in_950), .o(n_232) );
na02f40 g67631_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_105), .b(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .o(g67631_p) );
in01f40 g67631_u1 ( .a(g67631_p), .o(n_1107) );
no02f40 g67632_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .b(wishbone_slave_unit_fifos_wbr_be_in_266), .o(n_398) );
no02m20 g67633_u0 ( .a(wbs_cti_i_0_), .b(wbs_cti_i_2_), .o(n_272) );
na02f40 g67634_u0 ( .a(wbm_adr_o_18_), .b(wbm_adr_o_19_), .o(n_911) );
na02f10 g67635_u0 ( .a(wbu_addr_in_257), .b(wbu_addr_in_256), .o(n_893) );
in01f20 g67638_u0 ( .a(n_533), .o(n_534) );
na02f40 g67639_u0 ( .a(conf_wb_err_addr_in_960), .b(conf_wb_err_addr_in_961), .o(n_533) );
in01f04 g67640_u0 ( .a(n_16052), .o(n_1774) );
na02f20 g67642_u0 ( .a(pciu_am1_in_536), .b(parchk_pci_ad_reg_in_1231), .o(n_385) );
na02f40 g67644_u0 ( .a(n_16906), .b(n_391), .o(n_1200) );
no02s40 g67645_u0 ( .a(wbu_cache_line_size_in_211), .b(wbu_cache_line_size_in_210), .o(n_257) );
no02f20 g67646_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_), .o(n_386) );
na02f01 g67647_u0 ( .a(wbu_addr_in_277), .b(wbu_addr_in_276), .o(n_939) );
in01f03 g67651_u0 ( .a(n_1468), .o(n_13354) );
in01f10 g67654_u0 ( .a(n_1468), .o(n_7552) );
in01f06 g67657_u0 ( .a(n_1468), .o(n_7822) );
in01f20 g67662_u0 ( .a(n_1468), .o(n_12595) );
in01f40 g67663_u0 ( .a(n_532), .o(n_1468) );
no02f80 g67666_u0 ( .a(pci_target_unit_pci_target_sm_cnf_progress), .b(n_2314), .o(n_532) );
na02f10 g67667_u0 ( .a(wbm_adr_o_16_), .b(wbm_adr_o_17_), .o(n_921) );
na02f20 g67668_u0 ( .a(parchk_pci_ad_reg_in_1215), .b(pciu_am1_in_520), .o(n_231) );
no02s02 g67669_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_decode_count_1_), .b(wishbone_slave_unit_pci_initiator_sm_decode_count_2_), .o(n_1471) );
na02f20 g67670_u0 ( .a(parchk_pci_ad_reg_in_1217), .b(pciu_am1_in_522), .o(n_389) );
na02f40 g67671_u0 ( .a(pciu_am1_in_538), .b(parchk_pci_ad_reg_in_1233), .o(g67671_p) );
in01f20 g67671_u1 ( .a(g67671_p), .o(n_277) );
na02f40 g67672_u0 ( .a(conf_wb_err_addr_in_956), .b(conf_wb_err_addr_in_957), .o(g67672_p) );
in01f20 g67672_u1 ( .a(g67672_p), .o(n_913) );
no02f80 g67673_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_1), .b(wishbone_slave_unit_wishbone_slave_c_state), .o(n_1432) );
na02f80 g67675_u0 ( .a(pciu_bar1_in_389), .b(pciu_am1_in_527), .o(g67675_p) );
in01f20 g67675_u1 ( .a(g67675_p), .o(n_2866) );
no02f80 g67676_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_), .b(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_), .o(n_1416) );
na02f02 g67677_u0 ( .a(wbu_addr_in_273), .b(wbu_addr_in_272), .o(n_889) );
no02s01 g67678_u0 ( .a(n_1724), .b(n_2311), .o(n_2763) );
na02s02 g67680_u0 ( .a(wbu_bar2_in), .b(wbu_am2_in), .o(g67680_p) );
in01s04 g67680_u1 ( .a(g67680_p), .o(n_1332) );
na02f02 g67682_u0 ( .a(wbu_addr_in_261), .b(wbu_addr_in_262), .o(n_887) );
no02f40 g67684_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .o(n_230) );
in01f08 g67685_u0 ( .a(n_530), .o(n_531) );
na02f40 g67686_u0 ( .a(conf_wb_err_addr_in_967), .b(conf_wb_err_addr_in_968), .o(n_530) );
na02s40 g67688_u0 ( .a(wbu_bar1_in), .b(wbu_am1_in), .o(g67688_p) );
in01m10 g67688_u1 ( .a(g67688_p), .o(n_1330) );
na02f40 g67689_u0 ( .a(pciu_am1_in_530), .b(pciu_bar1_in_392), .o(g67689_p) );
in01f20 g67689_u1 ( .a(g67689_p), .o(n_2828) );
no02f20 g67690_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_), .o(n_420) );
na02f20 g67691_u0 ( .a(wbu_addr_in_259), .b(wbu_addr_in_258), .o(n_894) );
no02f20 g67692_u0 ( .a(n_497), .b(n_1023), .o(n_798) );
no02f01 g67694_u0 ( .a(n_978), .b(n_15302), .o(n_1251) );
no02f10 g67695_u0 ( .a(wbs_err_o), .b(wbs_rty_o), .o(n_3083) );
no02m20 g67698_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_57), .o(n_1440) );
na02f80 g67699_u0 ( .a(conf_wb_err_addr_in_948), .b(conf_wb_err_addr_in_949), .o(g67699_p) );
in01f40 g67699_u1 ( .a(g67699_p), .o(n_1165) );
in01f06 g67700_u0 ( .a(n_528), .o(n_529) );
na02f80 g67701_u0 ( .a(conf_wb_err_addr_in_966), .b(conf_wb_err_addr_in_967), .o(n_528) );
na02f80 g67702_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_3_), .b(n_1263), .o(n_906) );
no02f40 g67703_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .b(wishbone_slave_unit_fifos_wbr_be_in), .o(n_294) );
na02m20 g67704_u0 ( .a(wbm_adr_o_21_), .b(wbm_adr_o_20_), .o(n_910) );
na02f40 g67705_u0 ( .a(wbm_adr_o_9_), .b(wbm_adr_o_10_), .o(n_897) );
no02f20 g67706_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_), .o(n_409) );
na02f40 g67707_u0 ( .a(pciu_bar1_in_397), .b(pciu_am1_in_535), .o(g67707_p) );
in01f20 g67707_u1 ( .a(g67707_p), .o(n_2856) );
no02f04 g67709_u0 ( .a(n_526), .b(wishbone_slave_unit_del_sync_bc_out_reg_1__Q), .o(g67709_p) );
in01f02 g67709_u1 ( .a(g67709_p), .o(n_527) );
na02f80 g67710_u0 ( .a(conf_wb_err_addr_in_953), .b(conf_wb_err_addr_in_954), .o(n_885) );
na02f40 g67712_u0 ( .a(pciu_bar1_in_391), .b(pciu_am1_in_529), .o(g67712_p) );
in01f20 g67712_u1 ( .a(g67712_p), .o(n_2835) );
na02f08 g67713_u0 ( .a(parchk_pci_ad_reg_in_1213), .b(pciu_am1_in_518), .o(n_298) );
na02f10 g67714_u0 ( .a(wbm_adr_o_7_), .b(wbm_adr_o_8_), .o(n_977) );
na02f20 g67715_u0 ( .a(wbu_addr_in_262), .b(wbu_addr_in_263), .o(n_404) );
na02f20 g67716_u0 ( .a(wbm_adr_o_4_), .b(wbm_adr_o_5_), .o(n_405) );
na02f40 g67717_u0 ( .a(wbm_adr_o_17_), .b(wbm_adr_o_18_), .o(n_917) );
no02f80 g67720_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_), .o(n_407) );
no02s06 g67721_u0 ( .a(wbs_adr_i_2_), .b(wbs_adr_i_3_), .o(g67721_p) );
in01s03 g67721_u1 ( .a(g67721_p), .o(n_748) );
na02f10 g67722_u0 ( .a(pciu_am1_in_533), .b(parchk_pci_ad_reg_in_1228), .o(g67722_p) );
in01f08 g67722_u1 ( .a(g67722_p), .o(n_227) );
in01f01 g67723_u0 ( .a(n_8486), .o(n_2483) );
no02f01 g67724_u0 ( .a(n_2314), .b(n_2629), .o(n_8486) );
na02m80 g67725_u0 ( .a(wbs_cyc_i), .b(wbs_stb_i), .o(g67725_p) );
in01f10 g67725_u1 ( .a(g67725_p), .o(n_1347) );
na02f01 g67726_u0 ( .a(wbu_addr_in_279), .b(n_261), .o(n_524) );
no02f40 g67727_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(n_408) );
no02f20 g67730_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_), .o(n_364) );
na02f01 g67731_u0 ( .a(wbu_addr_in_276), .b(wbu_addr_in_275), .o(g67731_p) );
in01f02 g67731_u1 ( .a(g67731_p), .o(n_1285) );
no02f20 g67734_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_), .o(n_342) );
na02f40 g67735_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_5_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_6_), .o(g67735_p) );
in01f20 g67735_u1 ( .a(g67735_p), .o(n_1689) );
in01s02 g67736_u0 ( .a(n_522), .o(n_523) );
na02s04 g67737_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_12_), .b(pci_target_unit_del_sync_comp_cycle_count_13_), .o(n_522) );
na02f40 g67739_u0 ( .a(pciu_bar1_in_395), .b(pciu_am1_in_533), .o(g67739_p) );
in01f20 g67739_u1 ( .a(g67739_p), .o(n_2815) );
in01f20 g67741_u0 ( .a(n_881), .o(n_521) );
na02f80 g67742_u0 ( .a(conf_wb_err_addr_in_951), .b(conf_wb_err_addr_in_952), .o(n_881) );
no02f06 g67744_u0 ( .a(conf_wb_err_bc_in_847), .b(conf_wb_err_bc_in_848), .o(n_329) );
na02f10 g67745_u0 ( .a(n_653), .b(n_1724), .o(g67745_p) );
in01f08 g67745_u1 ( .a(g67745_p), .o(n_7044) );
na02f40 g67746_u0 ( .a(pciu_am1_in_524), .b(pciu_bar1_in_386), .o(g67746_p) );
in01f20 g67746_u1 ( .a(g67746_p), .o(n_2831) );
na02f20 g67747_u0 ( .a(pciu_bar1_in_401), .b(pciu_am1_in_539), .o(g67747_p) );
in01f10 g67747_u1 ( .a(g67747_p), .o(n_2851) );
na02f04 g67748_u0 ( .a(wbu_addr_in_257), .b(wbu_addr_in_258), .o(n_946) );
no02m06 g67749_u0 ( .a(pci_target_unit_wishbone_master_read_count_1_), .b(pci_target_unit_wishbone_master_read_count_0_), .o(n_987) );
no02f40 g67750_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_), .o(n_320) );
no02s01 g67751_u0 ( .a(pci_target_unit_pci_target_sm_n_2), .b(pci_target_unit_pci_target_sm_n_3), .o(n_520) );
na02f20 g67752_u0 ( .a(wbu_addr_in_255), .b(wbu_addr_in_256), .o(n_884) );
na02f40 g67753_u0 ( .a(wbu_addr_in_271), .b(wbu_addr_in_270), .o(n_902) );
na02f20 g67754_u0 ( .a(conf_wb_err_addr_in_950), .b(conf_wb_err_addr_in_951), .o(g67754_p) );
in01f10 g67754_u1 ( .a(g67754_p), .o(n_411) );
na02f08 g67755_u0 ( .a(pciu_am1_in_527), .b(FE_OFN1778_parchk_pci_ad_reg_in_1222), .o(n_300) );
na02f20 g67756_u0 ( .a(wbm_adr_o_19_), .b(wbm_adr_o_20_), .o(n_916) );
na02f40 g67757_u0 ( .a(conf_wb_err_addr_in_958), .b(conf_wb_err_addr_in_959), .o(g67757_p) );
in01f20 g67757_u1 ( .a(g67757_p), .o(n_912) );
na02s01 g67758_u0 ( .a(configuration_sync_command_bit6), .b(conf_pci_init_complete_out), .o(g67758_p) );
in01f02 g67758_u1 ( .a(g67758_p), .o(n_13766) );
na02f20 g67759_u0 ( .a(parchk_pci_ad_reg_in_1218), .b(pciu_am1_in_523), .o(n_413) );
in01m02 g67760_u0 ( .a(n_518), .o(n_519) );
na02f40 g67761_u0 ( .a(wbm_adr_o_26_), .b(wbm_adr_o_25_), .o(n_518) );
no02f40 g67762_u0 ( .a(pci_target_unit_pci_target_sm_n_2), .b(n_1628), .o(n_976) );
no02f80 g67763_u0 ( .a(wishbone_slave_unit_wishbone_slave_img_hit_1_), .b(wishbone_slave_unit_wishbone_slave_img_hit_0_), .o(g67763_p) );
in01f40 g67763_u1 ( .a(g67763_p), .o(n_412) );
no02m10 g67764_u0 ( .a(n_657), .b(pci_target_unit_pcit_if_req_req_pending_in), .o(n_791) );
na02f40 g67765_u0 ( .a(pciu_bar1_in_393), .b(pciu_am1_in_531), .o(g67765_p) );
in01f20 g67765_u1 ( .a(g67765_p), .o(n_2864) );
no02f10 g67766_u0 ( .a(n_16690), .b(n_2078), .o(n_1248) );
na02f01 g67768_u0 ( .a(n_16070), .b(n_440), .o(n_1215) );
na02m40 g67770_u0 ( .a(output_backup_devsel_out_reg_Q), .b(parchk_pci_trdy_en_in), .o(n_1505) );
no02f20 g67771_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .b(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .o(n_1315) );
no02s01 g67772_u0 ( .a(n_961), .b(n_333), .o(n_727) );
na02f04 g67773_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_1), .b(wishbone_slave_unit_wishbone_slave_c_state_2), .o(n_790) );
no02s01 g67774_u0 ( .a(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q), .b(wishbone_slave_unit_wishbone_slave_pref_en_reg_Q), .o(n_665) );
na02f20 g67775_u0 ( .a(parchk_pci_ad_reg_in_1216), .b(pciu_am1_in_521), .o(n_297) );
na02f40 g67778_u0 ( .a(pciu_am1_in_518), .b(pciu_bar1_in_380), .o(g67778_p) );
in01f10 g67778_u1 ( .a(g67778_p), .o(n_2838) );
na02f40 g67779_u0 ( .a(wbu_addr_in_269), .b(wbu_addr_in_268), .o(n_877) );
na02f20 g67780_u0 ( .a(wbu_addr_in_261), .b(wbu_addr_in_260), .o(n_918) );
na02f40 g67783_u0 ( .a(pciu_am1_in_537), .b(parchk_pci_ad_reg_in_1232), .o(g67783_p) );
in01f20 g67783_u1 ( .a(g67783_p), .o(n_302) );
na02f80 g67785_u0 ( .a(wbm_adr_o_11_), .b(wbm_adr_o_12_), .o(n_896) );
no02s20 g67786_u0 ( .a(wbu_cache_line_size_in_208), .b(wbu_cache_line_size_in_209), .o(n_432) );
no02f40 g67787_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_8_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_9_), .o(n_928) );
na02f20 g67788_u0 ( .a(parchk_pci_ad_reg_in_1219), .b(pciu_am1_in_524), .o(n_303) );
na02f04 g67791_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_3_), .b(pci_target_unit_wishbone_master_rty_counter_4_), .o(g67791_p) );
in01f02 g67791_u1 ( .a(g67791_p), .o(n_929) );
na02f20 g67792_u0 ( .a(wbm_adr_o_22_), .b(wbm_adr_o_23_), .o(n_941) );
in01f02 g67793_u0 ( .a(n_512), .o(n_513) );
na02f01 g67794_u0 ( .a(wbu_addr_in_274), .b(wbu_addr_in_273), .o(n_512) );
in01f02 g67797_u0 ( .a(n_16307), .o(n_1057) );
na02f40 g67799_u0 ( .a(pciu_bar1_in_400), .b(pciu_am1_in_538), .o(g67799_p) );
in01f20 g67799_u1 ( .a(g67799_p), .o(n_2854) );
no02f20 g67800_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .b(wishbone_slave_unit_fifos_wbr_be_in_265), .o(n_236) );
no02f02 g67801_u0 ( .a(n_16685), .b(n_15746), .o(n_2125) );
na02m01 g67802_u0 ( .a(n_1111), .b(wishbone_slave_unit_pcim_sm_be_in_557), .o(g67802_p) );
in01m02 g67802_u1 ( .a(g67802_p), .o(n_1013) );
na02f80 g67803_u0 ( .a(conf_wb_err_addr_in_944), .b(conf_wb_err_addr_in_943), .o(n_568) );
na02s10 g67804_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_3_), .b(pci_target_unit_del_sync_comp_cycle_count_4_), .o(g67804_p) );
in01m06 g67804_u1 ( .a(g67804_p), .o(n_1187) );
na02f20 g67805_u0 ( .a(conf_wb_err_addr_in_955), .b(conf_wb_err_addr_in_952), .o(n_306) );
na02m40 g67806_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_4_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_3_), .o(g67806_p) );
in01m10 g67806_u1 ( .a(g67806_p), .o(n_1186) );
na02f80 g67807_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_1_), .b(wishbone_slave_unit_del_sync_comp_cycle_count_0_), .o(g67807_p) );
in01f20 g67807_u1 ( .a(g67807_p), .o(n_947) );
in01m06 g67808_u0 ( .a(n_784), .o(n_785) );
na02m10 g67809_u0 ( .a(n_206), .b(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q), .o(n_784) );
no02f10 g67810_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_), .o(n_433) );
na02f40 g67811_u0 ( .a(conf_wb_err_addr_in_964), .b(conf_wb_err_addr_in_963), .o(n_904) );
na02f40 g67812_u0 ( .a(conf_wb_err_addr_in_965), .b(conf_wb_err_addr_in_966), .o(n_903) );
no02f40 g67813_u0 ( .a(n_3415), .b(pci_target_unit_fifos_pciw_whole_waddr_47), .o(n_1294) );
na02m20 g67814_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_8_), .b(pci_target_unit_del_sync_comp_cycle_count_9_), .o(g67814_p) );
in01f08 g67814_u1 ( .a(g67814_p), .o(n_937) );
na02f02 g67817_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_55), .b(wishbone_slave_unit_fifos_wbw_whole_waddr), .o(n_1109) );
no02f80 g67818_u0 ( .a(n_763), .b(n_15932), .o(n_2392) );
na02f40 g67820_u0 ( .a(conf_wb_err_addr_in_960), .b(conf_wb_err_addr_in_959), .o(n_890) );
na02f80 g67822_u0 ( .a(wbm_adr_o_13_), .b(wbm_adr_o_14_), .o(n_899) );
na02f10 g67823_u0 ( .a(pciu_am1_in_531), .b(parchk_pci_ad_reg_in_1226), .o(n_436) );
na02f10 g67824_u0 ( .a(pciu_am1_in_534), .b(parchk_pci_ad_reg_in_1229), .o(n_307) );
no02f06 g67826_u0 ( .a(wbs_ack_o), .b(n_16635), .o(n_783) );
na02f40 g67827_u0 ( .a(wishbone_slave_unit_wishbone_slave_del_addr_hit), .b(wishbone_slave_unit_wishbone_slave_del_completion_allow), .o(n_319) );
na02f40 g67828_u0 ( .a(pciu_bar1_in), .b(pciu_am1_in), .o(g67828_p) );
in01f10 g67828_u1 ( .a(g67828_p), .o(n_2844) );
in01m08 g67832_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260), .o(n_4403) );
in01f80 g67857_u0 ( .a(wbm_rty_i), .o(n_705) );
in01f20 g67868_u0 ( .a(n_1111), .o(n_2263) );
in01m10 g67877_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243), .o(n_3636) );
in01m10 g67885_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_), .o(n_4280) );
in01m08 g67936_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487), .o(n_28) );
in01f10 g67939_u0 ( .a(wishbone_slave_unit_pcim_sm_last_in), .o(n_5757) );
in01m10 g67945_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258), .o(n_156) );
in01m10 g67948_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_2_), .o(n_9) );
in01m10 g67969_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70), .o(n_4312) );
in01s04 g67991_u0 ( .a(n_689), .o(n_8876) );
in01f40 g67993_u0 ( .a(pci_target_unit_fifos_pcir_whole_waddr), .o(n_689) );
in01s01 g68021_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46), .o(n_3763) );
in01f02 g68029_u0 ( .a(n_1263), .o(n_221) );
in01s01 g68042_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236), .o(n_4399) );
in01f40 g68103_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_0_), .o(n_1280) );
in01s02 g68110_u0 ( .a(wbu_pci_drcomp_pending_in), .o(n_1816) );
in01f80 g68132_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_rdata_selector), .o(n_541) );
in01s01 g68160_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_0_), .o(n_321) );
in01s01 g68163_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582), .o(n_317) );
in01m01 g68172_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_mabort1), .o(n_188) );
in01s01 g68212_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310), .o(n_7373) );
in01s10 g68217_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_), .o(n_362) );
in01f20 g68225_u0 ( .a(n_324), .o(n_13447) );
in01f40 g68229_u0 ( .a(n_324), .o(n_504) );
in01f80 g68230_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_rdata_selector_14), .o(n_324) );
in01m10 g68239_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622), .o(n_323) );
in01m08 g68251_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43), .o(n_95) );
in01f10 g68277_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_), .o(n_276) );
in01f02 g68284_u0 ( .a(wbu_pciif_frame_out_in), .o(n_3022) );
in01s03 g68315_u0 ( .a(pci_target_unit_del_sync_addr_in_204), .o(n_2598) );
in01m06 g68318_u0 ( .a(wishbone_slave_unit_del_sync_req_done_reg), .o(n_325) );
in01m08 g68325_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6), .o(n_75) );
in01s01 g68332_u0 ( .a(pci_target_unit_fifos_inGreyCount_0_), .o(n_42) );
in01m08 g68346_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380), .o(n_74) );
in01s01 g68356_u0 ( .a(pci_frame_o), .o(n_67) );
in01f02 g68368_u0 ( .a(wbs_ack_o), .o(n_779) );
in01f04 g68369_u0 ( .a(n_326), .o(wbs_ack_o) );
in01f80 g68370_u0 ( .a(wbs_ack_o_1307), .o(n_326) );
in01f40 g68381_u0 ( .a(wishbone_slave_unit_wbs_sm_del_req_pending_in), .o(n_709) );
in01s04 g68389_u0 ( .a(pci_target_unit_del_sync_addr_in_209), .o(n_2512) );
in01s01 g68393_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183), .o(n_6) );
in01m08 g68398_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238), .o(n_4396) );
in01m08 g68401_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377), .o(n_139) );
in01m08 g68410_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376), .o(n_3665) );
in01f40 g68420_u0 ( .a(n_525), .o(n_1023) );
in01f80 g68421_u0 ( .a(conf_w_addr_in_939), .o(n_525) );
in01f80 g68423_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr), .o(n_2) );
in01m20 g68426_u0 ( .a(n_2), .o(n_8953) );
in01s01 g68439_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_0_), .o(n_282) );
in01f20 g68448_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_11_), .o(n_193) );
in01s01 g68452_u0 ( .a(configuration_set_isr_bit2), .o(n_72) );
in01m10 g68454_u0 ( .a(pci_target_unit_del_sync_addr_in_210), .o(n_2541) );
in01m10 g68465_u0 ( .a(pci_target_unit_del_sync_addr_in_212), .o(n_2503) );
in01f02 g68472_u0 ( .a(n_2314), .o(n_5755) );
in01f40 g68485_u0 ( .a(n_1061), .o(n_8511) );
in01m10 g68501_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247), .o(n_4410) );
in01f03 g68509_u0 ( .a(wbu_pciif_devsel_reg_in), .o(n_707) );
in01f20 g68515_u0 ( .a(n_551), .o(n_497) );
in01f80 g68516_u0 ( .a(conf_w_addr_in_938), .o(n_551) );
in01s01 g68522_u0 ( .a(n_333), .o(n_447) );
in01s01 g68523_u0 ( .a(parchk_pci_frame_en_in), .o(n_333) );
in01s01 g68548_u0 ( .a(configuration_pci_err_cs_bit0), .o(n_200) );
in01f08 g68550_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_), .o(n_160) );
in01f80 g68572_u0 ( .a(wishbone_slave_unit_fifos_wbw_whole_waddr_56), .o(n_349) );
in01f10 g68604_u0 ( .a(pci_target_unit_fifos_outGreyCount_0_), .o(n_202) );
in01s01 g68613_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237), .o(n_3738) );
in01s06 g68616_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466), .o(n_351) );
in01m06 g68622_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__248), .o(n_0) );
in01f40 g68642_u0 ( .a(wbu_addr_in_280), .o(n_539) );
in01f20 g68652_u0 ( .a(pciu_pciif_bckp_stop_in), .o(n_205) );
in01f08 g68658_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_1), .o(n_279) );
in01f40 g68674_u0 ( .a(parchk_pci_irdy_en_in), .o(n_961) );
in01m10 g68681_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51), .o(n_17) );
in01s03 g68683_u0 ( .a(wbs_bte_i_0_), .o(n_23) );
in01s03 g68703_u0 ( .a(pci_target_unit_del_sync_addr_in), .o(n_2671) );
in01s01 g68707_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309), .o(n_337) );
in01m10 g68759_u0 ( .a(pci_target_unit_del_sync_addr_in_211), .o(n_2507) );
in01f08 g68771_u0 ( .a(wbm_adr_o_2_), .o(n_208) );
in01s10 g68773_u0 ( .a(pci_target_unit_fifos_pciw_outTransactionCount_1_), .o(n_996) );
in01m10 g68776_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_12_), .o(n_206) );
in01f08 g68778_u0 ( .a(n_691), .o(n_692) );
in01m03 g68787_u0 ( .a(wishbone_slave_unit_pci_initiator_if_del_read_req), .o(n_691) );
in01m08 g68814_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358), .o(n_40) );
in01s20 g68832_u0 ( .a(n_2071), .o(n_3030) );
in01m10 g68839_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544), .o(n_263) );
in01m20 g68852_u0 ( .a(n_2648), .o(TIMEBOOST_net_5255) );
in01f40 g68853_u0 ( .a(n_15854), .o(n_2648) );
in01f40 g68866_u0 ( .a(n_573), .o(n_3415) );
in01f80 g68867_u0 ( .a(pci_target_unit_fifos_pciw_whole_waddr), .o(n_573) );
in01m40 g68882_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_), .o(n_148) );
in01m10 g68888_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_), .o(n_345) );
in01s01 g68917_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543), .o(n_354) );
in01f04 g68929_u0 ( .a(n_285), .o(n_574) );
in01f04 g68941_u0 ( .a(n_285), .o(n_2373) );
in01s02 g68942_u0 ( .a(conf_pci_init_complete_out), .o(n_285) );
in01s01 g68949_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in), .o(n_181) );
in01m10 g68961_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359), .o(n_4323) );
in01m08 g68971_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_2__231), .o(n_366) );
in01s01 g68991_u0 ( .a(n_15856), .o(n_2087) );
na02f08 g68_u0 ( .a(n_16566), .b(n_16105), .o(g68_p) );
in01f08 g68_u1 ( .a(g68_p), .o(n_16992) );
in01m08 g69007_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360), .o(n_119) );
in01f20 g69013_u0 ( .a(pci_target_unit_pci_target_if_keep_desconnect_wo_data_set), .o(n_8728) );
in01f40 g69023_u0 ( .a(pci_target_unit_wishbone_master_addr_into_cnt_reg), .o(n_168) );
in01f40 g69033_u0 ( .a(n_1628), .o(n_278) );
in01m10 g69050_u0 ( .a(pci_target_unit_del_sync_addr_in_205), .o(n_2515) );
in01f08 g69063_u0 ( .a(wishbone_slave_unit_wishbone_slave_c_state_2), .o(n_288) );
in01f06 g69074_u0 ( .a(n_15249), .o(n_7114) );
in01m10 g69089_u0 ( .a(pci_target_unit_del_sync_addr_in_207), .o(n_2526) );
in01m10 g69092_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484), .o(n_83) );
in01m08 g69098_u0 ( .a(pci_target_unit_pci_target_sm_wr_progress), .o(n_2311) );
in01f40 g69104_u0 ( .a(pci_target_unit_pcit_if_req_req_pending_in), .o(n_373) );
in01f40 g69114_u0 ( .a(wbu_addr_in_278), .o(n_261) );
in01m02 g69135_u0 ( .a(pciu_pciif_stop_reg_in), .o(n_378) );
in01f10 g69146_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_), .o(n_440) );
in01f40 g69180_u0 ( .a(pci_target_unit_pci_target_sm_n_3), .o(n_61) );
in01f40 g69207_u0 ( .a(wishbone_slave_unit_wishbone_slave_map), .o(n_1323) );
in01f10 g69209_u0 ( .a(n_15331), .o(n_2092) );
in01m08 g69218_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67), .o(n_38) );
in01m10 g69220_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177), .o(n_18) );
in01m08 g69230_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__265), .o(n_50) );
in01s01 g69252_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_3__270), .o(n_271) );
in01f10 g69259_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_), .o(n_76) );
in01f80 g69271_u0 ( .a(n_16284), .o(n_1519) );
in01s01 g69285_u0 ( .a(pci_target_unit_pcit_if_strd_addr_in_686), .o(n_85) );
in01f10 g69321_u0 ( .a(pci_target_unit_pci_target_sm_rd_progress), .o(n_243) );
in01f40 g69337_u0 ( .a(wishbone_slave_unit_pcim_sm_be_in_559), .o(n_57) );
in01f40 g69362_u0 ( .a(pci_target_unit_wbm_sm_pci_tar_burst_ok), .o(n_815) );
in01m10 g69364_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__365), .o(n_4429) );
in01s01 g69369_u0 ( .a(wishbone_slave_unit_pcim_if_del_req_in), .o(n_169) );
in01s10 g69378_u0 ( .a(pci_target_unit_del_sync_comp_rty_exp_reg), .o(n_1817) );
in01m08 g69418_u0 ( .a(wishbone_slave_unit_pcim_if_del_bc_in_382), .o(n_213) );
in01f80 g69428_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_106), .o(n_242) );
in01m10 g69431_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_8_), .o(n_882) );
in01m08 g69436_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522), .o(n_12) );
in01m10 g69457_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249), .o(n_3691) );
in01f01 g69489_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_9_), .o(n_1992) );
in01s03 g69505_u0 ( .a(pci_target_unit_del_sync_addr_in_206), .o(n_2499) );
in01f40 g69532_u0 ( .a(n_657), .o(n_565) );
in01s01 g69534_u0 ( .a(pci_resi_conf_soft_res_in), .o(n_123) );
in01m08 g69550_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_0__153), .o(n_384) );
in01f40 g69558_u0 ( .a(n_763), .o(n_2316) );
in01f80 g69561_u0 ( .a(n_629), .o(n_763) );
in01f80 g69562_u0 ( .a(n_16285), .o(n_629) );
in01m08 g69576_u0 ( .a(wishbone_slave_unit_pcim_if_del_bc_in_383), .o(n_211) );
in01m02 g69593_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_), .o(n_11) );
in01m01 g69609_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374), .o(n_65) );
in01m08 g69632_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509), .o(n_14) );
in01m10 g69640_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178), .o(n_27) );
in01s01 g69643_u0 ( .a(wbu_cache_line_size_in_207), .o(n_292) );
in01f20 g69650_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_), .o(n_135) );
in01m10 g69652_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342), .o(n_84) );
in01m08 g69673_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330), .o(n_26) );
in01m04 g69686_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_), .o(n_150) );
in01f40 g69707_u0 ( .a(n_391), .o(n_1104) );
in01f80 g69708_u0 ( .a(pci_target_unit_wishbone_master_c_state_0_), .o(n_391) );
in01s10 g69724_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_), .o(n_247) );
in01s01 g69746_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621), .o(n_393) );
in01s01 g69749_u0 ( .a(wbs_err_o), .o(n_471) );
in01f06 g69750_u0 ( .a(n_15204), .o(wbs_err_o) );
in01f40 g69754_u0 ( .a(wishbone_slave_unit_fifos_wbr_whole_waddr_104), .o(n_143) );
in01f80 g69761_u0 ( .a(n_1293), .o(n_1316) );
in01f40 g69775_u0 ( .a(n_2509), .o(n_396) );
in01m10 g69786_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583), .o(n_395) );
in01s01 g69794_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_decode_count_0_), .o(n_401) );
in01m10 g69797_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532), .o(n_15) );
in01m10 g69799_u0 ( .a(wishbone_slave_unit_pcim_if_del_we_in), .o(n_4078) );
in01s01 g69804_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465), .o(n_251) );
in01f10 g69834_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_), .o(n_46) );
in01m08 g69845_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56), .o(n_4394) );
in01m10 g69855_u0 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_), .o(n_397) );
in01s01 g69856_u0 ( .a(configuration_wb_err_cs_bit0), .o(n_24) );
in01f20 g69886_u0 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_10_), .o(n_245) );
in01s01 g69888_u0 ( .a(wishbone_slave_unit_fifos_inGreyCount_0_), .o(n_22) );
in01s01 g69901_u0 ( .a(pci_target_unit_pci_target_if_same_read_reg), .o(n_152) );
in01f80 g69904_u0 ( .a(pci_gnt_i), .o(n_47) );
in01s01 g69937_u0 ( .a(pci_devsel_i), .o(n_34) );
in01s01 g69939_u0 ( .a(wbm_cti_o_1_), .o(n_112) );
in01f20 g69962_u0 ( .a(n_2308), .o(n_2742) );
in01f80 g69963_u0 ( .a(n_15924), .o(n_2308) );
in01m01 g70007_u0 ( .a(pci_target_unit_del_sync_addr_in_208), .o(n_2544) );
in01f40 g70023_u0 ( .a(n_1117), .o(n_1174) );
in01s02 g70029_u0 ( .a(pci_target_unit_del_sync_comp_cycle_count_10_), .o(n_207) );
in01f80 g70054_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_), .o(n_104) );
in01s01 g70062_u0 ( .a(n_16175), .o(n_13608) );
in01f40 g70068_u0 ( .a(pci_target_unit_pci_target_sm_cnf_progress), .o(n_653) );
in01f20 g70083_u0 ( .a(n_1724), .o(n_2629) );
in01f40 g70086_u0 ( .a(n_978), .o(n_1724) );
in01m08 g70097_u0 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_1__192), .o(n_255) );
in01s01 g70100_u0 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_3_), .o(n_416) );
in01m20 g70132_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536), .o(n_4273) );
in01s01 g70154_u0 ( .a(wbm_ack_i), .o(n_1183) );
in01f80 g70183_u0 ( .a(pci_target_unit_wishbone_master_c_state_2_), .o(n_681) );
in01s01 g70191_u0 ( .a(FE_OCP_RBN2277_pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_), .o(n_358) );
in01m08 g70203_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__379), .o(n_4343) );
in01s02 g70209_u0 ( .a(pci_target_unit_fifos_pciw_inTransactionCount_1_), .o(n_852) );
in01f10 g70215_u0 ( .a(n_15330), .o(n_696) );
in01f01 g70227_u0 ( .a(wishbone_slave_unit_pcim_if_del_burst_in), .o(n_21) );
in01f04 g70251_u0 ( .a(wishbone_slave_unit_pcim_if_del_bc_in), .o(n_526) );
in01f40 g70258_u0 ( .a(conf_wb_err_bc_in_847), .o(n_715) );
in01f01 g70269_u0 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_), .o(n_425) );
in01s04 g70281_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271), .o(n_424) );
in01m10 g70305_u0 ( .a(n_1698), .o(n_2651) );
in01s40 g70310_u0 ( .a(parchk_pci_cbe_reg_in_1236), .o(n_1698) );
in01s01 g70414_u0 ( .a(pci_target_unit_pci_target_sm_rd_request), .o(n_177) );
in01m10 g70418_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62), .o(n_3608) );
in01m10 g70425_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__363), .o(n_3672) );
in01m10 g70441_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47), .o(n_36) );
in01m10 g70451_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59), .o(n_3616) );
in01f10 g70465_u0 ( .a(parchk_pci_trdy_en_in), .o(n_454) );
na02f04 g70_u0 ( .a(n_8860), .b(n_16566), .o(g70_p) );
in01f06 g70_u1 ( .a(g70_p), .o(n_15534) );
no02f02 g71_u0 ( .a(n_12151), .b(n_10669), .o(n_15527) );
in01f01 g73860_u0 ( .a(n_14967), .o(n_14965) );
in01f06 g73876_u0 ( .a(FE_OCPN1827_n_14995), .o(n_15001) );
na02f10 g73889_u0 ( .a(n_16311), .b(n_16394), .o(n_16798) );
na03f02 TIMEBOOST_cell_73531 ( .a(TIMEBOOST_net_17473), .b(FE_OFN1242_n_4092), .c(g63108_sb), .o(n_5854) );
no02f10 g73934_u0 ( .a(n_16287), .b(n_1408), .o(n_15125) );
no02f10 g73935_u0 ( .a(n_16291), .b(n_16033), .o(n_15128) );
na02f04 g73947_u0 ( .a(n_16156), .b(n_15388), .o(n_15142) );
oa12m02 g73970_u0 ( .a(n_15196), .b(n_15187), .c(FE_OFN2164_n_16301), .o(n_15197) );
ao12f02 g73971_u0 ( .a(n_14730), .b(n_14800), .c(wbm_dat_o_10_), .o(n_15187) );
na02f01 TIMEBOOST_cell_26099 ( .a(pci_target_unit_pcit_if_strd_addr_in_706), .b(FE_OFN785_n_2678), .o(TIMEBOOST_net_7154) );
na02f02 g73977_u0 ( .a(FE_OFN2164_n_16301), .b(wbm_dat_o_10_), .o(n_15196) );
in01f80 g73986_u0 ( .a(wbs_err_o_1309), .o(n_15204) );
no02f08 g73989_u0 ( .a(n_16284), .b(n_16285), .o(g73989_p) );
in01f08 g73989_u1 ( .a(g73989_p), .o(n_15210) );
in01f02 g73996_u0 ( .a(n_15389), .o(n_15217) );
in01f40 g74023_u0 ( .a(n_16501), .o(n_15249) );
na02f20 g74027_u0 ( .a(n_15260), .b(wishbone_slave_unit_pci_initiator_if_posted_write_req), .o(n_15261) );
na02f20 g74028_u0 ( .a(n_4718), .b(n_15805), .o(g74028_p) );
in01f20 g74028_u1 ( .a(g74028_p), .o(n_15260) );
in01f10 g74031_u0 ( .a(n_15260), .o(n_15262) );
na02f02 g74037_u0 ( .a(n_15994), .b(n_15275), .o(n_15276) );
in01f20 g74038_u0 ( .a(n_16287), .o(n_15275) );
in01f06 g74050_u0 ( .a(n_16002), .o(n_15291) );
na02m02 TIMEBOOST_cell_69618 ( .a(n_4447), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q), .o(TIMEBOOST_net_22017) );
na02f02 g74059_u0 ( .a(n_15614), .b(n_15292), .o(n_15301) );
in01s20 g74061_u0 ( .a(n_15295), .o(n_15302) );
na02s01 TIMEBOOST_cell_45191 ( .a(n_739), .b(wbu_addr_in_252), .o(TIMEBOOST_net_13490) );
no02f80 g74074_u0 ( .a(n_16964), .b(n_15313), .o(n_15314) );
in01f80 g74075_u0 ( .a(wbs_stb_i), .o(n_15313) );
na04f02 TIMEBOOST_cell_35122 ( .a(wbs_dat_o_12_), .b(g52506_sb), .c(wbs_wbb3_2_wbb2_dat_o_i_111), .d(FE_OFN1471_g52675_p), .o(n_13724) );
na02f80 g74082_u0 ( .a(n_2447), .b(n_2392), .o(n_15324) );
in01f20 g74087_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_1_), .o(n_15330) );
in01f20 g74088_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_0_), .o(n_15331) );
no02f80 g74121_u0 ( .a(parchk_pci_frame_en_in), .b(parchk_pci_frame_reg_in), .o(n_15365) );
in01f10 g74122_u0 ( .a(parchk_pci_frame_reg_in), .o(n_15295) );
na02f04 g74124_u0 ( .a(n_16560), .b(n_15372), .o(n_15373) );
no02f04 g74126_u0 ( .a(n_15370), .b(n_15371), .o(n_15372) );
in01f02 g74129_u0 ( .a(n_15371), .o(n_15376) );
na02f80 g74140_u0 ( .a(pci_target_unit_wishbone_master_rty_counter_5_), .b(pci_target_unit_wishbone_master_rty_counter_7_), .o(g74140_p) );
in01f40 g74140_u1 ( .a(g74140_p), .o(n_15385) );
na02f04 g74141_u0 ( .a(n_16980), .b(n_1445), .o(n_15388) );
na02f40 g74142_u0 ( .a(n_16154), .b(n_16150), .o(n_15390) );
in01f10 g74147_u0 ( .a(n_16495), .o(n_15397) );
na02f01 g74153_u0 ( .a(n_1724), .b(pci_target_unit_pci_target_sm_same_read_reg), .o(g74153_p) );
in01f02 g74153_u1 ( .a(g74153_p), .o(n_15405) );
na02f10 g74154_u0 ( .a(pci_target_unit_pci_target_sm_rd_from_fifo), .b(FE_OCPN1836_n_16798), .o(g74154_p) );
in01f08 g74154_u1 ( .a(g74154_p), .o(n_15406) );
no02f02 g74155_u0 ( .a(n_1435), .b(pci_target_unit_pci_target_sm_cnf_progress), .o(n_15407) );
na02f10 g74162_dup_u0 ( .a(n_16949), .b(n_16635), .o(g74162_dup_p) );
in01f10 g74162_dup_u1 ( .a(g74162_dup_p), .o(n_16855) );
na02f02 TIMEBOOST_cell_18457 ( .a(g75418_da), .b(g75418_db), .o(TIMEBOOST_net_5592) );
no02f20 g74173_u0 ( .a(n_15446), .b(n_15467), .o(n_15442) );
na02f04 g74174_u0 ( .a(n_15065), .b(n_2129), .o(g74174_p) );
in01f08 g74174_u1 ( .a(g74174_p), .o(n_15444) );
na02s01 TIMEBOOST_cell_43045 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q), .b(FE_OFN603_n_9687), .o(TIMEBOOST_net_12417) );
na02s01 TIMEBOOST_cell_51573 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q), .o(TIMEBOOST_net_16004) );
in01f06 g74183_u0 ( .a(n_16160), .o(n_15456) );
na02f20 g74191_u0 ( .a(n_15918), .b(n_15908), .o(n_15467) );
no02f10 g74197_u0 ( .a(n_15924), .b(n_15998), .o(n_15474) );
no02f04 g74218_u0 ( .a(n_15514), .b(n_15515), .o(n_15516) );
na03s02 TIMEBOOST_cell_73333 ( .a(FE_OFN229_n_9120), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q), .c(TIMEBOOST_net_20510), .o(TIMEBOOST_net_16995) );
na02s01 TIMEBOOST_cell_39185 ( .a(TIMEBOOST_net_11204), .b(g58040_db), .o(n_9748) );
in01f08 g74222_u0 ( .a(n_15514), .o(n_15517) );
in01f20 g74224_u0 ( .a(n_15518), .o(n_8747) );
no02f20 g74225_u0 ( .a(n_15397), .b(n_15403), .o(n_15518) );
ao12f02 g74239_u0 ( .a(n_15553), .b(n_14918), .c(n_16810), .o(n_16853) );
na02f02 g74240_u0 ( .a(n_15549), .b(n_15552), .o(n_15553) );
ao22f02 g74241_u0 ( .a(n_2831), .b(FE_OCPN1845_n_16427), .c(FE_OFN1063_n_15808), .d(configuration_pci_err_data_516), .o(n_15549) );
ao12f02 g74242_u0 ( .a(n_15551), .b(FE_OFN1069_n_15729), .c(configuration_wb_err_data_585), .o(n_15552) );
na02f04 g74243_u0 ( .a(n_16791), .b(pciu_bar0_in_363), .o(g74243_p) );
in01f02 g74243_u1 ( .a(g74243_p), .o(n_15551) );
no02f02 g74245_u0 ( .a(n_15594), .b(n_11739), .o(g74245_p) );
in01f02 g74245_u1 ( .a(g74245_p), .o(n_15565) );
oa22f01 g74248_u0 ( .a(n_15560), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252), .c(n_16572), .d(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291), .o(n_15562) );
in01f08 g74249_u0 ( .a(FE_OFN1502_n_15558), .o(n_15560) );
in01f08 g74251_u0 ( .a(n_16572), .o(n_15566) );
in01f08 g74252_u0 ( .a(n_15560), .o(n_15568) );
na02f02 g74266_u0 ( .a(n_9305), .b(n_15584), .o(n_15585) );
na02f02 g74267_u0 ( .a(FE_OFN1529_n_10853), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q), .o(n_15584) );
in01f06 g74268_u0 ( .a(FE_OFN1508_n_15587), .o(n_15589) );
na02f06 g74270_u0 ( .a(n_8867), .b(n_8866), .o(g74270_p) );
in01f04 g74270_u1 ( .a(g74270_p), .o(n_15587) );
na02f02 g74272_u0 ( .a(n_10144), .b(n_10728), .o(n_15592) );
na02f02 g74283_u0 ( .a(n_978), .b(n_15295), .o(g74283_p) );
in01f03 g74283_u1 ( .a(g74283_p), .o(n_15607) );
oa12f02 g74287_u0 ( .a(n_15607), .b(n_8819), .c(n_1513), .o(n_15614) );
in01f04 g74313_u0 ( .a(n_15373), .o(n_15638) );
in01f06 g74317_u0 ( .a(n_16560), .o(n_15645) );
na02f80 g74343_u0 ( .a(n_16871), .b(n_16864), .o(n_16940) );
no02f80 g74346_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_1_), .b(wishbone_slave_unit_pci_initiator_sm_cur_state_0_), .o(n_15680) );
no02f02 g74357_u0 ( .a(n_15919), .b(n_16911), .o(n_15689) );
ao12f02 g74359_u0 ( .a(n_15698), .b(n_14917), .c(n_16810), .o(n_15699) );
ao12f04 g74361_u0 ( .a(n_15694), .b(FE_OFN1069_n_15729), .c(configuration_wb_err_data_584), .o(n_15695) );
na02f08 g74363_u0 ( .a(n_16791), .b(pciu_bar0_in_362), .o(g74363_p) );
in01f04 g74363_u1 ( .a(g74363_p), .o(n_15694) );
na02s01 TIMEBOOST_cell_52777 ( .a(g58267_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q), .o(TIMEBOOST_net_16606) );
in01f02 g74388_u0 ( .a(n_15732), .o(n_15733) );
na03f02 TIMEBOOST_cell_73653 ( .a(TIMEBOOST_net_17398), .b(FE_OFN1207_n_6356), .c(g62986_sb), .o(n_5910) );
na03s01 TIMEBOOST_cell_41727 ( .a(g58425_sb), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q), .c(g58425_db), .o(n_9423) );
no02f40 g74406_u0 ( .a(n_1828), .b(n_1829), .o(n_15736) );
no02f20 g74407_u0 ( .a(n_15859), .b(n_15738), .o(n_15739) );
no02f10 g74408_u0 ( .a(wishbone_slave_unit_pci_initiator_if_del_read_req), .b(wishbone_slave_unit_pci_initiator_if_err_recovery), .o(g74408_p) );
in01f10 g74408_u1 ( .a(g74408_p), .o(n_15738) );
in01s01 g74409_u0 ( .a(wishbone_slave_unit_pci_initiator_if_err_recovery), .o(n_15741) );
na02f80 g74416_u0 ( .a(n_525), .b(n_2078), .o(n_15744) );
in01f04 g74423_u0 ( .a(n_15754), .o(n_15756) );
in01f20 g74424_u0 ( .a(n_15744), .o(n_15757) );
in01f06 g74428_u0 ( .a(n_8820), .o(n_15758) );
na02f02 g74429_u0 ( .a(n_4635), .b(n_3810), .o(g74429_p) );
in01f02 g74429_u1 ( .a(g74429_p), .o(n_15759) );
in01f04 g74430_u0 ( .a(n_2416), .o(n_15760) );
no02f20 g74433_u0 ( .a(n_1536), .b(n_1436), .o(n_15762) );
in01m40 g74434_u0 ( .a(parchk_pci_frame_en_in), .o(g74434_sb) );
in01f01 g74437_u0 ( .a(n_15758), .o(n_15769) );
no02s01 g74455_u0 ( .a(n_3320), .b(n_16512), .o(n_15788) );
no02f10 g74470_u0 ( .a(n_16763), .b(wishbone_slave_unit_pcim_sm_rdy_in), .o(g74470_p) );
in01f08 g74470_u1 ( .a(g74470_p), .o(n_15802) );
no02f40 g74471_u0 ( .a(wbu_pciif_devsel_reg_in), .b(parchk_pci_trdy_reg_in), .o(n_15805) );
no02f80 g74472_u0 ( .a(n_15988), .b(n_16936), .o(n_4718) );
na02f10 g74475_u0 ( .a(n_15128), .b(n_15125), .o(g74475_p) );
in01f10 g74475_u1 ( .a(g74475_p), .o(n_15808) );
na03f02 TIMEBOOST_cell_66937 ( .a(FE_OFN1753_n_12086), .b(TIMEBOOST_net_16013), .c(FE_OFN2210_n_11027), .o(n_12611) );
in01f40 g74518_u0 ( .a(parchk_pci_cbe_reg_in_1237), .o(n_15854) );
na02m80 g74520_u0 ( .a(n_1238), .b(n_15856), .o(n_15859) );
in01f80 g74522_u0 ( .a(wishbone_slave_unit_pci_initiator_if_del_write_req), .o(n_15856) );
na02f20 g74553_u0 ( .a(n_16462), .b(n_15824), .o(g74553_p) );
in01f10 g74553_u1 ( .a(g74553_p), .o(n_16599) );
na03f02 TIMEBOOST_cell_73790 ( .a(FE_OFN1602_n_13995), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q), .c(n_14163), .o(n_14481) );
in01f04 g74563_u1 ( .a(g74563_p), .o(n_15910) );
na02f20 g74573_u0 ( .a(FE_OCP_RBN2222_n_15347), .b(n_319), .o(n_15918) );
na02f08 g74575_u0 ( .a(n_16015), .b(n_16016), .o(n_15920) );
in01f20 g74576_u1 ( .a(g74576_p), .o(n_15931) );
na03f02 TIMEBOOST_cell_65164 ( .a(TIMEBOOST_net_16248), .b(g64144_sb), .c(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q), .o(TIMEBOOST_net_17323) );
na02f02 TIMEBOOST_cell_63049 ( .a(TIMEBOOST_net_20471), .b(FE_OFN1136_g64577_p), .o(TIMEBOOST_net_15128) );
na02f20 g74580_u0 ( .a(n_2016), .b(n_798), .o(g74580_p) );
in01f10 g74580_u1 ( .a(g74580_p), .o(n_15922) );
no02f20 g74581_u0 ( .a(n_16690), .b(n_629), .o(n_15923) );
in01f80 g74583_u0 ( .a(conf_w_addr_in_932), .o(n_15924) );
na02s01 TIMEBOOST_cell_18557 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q), .b(FE_OFN2079_n_8069), .o(TIMEBOOST_net_5642) );
in01f40 g74586_u0 ( .a(n_2078), .o(n_15932) );
na02f02 TIMEBOOST_cell_18646 ( .a(TIMEBOOST_net_5686), .b(n_8757), .o(g52401_db) );
no02f04 g74593_u0 ( .a(n_15939), .b(n_12716), .o(n_15940) );
in01f02 g74594_u0 ( .a(n_12924), .o(n_15939) );
no02f02 g74595_u0 ( .a(n_12717), .b(n_12461), .o(n_15941) );
na02f06 g74612_u0 ( .a(n_16334), .b(FE_OCP_RBN2227_g75174_p), .o(n_15969) );
ao12f10 g74627_u0 ( .a(n_1238), .b(n_15982), .c(n_15980), .o(n_15985) );
na02f10 g74628_u0 ( .a(n_15802), .b(wishbone_slave_unit_pci_initiator_if_write_req_int), .o(g74628_p) );
in01f08 g74628_u1 ( .a(g74628_p), .o(n_15980) );
in01f80 g74632_u0 ( .a(wishbone_slave_unit_pci_initiator_if_posted_write_req), .o(n_1238) );
in01f01 g74633_u0 ( .a(FE_OCPN1839_n_1238), .o(n_1041) );
in01f40 g74634_u0 ( .a(n_15981), .o(n_15988) );
in01f02 g74640_u0 ( .a(n_16290), .o(n_15994) );
na02f20 g74642_u0 ( .a(n_15996), .b(parchk_pci_cbe_reg_in_1236), .o(n_16326) );
in01m40 g74643_u0 ( .a(parchk_pci_cbe_reg_in_1237), .o(n_15996) );
no02f10 g74644_u0 ( .a(n_15744), .b(n_15924), .o(g74644_p) );
in01f10 g74644_u1 ( .a(g74644_p), .o(n_15999) );
no02f08 g74645_u0 ( .a(n_1291), .b(n_16289), .o(n_16002) );
in01f08 g74646_u0 ( .a(n_15998), .o(n_16003) );
na03f02 TIMEBOOST_cell_73479 ( .a(wbm_adr_o_4_), .b(g63203_sb), .c(g52450_sb), .o(TIMEBOOST_net_22955) );
na02f40 g74660_u0 ( .a(n_16942), .b(n_16635), .o(g74660_p) );
in01f20 g74660_u1 ( .a(g74660_p), .o(n_16016) );
na02f02 g74661_u0 ( .a(n_16914), .b(n_16021), .o(g74661_p) );
in01f02 g74661_u1 ( .a(g74661_p), .o(n_16022) );
in01f40 g74667_u0 ( .a(conf_w_addr_in_931), .o(n_16027) );
in01f08 g74668_u0 ( .a(n_16351), .o(n_16030) );
na02f40 g74673_u0 ( .a(n_629), .b(n_16284), .o(n_16033) );
in01f04 g74674_u0 ( .a(n_16034), .o(n_16036) );
no02f20 g74686_u0 ( .a(n_16048), .b(pci_target_unit_del_sync_bc_in_202), .o(n_16049) );
na02f40 g74687_u0 ( .a(n_16047), .b(pci_target_unit_del_sync_bc_in_201), .o(n_16048) );
in01f40 g74688_u0 ( .a(pci_target_unit_del_sync_bc_in_203), .o(n_16047) );
na02s01 g74689_u0 ( .a(FE_OFN2214_n_15366), .b(pci_target_unit_del_sync_bc_in_201), .o(g74689_p) );
no02f04 g74690_u0 ( .a(pci_target_unit_del_sync_bc_in_202), .b(pci_target_unit_del_sync_bc_in_203), .o(n_16052) );
na02f40 g74704_u0 ( .a(n_16066), .b(FE_OCPN1841_n_16089), .o(n_13221) );
in01f10 g74705_u0 ( .a(n_16486), .o(n_16066) );
in01f20 g74709_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_), .o(n_16070) );
no02f06 g74733_u0 ( .a(n_16573), .b(n_16577), .o(n_16105) );
no02f10 g74739_u0 ( .a(n_14981), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_), .o(g74739_p) );
in01f10 g74739_u1 ( .a(g74739_p), .o(n_16101) );
na02f10 g74740_u0 ( .a(n_14981), .b(n_16102), .o(n_16103) );
in01f20 g74741_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_), .o(n_16102) );
na02f10 g74749_u0 ( .a(n_16980), .b(n_16157), .o(g74749_p) );
in01s01 TIMEBOOST_cell_73862 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_), .o(TIMEBOOST_net_23427) );
no02f04 g74785_u0 ( .a(n_16152), .b(pci_target_unit_wbm_sm_pciw_fifo_control_in_86), .o(n_16153) );
na02f06 g74786_u0 ( .a(n_16150), .b(n_16151), .o(n_16152) );
na02f40 g74787_u0 ( .a(n_15385), .b(pci_target_unit_wishbone_master_rty_counter_6_), .o(g74787_p) );
in01f20 g74787_u1 ( .a(g74787_p), .o(n_16150) );
no03f80 g74788_u0 ( .a(n_705), .b(wbm_err_i), .c(wbm_ack_i), .o(n_16151) );
na02f02 TIMEBOOST_cell_4055 ( .a(TIMEBOOST_net_587), .b(n_3832), .o(n_4884) );
in01f20 g74793_u0 ( .a(n_1998), .o(n_16159) );
no02f40 g74794_u0 ( .a(n_819), .b(pci_target_unit_wishbone_master_c_state_2_), .o(n_16160) );
oa12f04 g74795_u0 ( .a(n_16160), .b(n_4642), .c(n_2387), .o(n_16162) );
ao12f04 g74796_u0 ( .a(n_16164), .b(n_2702), .c(n_4874), .o(n_16165) );
in01f02 g74797_u0 ( .a(n_16163), .o(n_16164) );
na02f10 g74798_u0 ( .a(n_16738), .b(n_16474), .o(n_16163) );
na02s02 TIMEBOOST_cell_42840 ( .a(TIMEBOOST_net_12314), .b(TIMEBOOST_net_8653), .o(n_9124) );
in01f08 g74800_u0 ( .a(n_16160), .o(n_16168) );
no02f02 g74802_u0 ( .a(n_14419), .b(n_16169), .o(n_16170) );
na04f04 TIMEBOOST_cell_24572 ( .a(n_9484), .b(g57472_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q), .d(FE_OFN2184_n_8567), .o(n_11262) );
in01f40 g74810_u0 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_), .o(n_16175) );
no02f08 g74818_u0 ( .a(n_16326), .b(n_16350), .o(n_16183) );
na03f06 g74828_u0 ( .a(n_16967), .b(n_16970), .c(n_16205), .o(n_16206) );
na02f02 g74838_u0 ( .a(n_16209), .b(n_16212), .o(n_16213) );
no02f02 g74839_u0 ( .a(n_16207), .b(n_16208), .o(n_16209) );
na02f02 TIMEBOOST_cell_71811 ( .a(TIMEBOOST_net_23113), .b(FE_OFN1770_n_14054), .o(n_14458) );
na04f04 TIMEBOOST_cell_24574 ( .a(n_9017), .b(g57485_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q), .d(FE_OFN2169_n_8567), .o(n_10332) );
no02f02 g74842_u0 ( .a(n_16210), .b(n_16211), .o(n_16212) );
na04f04 TIMEBOOST_cell_24318 ( .a(n_9655), .b(g57278_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q), .d(FE_OFN1425_n_8567), .o(n_11476) );
na02f02 g74850_u0 ( .a(n_16221), .b(n_16223), .o(n_16224) );
in01f02 g74851_u0 ( .a(n_16220), .o(n_16221) );
in01f02 g74853_u0 ( .a(n_16222), .o(n_16223) );
no02f02 g74856_u0 ( .a(n_16226), .b(n_16225), .o(n_16227) );
na02s01 g58354_u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q), .b(g58354_sb), .o(g58354_da) );
na04f04 TIMEBOOST_cell_24576 ( .a(n_9049), .b(g57367_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q), .d(FE_OFN2168_n_8567), .o(n_10383) );
na03m02 TIMEBOOST_cell_69984 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q), .b(FE_OFN2257_n_8060), .c(n_4522), .o(TIMEBOOST_net_22200) );
in01f02 g74859_u1 ( .a(g74859_p), .o(n_16228) );
in01f02 g74860_u0 ( .a(n_16229), .o(n_16230) );
na04f04 TIMEBOOST_cell_24578 ( .a(n_9572), .b(g57356_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q), .d(FE_OFN2190_n_8567), .o(n_11391) );
no02f02 g74866_u0 ( .a(n_16235), .b(n_16236), .o(n_16237) );
in01f02 g74867_u0 ( .a(n_13868), .o(n_16235) );
in01f02 g74868_u0 ( .a(n_14022), .o(n_16236) );
in01f02 g74869_u0 ( .a(n_16238), .o(n_16239) );
na04f04 TIMEBOOST_cell_24580 ( .a(n_9586), .b(g57341_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q), .d(FE_OFN2179_n_8567), .o(n_11410) );
na04m04 TIMEBOOST_cell_24582 ( .a(n_9129), .b(g57064_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q), .d(FE_OFN2167_n_8567), .o(n_10501) );
in01f02 g74872_u1 ( .a(g74872_p), .o(n_16241) );
no02f02 g74873_u0 ( .a(n_16242), .b(n_16243), .o(n_16244) );
na02f06 TIMEBOOST_cell_44993 ( .a(FE_OFN2069_n_15978), .b(wishbone_slave_unit_pcim_if_wbw_addr_data_in_400), .o(TIMEBOOST_net_13391) );
na04f04 TIMEBOOST_cell_24584 ( .a(n_8550), .b(g58606_sb), .c(n_251), .d(FE_OFN2182_n_8567), .o(n_8955) );
in01f02 g74879_u1 ( .a(g74879_p), .o(n_16248) );
no02f02 g74880_u0 ( .a(n_16249), .b(n_16250), .o(n_16251) );
na02m02 TIMEBOOST_cell_63943 ( .a(TIMEBOOST_net_20957), .b(FE_OFN1218_n_6886), .o(TIMEBOOST_net_15717) );
na04f04 TIMEBOOST_cell_24320 ( .a(n_9658), .b(g57276_sb), .c(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q), .d(FE_OFN1421_n_8567), .o(n_11478) );
in01f02 g74883_u0 ( .a(n_16252), .o(n_16253) );
na03f02 TIMEBOOST_cell_66410 ( .a(n_4723), .b(g63179_sb), .c(g63179_db), .o(n_7112) );
in01f02 g74886_u1 ( .a(g74886_p), .o(n_16255) );
no02f02 g74887_u0 ( .a(n_16256), .b(n_16257), .o(n_16258) );
na02s02 TIMEBOOST_cell_63227 ( .a(TIMEBOOST_net_20560), .b(FE_OFN233_n_9876), .o(TIMEBOOST_net_12818) );
na02f02 TIMEBOOST_cell_71437 ( .a(TIMEBOOST_net_22926), .b(n_15611), .o(n_14104) );
in01f02 g74890_u0 ( .a(n_16259), .o(n_16260) );
na02s01 TIMEBOOST_cell_43811 ( .a(FE_OFN211_n_9858), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q), .o(TIMEBOOST_net_12800) );
no02f10 g74892_u0 ( .a(n_16264), .b(n_16262), .o(n_16265) );
na02f40 g74893_u0 ( .a(n_15249), .b(pci_target_unit_wbm_sm_pci_tar_read_request), .o(n_16262) );
no02f80 g74894_u0 ( .a(FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_), .o(n_16264) );
in01f10 g74902_u0 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_), .o(n_16271) );
na03f02 TIMEBOOST_cell_35007 ( .a(TIMEBOOST_net_9575), .b(g57305_sb), .c(FE_OFN1370_n_8567), .o(n_11446) );
no02f80 g74907_u0 ( .a(pci_target_unit_pcit_if_strd_bc_in), .b(pci_target_unit_pcit_if_strd_bc_in_717), .o(n_16275) );
na03f02 TIMEBOOST_cell_53469 ( .a(n_1912), .b(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q), .c(FE_OFN2084_n_8407), .o(TIMEBOOST_net_16952) );
in01f80 g74916_u0 ( .a(conf_w_addr_in_937), .o(n_16284) );
in01f80 g74917_u0 ( .a(conf_w_addr_in_933), .o(n_16285) );
no02f10 g74920_u0 ( .a(n_16003), .b(n_15924), .o(g74920_p) );
in01f10 g74920_u1 ( .a(g74920_p), .o(n_16290) );
na02f10 g74921_u0 ( .a(n_16690), .b(conf_w_addr_in_938), .o(n_16291) );
na02f20 g74929_u0 ( .a(n_16293), .b(n_168), .o(n_13363) );
no02f08 g74930_u0 ( .a(n_14837), .b(n_12858), .o(g74930_p) );
in01f08 g74930_u1 ( .a(g74930_p), .o(n_16293) );
in01f10 g74932_u0 ( .a(n_16300), .o(n_16301) );
in01f08 g74933_u0 ( .a(n_16299), .o(n_16300) );
in01f01 g74935_u0 ( .a(n_16300), .o(n_16305) );
in01f10 g74936_u0 ( .a(n_13363), .o(n_16306) );
oa12f08 g74939_u0 ( .a(n_16354), .b(n_15958), .c(n_15960), .o(n_16309) );
na02f02 TIMEBOOST_cell_39663 ( .a(TIMEBOOST_net_11443), .b(g63109_sb), .o(n_5038) );
no02f08 g74961_u0 ( .a(n_2440), .b(FE_OFN996_n_15366), .o(g74961_p) );
in01f06 g74961_u1 ( .a(g74961_p), .o(n_16330) );
in01f04 g74962_u0 ( .a(n_16325), .o(n_16332) );
na02m02 TIMEBOOST_cell_30763 ( .a(n_9602), .b(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q), .o(TIMEBOOST_net_9486) );
na02f04 g74965_u0 ( .a(n_16334), .b(n_16364), .o(n_11767) );
na02f06 g74967_u0 ( .a(n_16550), .b(n_16368), .o(g74967_p) );
in01f06 g74967_u1 ( .a(g74967_p), .o(n_16334) );
na02f10 g74981_u0 ( .a(n_16351), .b(conf_w_addr_in), .o(g74981_p) );
in01f08 g74981_u1 ( .a(g74981_p), .o(n_16352) );
in01f80 g74983_u0 ( .a(parchk_pci_cbe_reg_in), .o(n_16350) );
in01f40 g74984_u0 ( .a(n_16354), .o(n_2071) );
in01f40 g74985_u0 ( .a(n_16350), .o(n_16354) );
na02f02 g74989_u0 ( .a(n_16474), .b(pci_target_unit_wbm_sm_pci_tar_burst_ok), .o(n_16358) );
no02f08 g74995_u0 ( .a(n_16076), .b(n_16444), .o(n_16364) );
na02f06 g74996_u0 ( .a(n_16368), .b(n_16554), .o(g74996_p) );
in01f06 g75021_u0 ( .a(n_16183), .o(n_16389) );
in01f40 g75022_u0 ( .a(conf_w_addr_in), .o(n_16390) );
na02f10 g75023_u0 ( .a(n_16352), .b(n_16388), .o(n_16392) );
in01f10 g75024_u0 ( .a(conf_w_addr_in), .o(g75024_sb) );
na02f02 g55236_u0 ( .a(FE_OCPN1827_n_14995), .b(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q), .o(n_12115) );
na02s01 TIMEBOOST_cell_30967 ( .a(wishbone_slave_unit_del_sync_addr_out_reg_19__Q), .b(FE_OFN264_n_9849), .o(TIMEBOOST_net_9588) );
no02f02 g75025_u0 ( .a(n_16398), .b(n_16400), .o(n_16401) );
in01f02 g75027_u0 ( .a(n_12600), .o(n_16395) );
no02f02 g75028_u0 ( .a(n_12597), .b(n_16396), .o(n_16397) );
in01f02 g75029_u0 ( .a(n_11887), .o(n_16396) );
in01f02 g75030_u0 ( .a(n_16399), .o(n_16400) );
no02f02 g75031_u0 ( .a(n_12599), .b(n_12598), .o(n_16399) );
na02s02 TIMEBOOST_cell_70257 ( .a(TIMEBOOST_net_22336), .b(FE_OFN542_n_9690), .o(TIMEBOOST_net_14942) );
in01f02 g75034_u0 ( .a(n_12754), .o(n_16402) );
in01f02 g75036_u0 ( .a(n_12752), .o(n_16404) );
no02f02 g75038_u0 ( .a(n_16412), .b(n_16408), .o(n_16413) );
na03f02 TIMEBOOST_cell_73131 ( .a(g64097_sb), .b(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q), .c(TIMEBOOST_net_14710), .o(TIMEBOOST_net_20466) );
in01m20 TIMEBOOST_cell_17843 ( .a(TIMEBOOST_net_5254), .o(n_2044) );
no02f02 g75041_u0 ( .a(n_12507), .b(n_12685), .o(n_16409) );
in01f02 g75042_u0 ( .a(n_12686), .o(n_16410) );
na02f01 g75054_u0 ( .a(n_16427), .b(n_16428), .o(n_16429) );
in01f06 g75056_u0 ( .a(n_16425), .o(n_16427) );
no02f20 g75058_u0 ( .a(n_16289), .b(n_16538), .o(n_16424) );
na02f40 g75059_u0 ( .a(pciu_am1_in_521), .b(pciu_bar1_in_383), .o(g75059_p) );
in01f20 g75059_u1 ( .a(g75059_p), .o(n_16428) );
na02f80 g75061_u0 ( .a(FE_OCP_RBN2269_pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_), .b(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_), .o(g75061_p) );
na02f10 g75066_u0 ( .a(n_16437), .b(n_16438), .o(n_16439) );
no02f40 g75067_u0 ( .a(n_16435), .b(n_16436), .o(g75067_p) );
in01f10 g75067_u1 ( .a(g75067_p), .o(n_16437) );
na02f80 g75069_u0 ( .a(n_7398), .b(n_6943), .o(n_16436) );
no02f08 g75071_u0 ( .a(n_16441), .b(n_16444), .o(n_16445) );
in01f06 g75072_u0 ( .a(n_16523), .o(g75072_sb) );
na02f08 g75072_u2 ( .a(n_16523), .b(n_16071), .o(g75072_db) );
na02m10 TIMEBOOST_cell_70096 ( .a(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_), .b(n_1293), .o(TIMEBOOST_net_22256) );
na02f10 g75073_u0 ( .a(n_16564), .b(n_16442), .o(n_16444) );
na03m02 TIMEBOOST_cell_65763 ( .a(TIMEBOOST_net_11075), .b(TIMEBOOST_net_8288), .c(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q), .o(TIMEBOOST_net_17405) );
na02f02 g59798_u2 ( .a(n_4688), .b(FE_OFN1700_n_5751), .o(g59798_db) );
in01f04 g75081_u1 ( .a(g75081_p), .o(n_16459) );
na03f02 TIMEBOOST_cell_73435 ( .a(TIMEBOOST_net_17458), .b(FE_OFN1293_n_4098), .c(g62667_sb), .o(n_6204) );
no02f08 g75083_u0 ( .a(n_1779), .b(wishbone_slave_unit_wishbone_slave_wb_conf_hit), .o(n_16451) );
na02f06 g75084_u0 ( .a(n_15014), .b(n_16021), .o(g75084_p) );
in01f08 g75084_u1 ( .a(g75084_p), .o(n_16452) );
no02f20 g75086_u0 ( .a(n_943), .b(wishbone_slave_unit_wishbone_slave_c_state_2), .o(n_14526) );
na02f06 g75088_u0 ( .a(n_7398), .b(n_6989), .o(g75088_p) );
in01f04 g75088_u1 ( .a(g75088_p), .o(n_16456) );
in01f20 g75090_u0 ( .a(n_14526), .o(n_16460) );
na02f40 g75114_u0 ( .a(n_16485), .b(n_16486), .o(n_16487) );
no02f20 g75115_u0 ( .a(n_15985), .b(n_15979), .o(n_16485) );
na02f40 g75117_u0 ( .a(n_1434), .b(n_1231), .o(n_16089) );
na02f10 g75119_u0 ( .a(n_16495), .b(n_16496), .o(n_16497) );
ao12f20 g75121_u0 ( .a(n_1539), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_), .o(n_16490) );
ao12f40 g75122_u0 ( .a(n_16491), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_), .o(n_16492) );
no02f80 g75123_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_), .o(n_16491) );
ao12f40 g75124_u0 ( .a(n_16493), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_), .c(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_), .o(n_16494) );
no02f80 g75125_u0 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_), .b(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_), .o(n_16493) );
na02f80 g75126_u0 ( .a(n_2597), .b(n_565), .o(g75126_p) );
in01f40 g75126_u1 ( .a(g75126_p), .o(n_16496) );
in01f08 g75131_u0 ( .a(n_16503), .o(n_16504) );
na02f08 g75138_u0 ( .a(n_16280), .b(pciu_cache_lsize_not_zero_in), .o(n_16507) );
in01s01 g75140_u0 ( .a(n_16507), .o(n_16512) );
in01f40 g75146_u0 ( .a(pci_target_unit_wishbone_master_retried), .o(n_16516) );
na02f10 g75147_u0 ( .a(n_16521), .b(FE_OCPN1823_n_16560), .o(n_16523) );
na02f08 g75148_u0 ( .a(n_16524), .b(n_16520), .o(n_16521) );
na02f10 g75151_u0 ( .a(n_15638), .b(FE_OCP_RBN2223_n_15347), .o(n_16524) );
no02f08 g75159_u0 ( .a(n_16533), .b(n_16534), .o(n_16535) );
in01f08 g75160_u0 ( .a(n_14981), .o(g75160_sb) );
na02m01 TIMEBOOST_cell_47947 ( .a(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q), .b(pci_target_unit_fifos_pcir_data_in_161), .o(TIMEBOOST_net_14191) );
na02f10 g75160_u2 ( .a(n_14981), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_), .o(g75160_db) );
in01f08 g75162_u0 ( .a(n_14981), .o(g75162_sb) );
na02f10 g75162_u2 ( .a(n_14981), .b(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_), .o(g75162_db) );
na02m04 TIMEBOOST_cell_54000 ( .a(TIMEBOOST_net_17217), .b(FE_OFN918_n_4725), .o(TIMEBOOST_net_14286) );
in01f08 g75163_u0 ( .a(n_16534), .o(n_16536) );
in01f10 g75164_u0 ( .a(n_16533), .o(n_16537) );
na02f08 g75165_u0 ( .a(n_16541), .b(n_16542), .o(g75165_p) );
in01f08 g75165_u1 ( .a(g75165_p), .o(n_16543) );
in01f06 g75166_u0 ( .a(n_16540), .o(n_16541) );
in01f08 g75168_u0 ( .a(FE_OCPN1852_n_16538), .o(n_16539) );
na02f40 g75169_u0 ( .a(n_16695), .b(conf_w_addr_in_938), .o(n_16538) );
no02f08 g75170_u0 ( .a(n_16290), .b(n_15744), .o(n_16542) );
na02f01 g75171_u0 ( .a(n_763), .b(n_1519), .o(n_16544) );
na02f04 g75173_u0 ( .a(n_16552), .b(FE_OCP_RBN2226_g75174_p), .o(n_16553) );
na02f06 g75174_u0 ( .a(n_16441), .b(n_16444), .o(g75174_p) );
na03f01 TIMEBOOST_cell_72415 ( .a(TIMEBOOST_net_13997), .b(wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q), .c(wbu_addr_in_270), .o(n_9844) );
na04f04 TIMEBOOST_cell_24803 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q), .b(g58834_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q), .d(FE_OFN2156_n_16439), .o(n_8603) );
na02f01 TIMEBOOST_cell_39457 ( .a(TIMEBOOST_net_11340), .b(FE_OFN1124_g64577_p), .o(n_5505) );
na04f04 TIMEBOOST_cell_24812 ( .a(wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q), .b(g58825_sb), .c(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q), .d(FE_OFN2153_n_16439), .o(n_8616) );
na04m06 TIMEBOOST_cell_72573 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q), .b(n_3739), .c(FE_OFN661_n_4392), .d(g64936_sb), .o(n_3677) );
na02f04 g75181_u2 ( .a(n_16273), .b(n_160), .o(g75181_db) );
na02f08 g75194_u0 ( .a(n_16566), .b(n_16579), .o(n_16572) );
no02f10 g75195_u0 ( .a(n_16536), .b(n_16537), .o(n_16566) );
na02f08 g75200_u0 ( .a(n_16573), .b(n_16578), .o(g75200_p) );
in01f08 g75200_u1 ( .a(g75200_p), .o(n_16579) );
na02f20 g75201_u0 ( .a(n_16101), .b(n_16103), .o(n_16573) );
na02f40 g75205_u0 ( .a(n_16487), .b(n_16089), .o(n_14981) );
in01f10 g75221_u0 ( .a(n_9256), .o(n_16637) );
in01f06 g75235_u0 ( .a(n_16690), .o(n_16685) );
in01f80 g75244_u0 ( .a(n_16695), .o(n_16690) );
in01f04 g75246_u0 ( .a(n_16695), .o(n_16696) );
in01f80 g75247_u0 ( .a(conf_w_addr_in_935), .o(n_16695) );
in01f08 g75259_u0 ( .a(n_8940), .o(n_16698) );
in01f10 g75272_u0 ( .a(FE_OCP_RBN2003_FE_OFN1026_n_16760), .o(n_16738) );
in01f08 g75277_u0 ( .a(n_16738), .o(TIMEBOOST_net_6736) );
in01f04 g75295_u0 ( .a(n_9170), .o(n_16779) );
in01s01 g75316_u0 ( .a(n_16818), .o(n_16816) );
na02f20 g75332_u0 ( .a(n_16952), .b(n_16635), .o(g75332_p) );
in01f20 g75332_u1 ( .a(g75332_p), .o(n_16854) );
in01f20 g75337_u0 ( .a(n_16864), .o(n_16860) );
in01f80 g75341_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_3_), .o(n_16864) );
in01f10 g75343_u0 ( .a(n_16871), .o(n_16867) );
in01f80 g75350_u0 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_2_), .o(n_16871) );
in01s01 g75351_u0 ( .a(n_16980), .o(n_16876) );
in01f06 g75362_u0 ( .a(n_16888), .o(n_16891) );
in01f10 g75365_u0 ( .a(n_16906), .o(n_16904) );
in01f80 g75367_u0 ( .a(pci_target_unit_wishbone_master_c_state_1_), .o(n_16906) );
in01f06 g75368_u0 ( .a(n_16910), .o(wbs_rty_o) );
in01f80 g75371_u0 ( .a(wbs_rty_o_1308), .o(n_16910) );
in01s01 g75372_u0 ( .a(n_16914), .o(n_16911) );
in01f40 g75386_u0 ( .a(n_16940), .o(n_16936) );
in01m08 g75393_u0 ( .a(FE_OCPN1832_n_16949), .o(n_16945) );
in01f20 g75399_u0 ( .a(n_16942), .o(n_16949) );
in01f80 g75400_u0 ( .a(n_16952), .o(n_16942) );
in01f80 g75401_u0 ( .a(wbu_we_in), .o(n_16952) );
na02f06 g75413_u2 ( .a(n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q), .o(g75413_db) );
na02f06 g75416_u2 ( .a(n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q), .o(g75416_db) );
na03s01 TIMEBOOST_cell_64713 ( .a(pci_target_unit_del_sync_addr_in_233), .b(g66415_sb), .c(g66420_db), .o(n_2510) );
na02f10 g75418_u1 ( .a(FE_OCP_RBN1956_n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q), .o(g75418_da) );
na02f08 g75418_u2 ( .a(n_16981), .b(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q), .o(g75418_db) );
na02f10 g75420_u0 ( .a(n_16131), .b(n_16980), .o(n_16981) );
na02f08 g75421_u0 ( .a(n_16976), .b(n_16977), .o(n_16131) );
no02f08 g75423_u0 ( .a(n_3421), .b(n_15117), .o(n_16977) );
na02f08 g75_u0 ( .a(n_8867), .b(n_16579), .o(g75_p) );
in01f08 g75_u1 ( .a(g75_p), .o(n_15558) );
in01s01 g78_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291), .o(n_15567) );
in01s01 g79_u0 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252), .o(n_15569) );
na02f80 g7_u0 ( .a(n_16635), .b(n_16818), .o(n_15371) );
no02f80 g9_u0 ( .a(n_16963), .b(FE_OCP_RBN1918_wbs_cti_i_1_), .o(n_16964) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_ack_o_reg_u0 ( .ck(ispd_clk), .d(n_10441), .o(wbs_ack_o_1307) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_0__u0 ( .ck(ispd_clk), .d(n_4106), .o(wbu_addr_in) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_10__u0 ( .ck(ispd_clk), .d(n_11876), .o(wbu_addr_in_259) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_11__u0 ( .ck(ispd_clk), .d(n_11878), .o(wbu_addr_in_260) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_12__u0 ( .ck(ispd_clk), .d(n_11875), .o(wbu_addr_in_261) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_13__u0 ( .ck(ispd_clk), .d(n_11874), .o(wbu_addr_in_262) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_14__u0 ( .ck(ispd_clk), .d(n_11872), .o(wbu_addr_in_263) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_15__u0 ( .ck(ispd_clk), .d(n_11873), .o(wbu_addr_in_264) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_16__u0 ( .ck(ispd_clk), .d(n_11871), .o(wbu_addr_in_265) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_17__u0 ( .ck(ispd_clk), .d(n_11870), .o(wbu_addr_in_266) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_18__u0 ( .ck(ispd_clk), .d(n_11869), .o(wbu_addr_in_267) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_19__u0 ( .ck(ispd_clk), .d(n_11868), .o(wbu_addr_in_268) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_1__u0 ( .ck(ispd_clk), .d(n_4105), .o(wbu_addr_in_250) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_20__u0 ( .ck(ispd_clk), .d(n_11867), .o(wbu_addr_in_269) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_21__u0 ( .ck(ispd_clk), .d(n_11866), .o(wbu_addr_in_270) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_22__u0 ( .ck(ispd_clk), .d(n_11865), .o(wbu_addr_in_271) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_23__u0 ( .ck(ispd_clk), .d(n_11864), .o(wbu_addr_in_272) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_24__u0 ( .ck(ispd_clk), .d(n_11863), .o(wbu_addr_in_273) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_25__u0 ( .ck(ispd_clk), .d(n_11862), .o(wbu_addr_in_274) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_26__u0 ( .ck(ispd_clk), .d(n_11861), .o(wbu_addr_in_275) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_27__u0 ( .ck(ispd_clk), .d(n_11860), .o(wbu_addr_in_276) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_28__u0 ( .ck(ispd_clk), .d(n_11859), .o(wbu_addr_in_277) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23400), .o(i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__Q) );
in01f40 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__u1 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_29__Q), .o(wbu_addr_in_278) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_2__u0 ( .ck(ispd_clk), .d(n_11858), .o(wbu_addr_in_251) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_30__u0 ( .ck(ispd_clk), .d(n_11857), .o(wbu_addr_in_279) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23402), .o(i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__Q) );
in01f40 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__u1 ( .a(i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_31__Q), .o(wbu_addr_in_280) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_3__u0 ( .ck(ispd_clk), .d(n_11854), .o(wbu_addr_in_252) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_4__u0 ( .ck(ispd_clk), .d(n_11853), .o(wbu_addr_in_253) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_5__u0 ( .ck(ispd_clk), .d(n_11852), .o(wbu_addr_in_254) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_6__u0 ( .ck(ispd_clk), .d(n_11851), .o(wbu_addr_in_255) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_7__u0 ( .ck(ispd_clk), .d(n_11850), .o(wbu_addr_in_256) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_8__u0 ( .ck(ispd_clk), .d(n_11848), .o(wbu_addr_in_257) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_adr_o_reg_9__u0 ( .ck(ispd_clk), .d(n_11849), .o(wbu_addr_in_258) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_cab_o_reg_u0 ( .ck(ispd_clk), .d(n_5723), .o(n_16818) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_cyc_o_reg_u0 ( .ck(ispd_clk), .d(n_12169), .o(n_16635) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__u0 ( .ck(ispd_clk), .d(n_7147), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_0__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__u0 ( .ck(ispd_clk), .d(n_7145), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_10__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__u0 ( .ck(ispd_clk), .d(n_7193), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_11__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__u0 ( .ck(ispd_clk), .d(n_7191), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_12__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__u0 ( .ck(ispd_clk), .d(n_7189), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_13__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__u0 ( .ck(ispd_clk), .d(n_7143), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_14__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__u0 ( .ck(ispd_clk), .d(n_7151), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_15__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__u0 ( .ck(ispd_clk), .d(n_7177), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_16__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__u0 ( .ck(ispd_clk), .d(n_7187), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_17__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__u0 ( .ck(ispd_clk), .d(n_7149), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_18__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__u0 ( .ck(ispd_clk), .d(n_7157), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_19__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__u0 ( .ck(ispd_clk), .d(n_7197), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_1__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__u0 ( .ck(ispd_clk), .d(n_7141), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_20__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__u0 ( .ck(ispd_clk), .d(n_7185), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_21__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__u0 ( .ck(ispd_clk), .d(n_7139), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_22__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__u0 ( .ck(ispd_clk), .d(n_7195), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_23__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__u0 ( .ck(ispd_clk), .d(n_7182), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_24__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__u0 ( .ck(ispd_clk), .d(n_7203), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_25__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__u0 ( .ck(ispd_clk), .d(n_7205), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_26__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__u0 ( .ck(ispd_clk), .d(n_7180), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_27__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__u0 ( .ck(ispd_clk), .d(n_7207), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_28__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__u0 ( .ck(ispd_clk), .d(n_7174), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_29__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__u0 ( .ck(ispd_clk), .d(n_7171), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_2__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__u0 ( .ck(ispd_clk), .d(n_7168), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_30__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__u0 ( .ck(ispd_clk), .d(n_7165), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_31__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__u0 ( .ck(ispd_clk), .d(n_7163), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_3__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__u0 ( .ck(ispd_clk), .d(n_7161), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_4__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__u0 ( .ck(ispd_clk), .d(n_7159), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_5__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__u0 ( .ck(ispd_clk), .d(n_7209), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_6__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__u0 ( .ck(ispd_clk), .d(n_7155), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_7__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__u0 ( .ck(ispd_clk), .d(n_7200), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_8__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__u0 ( .ck(ispd_clk), .d(n_7153), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_reg_9__Q) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid_reg_u0 ( .ck(ispd_clk), .d(n_11844), .o(i_pci_wbs_wbb3_2_wbb2_wbs_dat_i_o_valid) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_0__u0 ( .ck(ispd_clk), .d(n_13727), .o(wbs_dat_o_0_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_10__u0 ( .ck(ispd_clk), .d(n_13823), .o(wbs_dat_o_10_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_11__u0 ( .ck(ispd_clk), .d(n_13822), .o(wbs_dat_o_11_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_12__u0 ( .ck(ispd_clk), .d(n_13724), .o(wbs_dat_o_12_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_13__u0 ( .ck(ispd_clk), .d(n_13719), .o(wbs_dat_o_13_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_14__u0 ( .ck(ispd_clk), .d(n_13717), .o(wbs_dat_o_14_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_15__u0 ( .ck(ispd_clk), .d(n_13744), .o(wbs_dat_o_15_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_16__u0 ( .ck(ispd_clk), .d(n_13816), .o(wbs_dat_o_16_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_17__u0 ( .ck(ispd_clk), .d(n_13712), .o(wbs_dat_o_17_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_18__u0 ( .ck(ispd_clk), .d(n_13815), .o(wbs_dat_o_18_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_19__u0 ( .ck(ispd_clk), .d(n_13812), .o(wbs_dat_o_19_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_1__u0 ( .ck(ispd_clk), .d(n_13809), .o(wbs_dat_o_1_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_20__u0 ( .ck(ispd_clk), .d(n_13709), .o(wbs_dat_o_20_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_21__u0 ( .ck(ispd_clk), .d(n_13806), .o(wbs_dat_o_21_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_22__u0 ( .ck(ispd_clk), .d(n_13798), .o(wbs_dat_o_22_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_23__u0 ( .ck(ispd_clk), .d(n_13705), .o(wbs_dat_o_23_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_24__u0 ( .ck(ispd_clk), .d(n_13740), .o(wbs_dat_o_24_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_25__u0 ( .ck(ispd_clk), .d(n_13738), .o(wbs_dat_o_25_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_26__u0 ( .ck(ispd_clk), .d(n_13698), .o(wbs_dat_o_26_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_27__u0 ( .ck(ispd_clk), .d(n_13735), .o(wbs_dat_o_27_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_28__u0 ( .ck(ispd_clk), .d(n_13697), .o(wbs_dat_o_28_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_29__u0 ( .ck(ispd_clk), .d(n_13696), .o(wbs_dat_o_29_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_2__u0 ( .ck(ispd_clk), .d(n_13734), .o(wbs_dat_o_2_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_30__u0 ( .ck(ispd_clk), .d(n_13794), .o(wbs_dat_o_30_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_31__u0 ( .ck(ispd_clk), .d(n_13694), .o(wbs_dat_o_31_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_3__u0 ( .ck(ispd_clk), .d(n_13693), .o(wbs_dat_o_3_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_4__u0 ( .ck(ispd_clk), .d(n_13688), .o(wbs_dat_o_4_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_5__u0 ( .ck(ispd_clk), .d(n_13793), .o(wbs_dat_o_5_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_6__u0 ( .ck(ispd_clk), .d(n_13792), .o(wbs_dat_o_6_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_7__u0 ( .ck(ispd_clk), .d(n_13687), .o(wbs_dat_o_7_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_8__u0 ( .ck(ispd_clk), .d(n_13686), .o(wbs_dat_o_8_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_dat_o_o_reg_9__u0 ( .ck(ispd_clk), .d(n_13685), .o(wbs_dat_o_9_) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_err_o_reg_u0 ( .ck(ispd_clk), .d(n_8874), .o(wbs_err_o_1309) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_rty_o_reg_u0 ( .ck(ispd_clk), .d(n_8583), .o(wbs_rty_o_1308) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg_0__u0 ( .ck(ispd_clk), .d(n_4104), .o(wbu_sel_in) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg_1__u0 ( .ck(ispd_clk), .d(n_4103), .o(wbu_sel_in_312) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg_2__u0 ( .ck(ispd_clk), .d(n_4102), .o(wbu_sel_in_313) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_sel_o_reg_3__u0 ( .ck(ispd_clk), .d(n_4101), .o(wbu_sel_in_314) );
ms00f80 i_pci_wbs_wbb3_2_wbb2_wbs_we_o_reg_u0 ( .ck(ispd_clk), .d(n_4100), .o(wbu_we_in) );
ms00f80 input_register_pci_ad_reg_out_reg_0__u0 ( .ck(ispd_clk), .d(n_1654), .o(parchk_pci_ad_reg_in) );
ms00f80 input_register_pci_ad_reg_out_reg_10__u0 ( .ck(ispd_clk), .d(n_1497), .o(parchk_pci_ad_reg_in_1214) );
ms00f80 input_register_pci_ad_reg_out_reg_11__u0 ( .ck(ispd_clk), .d(n_1429), .o(parchk_pci_ad_reg_in_1215) );
ms00f80 input_register_pci_ad_reg_out_reg_12__u0 ( .ck(ispd_clk), .d(n_1647), .o(parchk_pci_ad_reg_in_1216) );
ms00f80 input_register_pci_ad_reg_out_reg_13__u0 ( .ck(ispd_clk), .d(n_1685), .o(parchk_pci_ad_reg_in_1217) );
ms00f80 input_register_pci_ad_reg_out_reg_14__u0 ( .ck(ispd_clk), .d(n_1502), .o(parchk_pci_ad_reg_in_1218) );
ms00f80 input_register_pci_ad_reg_out_reg_15__u0 ( .ck(ispd_clk), .d(n_1634), .o(parchk_pci_ad_reg_in_1219) );
ms00f80 input_register_pci_ad_reg_out_reg_16__u0 ( .ck(ispd_clk), .d(n_1499), .o(parchk_pci_ad_reg_in_1220) );
ms00f80 input_register_pci_ad_reg_out_reg_17__u0 ( .ck(ispd_clk), .d(n_1652), .o(parchk_pci_ad_reg_in_1221) );
ms00f80 input_register_pci_ad_reg_out_reg_18__u0 ( .ck(ispd_clk), .d(n_1428), .o(parchk_pci_ad_reg_in_1222) );
ms00f80 input_register_pci_ad_reg_out_reg_19__u0 ( .ck(ispd_clk), .d(n_1274), .o(parchk_pci_ad_reg_in_1223) );
ms00f80 input_register_pci_ad_reg_out_reg_1__u0 ( .ck(ispd_clk), .d(n_1272), .o(parchk_pci_ad_reg_in_1205) );
ms00f80 input_register_pci_ad_reg_out_reg_20__u0 ( .ck(ispd_clk), .d(n_1495), .o(parchk_pci_ad_reg_in_1224) );
ms00f80 input_register_pci_ad_reg_out_reg_21__u0 ( .ck(ispd_clk), .d(n_1431), .o(parchk_pci_ad_reg_in_1225) );
ms00f80 input_register_pci_ad_reg_out_reg_22__u0 ( .ck(ispd_clk), .d(n_1474), .o(parchk_pci_ad_reg_in_1226) );
ms00f80 input_register_pci_ad_reg_out_reg_23__u0 ( .ck(ispd_clk), .d(n_1681), .o(parchk_pci_ad_reg_in_1227) );
ms00f80 input_register_pci_ad_reg_out_reg_24__u0 ( .ck(ispd_clk), .d(n_1503), .o(parchk_pci_ad_reg_in_1228) );
ms00f80 input_register_pci_ad_reg_out_reg_25__u0 ( .ck(ispd_clk), .d(n_1704), .o(parchk_pci_ad_reg_in_1229) );
ms00f80 input_register_pci_ad_reg_out_reg_26__u0 ( .ck(ispd_clk), .d(n_1444), .o(parchk_pci_ad_reg_in_1230) );
ms00f80 input_register_pci_ad_reg_out_reg_27__u0 ( .ck(ispd_clk), .d(n_1483), .o(parchk_pci_ad_reg_in_1231) );
ms00f80 input_register_pci_ad_reg_out_reg_28__u0 ( .ck(ispd_clk), .d(n_1501), .o(parchk_pci_ad_reg_in_1232) );
ms00f80 input_register_pci_ad_reg_out_reg_29__u0 ( .ck(ispd_clk), .d(n_1677), .o(parchk_pci_ad_reg_in_1233) );
ms00f80 input_register_pci_ad_reg_out_reg_2__u0 ( .ck(ispd_clk), .d(n_1277), .o(parchk_pci_ad_reg_in_1206) );
ms00f80 input_register_pci_ad_reg_out_reg_30__u0 ( .ck(ispd_clk), .d(n_1640), .o(n_2509) );
ms00f80 input_register_pci_ad_reg_out_reg_31__u0 ( .ck(ispd_clk), .d(n_1470), .o(parchk_pci_ad_reg_in_1235) );
ms00f80 input_register_pci_ad_reg_out_reg_3__u0 ( .ck(ispd_clk), .d(n_1649), .o(parchk_pci_ad_reg_in_1207) );
ms00f80 input_register_pci_ad_reg_out_reg_4__u0 ( .ck(ispd_clk), .d(n_1683), .o(parchk_pci_ad_reg_in_1208) );
ms00f80 input_register_pci_ad_reg_out_reg_5__u0 ( .ck(ispd_clk), .d(n_1411), .o(parchk_pci_ad_reg_in_1209) );
ms00f80 input_register_pci_ad_reg_out_reg_6__u0 ( .ck(ispd_clk), .d(n_1276), .o(parchk_pci_ad_reg_in_1210) );
ms00f80 input_register_pci_ad_reg_out_reg_7__u0 ( .ck(ispd_clk), .d(n_1614), .o(parchk_pci_ad_reg_in_1211) );
ms00f80 input_register_pci_ad_reg_out_reg_8__u0 ( .ck(ispd_clk), .d(n_1275), .o(parchk_pci_ad_reg_in_1212) );
ms00f80 input_register_pci_ad_reg_out_reg_9__u0 ( .ck(ispd_clk), .d(n_1641), .o(parchk_pci_ad_reg_in_1213) );
ms00f80 input_register_pci_cbe_reg_out_reg_0__u0 ( .ck(ispd_clk), .d(n_3118), .o(parchk_pci_cbe_reg_in) );
ms00f80 input_register_pci_cbe_reg_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2564), .o(parchk_pci_cbe_reg_in_1236) );
ms00f80 input_register_pci_cbe_reg_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2568), .o(parchk_pci_cbe_reg_in_1237) );
ms00f80 input_register_pci_cbe_reg_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2567), .o(parchk_pci_cbe_reg_in_1238) );
ms00f80 input_register_pci_devsel_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2374), .o(wbu_pciif_devsel_reg_in) );
ms00f80 input_register_pci_frame_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2372), .o(parchk_pci_frame_reg_in) );
ms00f80 input_register_pci_idsel_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_1452), .o(pciu_pciif_idsel_reg_in) );
ms00f80 input_register_pci_irdy_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2471), .o(n_657) );
ms00f80 input_register_pci_stop_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2147), .o(pciu_pciif_stop_reg_in) );
ms00f80 input_register_pci_trdy_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_2718), .o(parchk_pci_trdy_reg_in) );
ms00f80 output_backup_ad_out_reg_0__u0 ( .ck(ispd_clk), .d(n_13908), .o(parchk_pci_ad_out_in) );
ms00f80 output_backup_ad_out_reg_10__u0 ( .ck(ispd_clk), .d(n_14320), .o(parchk_pci_ad_out_in_1177) );
ms00f80 output_backup_ad_out_reg_11__u0 ( .ck(ispd_clk), .d(n_14316), .o(parchk_pci_ad_out_in_1178) );
ms00f80 output_backup_ad_out_reg_12__u0 ( .ck(ispd_clk), .d(n_14318), .o(parchk_pci_ad_out_in_1179) );
ms00f80 output_backup_ad_out_reg_13__u0 ( .ck(ispd_clk), .d(n_14314), .o(parchk_pci_ad_out_in_1180) );
ms00f80 output_backup_ad_out_reg_14__u0 ( .ck(ispd_clk), .d(n_14312), .o(parchk_pci_ad_out_in_1181) );
ms00f80 output_backup_ad_out_reg_15__u0 ( .ck(ispd_clk), .d(n_14310), .o(parchk_pci_ad_out_in_1182) );
ms00f80 output_backup_ad_out_reg_16__u0 ( .ck(ispd_clk), .d(n_14383), .o(parchk_pci_ad_out_in_1183) );
ms00f80 output_backup_ad_out_reg_17__u0 ( .ck(ispd_clk), .d(n_14382), .o(parchk_pci_ad_out_in_1184) );
ms00f80 output_backup_ad_out_reg_18__u0 ( .ck(ispd_clk), .d(n_14381), .o(parchk_pci_ad_out_in_1185) );
ms00f80 output_backup_ad_out_reg_19__u0 ( .ck(ispd_clk), .d(n_14380), .o(parchk_pci_ad_out_in_1186) );
ms00f80 output_backup_ad_out_reg_1__u0 ( .ck(ispd_clk), .d(n_14094), .o(parchk_pci_ad_out_in_1168) );
ms00f80 output_backup_ad_out_reg_20__u0 ( .ck(ispd_clk), .d(n_14379), .o(parchk_pci_ad_out_in_1187) );
ms00f80 output_backup_ad_out_reg_21__u0 ( .ck(ispd_clk), .d(n_14093), .o(parchk_pci_ad_out_in_1188) );
ms00f80 output_backup_ad_out_reg_22__u0 ( .ck(ispd_clk), .d(n_14378), .o(parchk_pci_ad_out_in_1189) );
ms00f80 output_backup_ad_out_reg_23__u0 ( .ck(ispd_clk), .d(n_14377), .o(parchk_pci_ad_out_in_1190) );
ms00f80 output_backup_ad_out_reg_24__u0 ( .ck(ispd_clk), .d(n_14376), .o(parchk_pci_ad_out_in_1191) );
ms00f80 output_backup_ad_out_reg_25__u0 ( .ck(ispd_clk), .d(n_13831), .o(parchk_pci_ad_out_in_1192) );
ms00f80 output_backup_ad_out_reg_26__u0 ( .ck(ispd_clk), .d(n_14078), .o(parchk_pci_ad_out_in_1193) );
ms00f80 output_backup_ad_out_reg_27__u0 ( .ck(ispd_clk), .d(n_14375), .o(parchk_pci_ad_out_in_1194) );
ms00f80 output_backup_ad_out_reg_28__u0 ( .ck(ispd_clk), .d(n_14374), .o(parchk_pci_ad_out_in_1195) );
ms00f80 output_backup_ad_out_reg_29__u0 ( .ck(ispd_clk), .d(n_14373), .o(parchk_pci_ad_out_in_1196) );
ms00f80 output_backup_ad_out_reg_2__u0 ( .ck(ispd_clk), .d(n_14372), .o(parchk_pci_ad_out_in_1169) );
ms00f80 output_backup_ad_out_reg_30__u0 ( .ck(ispd_clk), .d(n_14088), .o(parchk_pci_ad_out_in_1197) );
ms00f80 output_backup_ad_out_reg_31__u0 ( .ck(ispd_clk), .d(n_14531), .o(parchk_pci_ad_out_in_1198) );
ms00f80 output_backup_ad_out_reg_3__u0 ( .ck(ispd_clk), .d(n_14371), .o(parchk_pci_ad_out_in_1170) );
ms00f80 output_backup_ad_out_reg_4__u0 ( .ck(ispd_clk), .d(n_14370), .o(parchk_pci_ad_out_in_1171) );
ms00f80 output_backup_ad_out_reg_5__u0 ( .ck(ispd_clk), .d(n_14369), .o(parchk_pci_ad_out_in_1172) );
ms00f80 output_backup_ad_out_reg_6__u0 ( .ck(ispd_clk), .d(n_14368), .o(parchk_pci_ad_out_in_1173) );
ms00f80 output_backup_ad_out_reg_7__u0 ( .ck(ispd_clk), .d(n_14367), .o(parchk_pci_ad_out_in_1174) );
ms00f80 output_backup_ad_out_reg_8__u0 ( .ck(ispd_clk), .d(n_14366), .o(parchk_pci_ad_out_in_1175) );
ms00f80 output_backup_ad_out_reg_9__u0 ( .ck(ispd_clk), .d(n_14365), .o(parchk_pci_ad_out_in_1176) );
ms00f80 output_backup_cbe_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7135), .o(parchk_pci_cbe_en_in) );
ms00f80 output_backup_cbe_out_reg_0__u0 ( .ck(ispd_clk), .d(n_14397), .o(parchk_pci_cbe_out_in) );
ms00f80 output_backup_cbe_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23404), .o(parchk_pci_cbe_out_in_1202) );
ms00f80 output_backup_cbe_out_reg_2__u0 ( .ck(ispd_clk), .d(n_14396), .o(parchk_pci_cbe_out_in_1203) );
ms00f80 output_backup_cbe_out_reg_3__u0 ( .ck(ispd_clk), .d(n_14394), .o(parchk_pci_cbe_out_in_1204) );
ms00f80 output_backup_devsel_out_reg_u0 ( .ck(ispd_clk), .d(n_14616), .o(output_backup_devsel_out_reg_Q) );
ms00f80 output_backup_frame_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7210), .o(parchk_pci_frame_en_in) );
ms00f80 output_backup_frame_out_reg_u0 ( .ck(ispd_clk), .d(n_8752), .o(wbu_pciif_frame_out_in) );
ms00f80 output_backup_irdy_en_out_reg_u0 ( .ck(ispd_clk), .d(n_447), .o(parchk_pci_irdy_en_in) );
ms00f80 output_backup_irdy_out_reg_u0 ( .ck(ispd_clk), .d(n_2900), .o(out_bckp_irdy_out) );
ms00f80 output_backup_mas_ad_en_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23406), .o(n_14905) );
ms00f80 output_backup_par_en_out_reg_u0 ( .ck(ispd_clk), .d(n_12954), .o(output_backup_par_en_out_reg_Q) );
in01m80 output_backup_par_en_out_reg_u1 ( .a(output_backup_par_en_out_reg_Q), .o(parchk_pci_par_en_in) );
ms00f80 output_backup_par_out_reg_u0 ( .ck(ispd_clk), .d(n_8576), .o(output_backup_par_out_reg_Q) );
ms00f80 output_backup_perr_en_out_reg_u0 ( .ck(ispd_clk), .d(n_14572), .o(out_bckp_perr_en_out) );
ms00f80 output_backup_perr_out_reg_u0 ( .ck(ispd_clk), .d(n_13918), .o(output_backup_perr_out_reg_Q) );
in01s01 output_backup_perr_out_reg_u1 ( .a(output_backup_perr_out_reg_Q), .o(parchk_pci_perr_out_in) );
ms00f80 output_backup_serr_en_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23408), .o(output_backup_serr_en_out_reg_Q) );
in01s01 output_backup_serr_en_out_reg_u1 ( .a(output_backup_serr_en_out_reg_Q), .o(parchk_pci_serr_en_in) );
ms00f80 output_backup_serr_out_reg_u0 ( .ck(ispd_clk), .d(n_13917), .o(parchk_pci_serr_out_in) );
ms00f80 output_backup_stop_out_reg_u0 ( .ck(ispd_clk), .d(n_14617), .o(output_backup_stop_out_reg_Q) );
in01f40 output_backup_stop_out_reg_u1 ( .a(output_backup_stop_out_reg_Q), .o(pciu_pciif_bckp_stop_in) );
ms00f80 output_backup_tar_ad_en_out_reg_u0 ( .ck(ispd_clk), .d(n_11448), .o(output_backup_tar_ad_en_out_reg_Q) );
in01f80 output_backup_tar_ad_en_out_reg_u1 ( .a(output_backup_tar_ad_en_out_reg_Q), .o(n_13784) );
ms00f80 output_backup_trdy_en_out_reg_u0 ( .ck(ispd_clk), .d(n_8875), .o(parchk_pci_trdy_en_in) );
ms00f80 output_backup_trdy_out_reg_u0 ( .ck(ispd_clk), .d(n_14622), .o(output_backup_trdy_out_reg_Q) );
ms00f80 parity_checker_check_for_serr_on_second_reg_u0 ( .ck(ispd_clk), .d(n_3794), .o(parity_checker_check_for_serr_on_second_reg_Q) );
in01m08 parity_checker_check_for_serr_on_second_reg_u1 ( .a(parity_checker_check_for_serr_on_second_reg_Q), .o(parity_checker_check_for_serr_on_second) );
ms00f80 parity_checker_check_perr_reg_u0 ( .ck(ispd_clk), .d(g54038_sb), .o(parity_checker_check_perr_reg_Q) );
in01s01 parity_checker_check_perr_reg_u1 ( .a(parity_checker_check_perr_reg_Q), .o(parity_checker_check_perr) );
ms00f80 parity_checker_frame_and_irdy_en_prev_prev_reg_u0 ( .ck(ispd_clk), .d(parity_checker_frame_and_irdy_en_prev), .o(parity_checker_frame_and_irdy_en_prev_prev) );
ms00f80 parity_checker_frame_and_irdy_en_prev_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23410), .o(parity_checker_frame_and_irdy_en_prev) );
ms00f80 parity_checker_frame_dec2_reg_u0 ( .ck(ispd_clk), .d(n_15302), .o(parity_checker_frame_dec2) );
ms00f80 parity_checker_master_perr_report_reg_u0 ( .ck(ispd_clk), .d(parity_checker_frame_and_irdy_en_prev_prev), .o(parity_checker_master_perr_report_reg_Q) );
in01s01 parity_checker_master_perr_report_reg_u1 ( .a(parity_checker_master_perr_report_reg_Q), .o(parity_checker_master_perr_report) );
ms00f80 parity_checker_perr_en_crit_gen_perr_en_reg_out_reg_u0 ( .ck(ispd_clk), .d(n_14386), .o(parity_checker_pci_perr_en_reg) );
ms00f80 parity_checker_perr_sampled_reg_u0 ( .ck(ispd_clk), .d(n_14765), .o(parity_checker_perr_sampled) );
ms00f80 pci_io_mux_ad_iob0_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_13911), .o(pci_ad_o_0_) );
ms00f80 pci_io_mux_ad_iob0_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_0_) );
ms00f80 pci_io_mux_ad_iob10_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14364), .o(pci_ad_o_10_) );
ms00f80 pci_io_mux_ad_iob10_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_10_) );
ms00f80 pci_io_mux_ad_iob11_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14363), .o(pci_ad_o_11_) );
ms00f80 pci_io_mux_ad_iob11_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_11_) );
ms00f80 pci_io_mux_ad_iob12_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14362), .o(pci_ad_o_12_) );
ms00f80 pci_io_mux_ad_iob12_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_12_) );
ms00f80 pci_io_mux_ad_iob13_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14361), .o(pci_ad_o_13_) );
ms00f80 pci_io_mux_ad_iob13_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_13_) );
ms00f80 pci_io_mux_ad_iob14_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14360), .o(pci_ad_o_14_) );
ms00f80 pci_io_mux_ad_iob14_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_14_) );
ms00f80 pci_io_mux_ad_iob15_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14359), .o(pci_ad_o_15_) );
ms00f80 pci_io_mux_ad_iob15_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_15_) );
ms00f80 pci_io_mux_ad_iob16_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14358), .o(pci_ad_o_16_) );
ms00f80 pci_io_mux_ad_iob16_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_16_) );
ms00f80 pci_io_mux_ad_iob17_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14356), .o(pci_ad_o_17_) );
ms00f80 pci_io_mux_ad_iob17_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_17_) );
ms00f80 pci_io_mux_ad_iob18_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14354), .o(pci_ad_o_18_) );
ms00f80 pci_io_mux_ad_iob18_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_18_) );
ms00f80 pci_io_mux_ad_iob19_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14352), .o(pci_ad_o_19_) );
ms00f80 pci_io_mux_ad_iob19_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_19_) );
ms00f80 pci_io_mux_ad_iob1_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14086), .o(pci_ad_o_1_) );
ms00f80 pci_io_mux_ad_iob1_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_1_) );
ms00f80 pci_io_mux_ad_iob20_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14350), .o(pci_ad_o_20_) );
ms00f80 pci_io_mux_ad_iob20_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_20_) );
ms00f80 pci_io_mux_ad_iob21_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14084), .o(pci_ad_o_21_) );
ms00f80 pci_io_mux_ad_iob21_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_21_) );
ms00f80 pci_io_mux_ad_iob22_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14348), .o(pci_ad_o_22_) );
ms00f80 pci_io_mux_ad_iob22_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_22_) );
ms00f80 pci_io_mux_ad_iob23_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14342), .o(pci_ad_o_23_) );
ms00f80 pci_io_mux_ad_iob23_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_23_) );
ms00f80 pci_io_mux_ad_iob24_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14346), .o(pci_ad_o_24_) );
ms00f80 pci_io_mux_ad_iob24_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_24_) );
ms00f80 pci_io_mux_ad_iob25_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_13830), .o(pci_ad_o_25_) );
ms00f80 pci_io_mux_ad_iob25_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_25_) );
ms00f80 pci_io_mux_ad_iob26_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14077), .o(pci_ad_o_26_) );
ms00f80 pci_io_mux_ad_iob26_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_26_) );
ms00f80 pci_io_mux_ad_iob27_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14344), .o(pci_ad_o_27_) );
ms00f80 pci_io_mux_ad_iob27_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_27_) );
ms00f80 pci_io_mux_ad_iob28_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14338), .o(pci_ad_o_28_) );
ms00f80 pci_io_mux_ad_iob28_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_28_) );
ms00f80 pci_io_mux_ad_iob29_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14340), .o(pci_ad_o_29_) );
ms00f80 pci_io_mux_ad_iob29_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_29_) );
ms00f80 pci_io_mux_ad_iob2_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14336), .o(pci_ad_o_2_) );
ms00f80 pci_io_mux_ad_iob2_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_2_) );
ms00f80 pci_io_mux_ad_iob30_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14082), .o(pci_ad_o_30_) );
ms00f80 pci_io_mux_ad_iob30_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1506_n_15768), .o(pci_ad_oe_o_30_) );
ms00f80 pci_io_mux_ad_iob31_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14530), .o(pci_ad_o_31_) );
ms00f80 pci_io_mux_ad_iob31_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_31_) );
ms00f80 pci_io_mux_ad_iob3_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14334), .o(pci_ad_o_3_) );
ms00f80 pci_io_mux_ad_iob3_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_3_) );
ms00f80 pci_io_mux_ad_iob4_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14332), .o(pci_ad_o_4_) );
ms00f80 pci_io_mux_ad_iob4_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_4_) );
ms00f80 pci_io_mux_ad_iob5_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14330), .o(pci_ad_o_5_) );
ms00f80 pci_io_mux_ad_iob5_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_5_) );
ms00f80 pci_io_mux_ad_iob6_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14328), .o(pci_ad_o_6_) );
ms00f80 pci_io_mux_ad_iob6_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_6_) );
ms00f80 pci_io_mux_ad_iob7_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14326), .o(pci_ad_o_7_) );
ms00f80 pci_io_mux_ad_iob7_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_7_) );
ms00f80 pci_io_mux_ad_iob8_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14324), .o(pci_ad_o_8_) );
ms00f80 pci_io_mux_ad_iob8_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_8_) );
ms00f80 pci_io_mux_ad_iob9_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14322), .o(pci_ad_o_9_) );
ms00f80 pci_io_mux_ad_iob9_en_out_reg_u0 ( .ck(ispd_clk), .d(FE_OFN1505_n_15768), .o(pci_ad_oe_o_9_) );
ms00f80 pci_io_mux_cbe_iob0_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14393), .o(pci_cbe_o_0_) );
ms00f80 pci_io_mux_cbe_iob0_en_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23412), .o(pci_cbe_oe_o_0_) );
ms00f80 pci_io_mux_cbe_iob1_dat_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23414), .o(pci_cbe_o_1_) );
ms00f80 pci_io_mux_cbe_iob1_en_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23416), .o(pci_cbe_oe_o_1_) );
ms00f80 pci_io_mux_cbe_iob2_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14391), .o(pci_cbe_o_2_) );
ms00f80 pci_io_mux_cbe_iob2_en_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23418), .o(pci_cbe_oe_o_2_) );
ms00f80 pci_io_mux_cbe_iob3_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14388), .o(pci_cbe_o_3_) );
ms00f80 pci_io_mux_cbe_iob3_en_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23420), .o(pci_cbe_oe_o_3_) );
ms00f80 pci_io_mux_devsel_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14616), .o(pci_devsel_o) );
ms00f80 pci_io_mux_devsel_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_8934), .o(pci_devsel_oe_o) );
ms00f80 pci_io_mux_frame_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_8751), .o(pci_frame_o) );
ms00f80 pci_io_mux_frame_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_7211), .o(pci_frame_oe_o) );
ms00f80 pci_io_mux_irdy_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_2900), .o(pci_irdy_o) );
ms00f80 pci_io_mux_irdy_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_333), .o(pci_irdy_oe_o) );
ms00f80 pci_io_mux_par_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_8576), .o(pci_par_o) );
ms00f80 pci_io_mux_par_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_12855), .o(pci_par_oe_o) );
ms00f80 pci_io_mux_perr_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_13918), .o(pci_perr_o) );
ms00f80 pci_io_mux_perr_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_14571), .o(pci_perr_oe_o) );
ms00f80 pci_io_mux_req_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_2246), .o(pci_req_o) );
ms00f80 pci_io_mux_req_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_285), .o(pci_req_oe_o) );
ms00f80 pci_io_mux_serr_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_13917), .o(pci_serr_o) );
ms00f80 pci_io_mux_serr_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_13758), .o(pci_serr_oe_o) );
ms00f80 pci_io_mux_stop_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(n_14617), .o(pci_stop_o) );
ms00f80 pci_io_mux_stop_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_8934), .o(pci_stop_oe_o) );
ms00f80 pci_io_mux_trdy_iob_dat_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23422), .o(pci_trdy_o) );
ms00f80 pci_io_mux_trdy_iob_en_out_reg_u0 ( .ck(ispd_clk), .d(n_8934), .o(pci_trdy_oe_o) );
ms00f80 pci_resets_and_interrupts_inta_en_out_reg_u0 ( .ck(ispd_clk), .d(n_3315), .o(pci_inta_oe_o) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_0__u0 ( .ck(ispd_clk), .d(n_2672), .o(pci_target_unit_pcit_if_strd_addr_in) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_10__u0 ( .ck(ispd_clk), .d(n_2632), .o(pci_target_unit_pcit_if_strd_addr_in_695) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_11__u0 ( .ck(ispd_clk), .d(n_2635), .o(pci_target_unit_pcit_if_strd_addr_in_696) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_12__u0 ( .ck(ispd_clk), .d(n_2660), .o(pci_target_unit_pcit_if_strd_addr_in_697) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_13__u0 ( .ck(ispd_clk), .d(n_2658), .o(pci_target_unit_pcit_if_strd_addr_in_698) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_14__u0 ( .ck(ispd_clk), .d(n_2668), .o(pci_target_unit_pcit_if_strd_addr_in_699) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_15__u0 ( .ck(ispd_clk), .d(n_2673), .o(pci_target_unit_pcit_if_strd_addr_in_700) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_16__u0 ( .ck(ispd_clk), .d(n_2679), .o(pci_target_unit_pcit_if_strd_addr_in_701) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_17__u0 ( .ck(ispd_clk), .d(n_2636), .o(pci_target_unit_pcit_if_strd_addr_in_702) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_18__u0 ( .ck(ispd_clk), .d(n_2634), .o(pci_target_unit_pcit_if_strd_addr_in_703) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_19__u0 ( .ck(ispd_clk), .d(n_2638), .o(pci_target_unit_pcit_if_strd_addr_in_704) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2653), .o(pci_target_unit_pcit_if_strd_addr_in_686) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_20__u0 ( .ck(ispd_clk), .d(n_2646), .o(pci_target_unit_pcit_if_strd_addr_in_705) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_21__u0 ( .ck(ispd_clk), .d(n_2661), .o(pci_target_unit_pcit_if_strd_addr_in_706) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_22__u0 ( .ck(ispd_clk), .d(n_2659), .o(pci_target_unit_pcit_if_strd_addr_in_707) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_23__u0 ( .ck(ispd_clk), .d(n_2664), .o(pci_target_unit_pcit_if_strd_addr_in_708) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_24__u0 ( .ck(ispd_clk), .d(n_2665), .o(pci_target_unit_pcit_if_strd_addr_in_709) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_25__u0 ( .ck(ispd_clk), .d(n_2666), .o(pci_target_unit_pcit_if_strd_addr_in_710) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_26__u0 ( .ck(ispd_clk), .d(n_2669), .o(pci_target_unit_pcit_if_strd_addr_in_711) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_27__u0 ( .ck(ispd_clk), .d(n_2670), .o(pci_target_unit_pcit_if_strd_addr_in_712) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_28__u0 ( .ck(ispd_clk), .d(n_2674), .o(pci_target_unit_pcit_if_strd_addr_in_713) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_29__u0 ( .ck(ispd_clk), .d(n_2637), .o(pci_target_unit_pcit_if_strd_addr_in_714) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2640), .o(pci_target_unit_pcit_if_strd_addr_in_687) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_30__u0 ( .ck(ispd_clk), .d(n_2641), .o(pci_target_unit_pcit_if_strd_addr_in_715) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_31__u0 ( .ck(ispd_clk), .d(n_2656), .o(pci_target_unit_pcit_if_strd_addr_in_716) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2655), .o(pci_target_unit_pcit_if_strd_addr_in_688) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_4__u0 ( .ck(ispd_clk), .d(n_2639), .o(pci_target_unit_pcit_if_strd_addr_in_689) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_5__u0 ( .ck(ispd_clk), .d(n_2633), .o(pci_target_unit_pcit_if_strd_addr_in_690) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_6__u0 ( .ck(ispd_clk), .d(n_2645), .o(pci_target_unit_pcit_if_strd_addr_in_691) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_7__u0 ( .ck(ispd_clk), .d(n_2663), .o(pci_target_unit_pcit_if_strd_addr_in_692) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_8__u0 ( .ck(ispd_clk), .d(n_2667), .o(pci_target_unit_pcit_if_strd_addr_in_693) );
ms00f80 pci_target_unit_del_sync_addr_out_reg_9__u0 ( .ck(ispd_clk), .d(n_2654), .o(pci_target_unit_pcit_if_strd_addr_in_694) );
ms00f80 pci_target_unit_del_sync_bc_out_reg_0__u0 ( .ck(ispd_clk), .d(n_2644), .o(pci_target_unit_pcit_if_strd_bc_in) );
ms00f80 pci_target_unit_del_sync_bc_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2657), .o(pci_target_unit_pcit_if_strd_bc_in_717) );
ms00f80 pci_target_unit_del_sync_bc_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2662), .o(pci_target_unit_pcit_if_strd_bc_in_718) );
ms00f80 pci_target_unit_del_sync_bc_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2677), .o(pci_target_unit_pcit_if_strd_bc_in_719) );
ms00f80 pci_target_unit_del_sync_be_out_reg_0__u0 ( .ck(ispd_clk), .d(n_3031), .o(pci_target_unit_del_sync_be_out_reg_0__Q) );
ms00f80 pci_target_unit_del_sync_be_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2652), .o(pci_target_unit_del_sync_be_out_reg_1__Q) );
ms00f80 pci_target_unit_del_sync_be_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2649), .o(pci_target_unit_del_sync_be_out_reg_2__Q) );
ms00f80 pci_target_unit_del_sync_be_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2643), .o(pci_target_unit_del_sync_be_out_reg_3__Q) );
ms00f80 pci_target_unit_del_sync_burst_out_reg_u0 ( .ck(ispd_clk), .d(n_2676), .o(pci_target_unit_wbm_sm_pci_tar_burst_ok) );
ms00f80 pci_target_unit_del_sync_comp_comp_pending_reg_u0 ( .ck(ispd_clk), .d(n_7699), .o(wbu_pci_drcomp_pending_in) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_0__u0 ( .ck(ispd_clk), .d(n_2932), .o(pci_target_unit_del_sync_comp_cycle_count_0_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_10__u0 ( .ck(ispd_clk), .d(n_3171), .o(pci_target_unit_del_sync_comp_cycle_count_10_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_11__u0 ( .ck(ispd_clk), .d(n_3355), .o(pci_target_unit_del_sync_comp_cycle_count_11_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_12__u0 ( .ck(ispd_clk), .d(n_4153), .o(pci_target_unit_del_sync_comp_cycle_count_12_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_13__u0 ( .ck(ispd_clk), .d(n_3162), .o(pci_target_unit_del_sync_comp_cycle_count_13_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_14__u0 ( .ck(ispd_clk), .d(n_3490), .o(pci_target_unit_del_sync_comp_cycle_count_14_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_15__u0 ( .ck(ispd_clk), .d(n_3497), .o(pci_target_unit_del_sync_comp_cycle_count_15_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_16__u0 ( .ck(ispd_clk), .d(n_5744), .o(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_1__u0 ( .ck(ispd_clk), .d(n_2938), .o(pci_target_unit_del_sync_comp_cycle_count_1_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_2__u0 ( .ck(ispd_clk), .d(n_2953), .o(pci_target_unit_del_sync_comp_cycle_count_2_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_3__u0 ( .ck(ispd_clk), .d(n_2748), .o(pci_target_unit_del_sync_comp_cycle_count_3_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_4__u0 ( .ck(ispd_clk), .d(n_2774), .o(pci_target_unit_del_sync_comp_cycle_count_4_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_5__u0 ( .ck(ispd_clk), .d(n_2937), .o(pci_target_unit_del_sync_comp_cycle_count_5_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_6__u0 ( .ck(ispd_clk), .d(n_2980), .o(pci_target_unit_del_sync_comp_cycle_count_6_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_7__u0 ( .ck(ispd_clk), .d(n_2757), .o(pci_target_unit_del_sync_comp_cycle_count_7_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_8__u0 ( .ck(ispd_clk), .d(n_3028), .o(pci_target_unit_del_sync_comp_cycle_count_8_) );
ms00f80 pci_target_unit_del_sync_comp_cycle_count_reg_9__u0 ( .ck(ispd_clk), .d(n_2952), .o(pci_target_unit_del_sync_comp_cycle_count_9_) );
ms00f80 pci_target_unit_del_sync_comp_done_reg_clr_reg_u0 ( .ck(ispd_clk), .d(n_2146), .o(pci_target_unit_del_sync_comp_done_reg_clr_reg_Q) );
in01s01 pci_target_unit_del_sync_comp_done_reg_clr_reg_u1 ( .a(pci_target_unit_del_sync_comp_done_reg_clr_reg_Q), .o(pci_target_unit_del_sync_comp_done_reg_clr) );
ms00f80 pci_target_unit_del_sync_comp_done_reg_main_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_sync_comp_done), .o(pci_target_unit_del_sync_comp_done_reg_main_reg_Q) );
in01s03 pci_target_unit_del_sync_comp_done_reg_main_reg_u1 ( .a(pci_target_unit_del_sync_comp_done_reg_main_reg_Q), .o(pci_target_unit_del_sync_comp_done_reg_main) );
ms00f80 pci_target_unit_del_sync_comp_flush_out_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_comp_cycle_count_reg_16__Q), .o(pci_target_unit_del_sync_comp_flush_out_reg_Q) );
in01s01 pci_target_unit_del_sync_comp_flush_out_reg_u1 ( .a(pci_target_unit_del_sync_comp_flush_out_reg_Q), .o(pci_target_unit_pcit_if_comp_flush_in) );
ms00f80 pci_target_unit_del_sync_comp_req_pending_reg_u0 ( .ck(ispd_clk), .d(n_7706), .o(pci_target_unit_wbm_sm_pci_tar_read_request) );
ms00f80 pci_target_unit_del_sync_comp_rty_exp_clr_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_sync_comp_rty_exp_clr), .o(pci_target_unit_del_sync_comp_rty_exp_clr_reg_Q) );
in01s01 pci_target_unit_del_sync_comp_rty_exp_clr_reg_u1 ( .a(pci_target_unit_del_sync_comp_rty_exp_clr_reg_Q), .o(pci_target_unit_del_sync_comp_rty_exp_clr) );
ms00f80 pci_target_unit_del_sync_comp_rty_exp_reg_reg_u0 ( .ck(ispd_clk), .d(n_4711), .o(pci_target_unit_del_sync_comp_rty_exp_reg) );
ms00f80 pci_target_unit_del_sync_comp_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wbu_pci_drcomp_pending_in), .o(TIMEBOOST_net_21227) );
ms00f80 pci_target_unit_del_sync_done_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_req_done_reg), .o(pci_target_unit_del_sync_sync_comp_done) );
ms00f80 pci_target_unit_del_sync_req_comp_pending_reg_u0 ( .ck(ispd_clk), .d(n_3796), .o(pci_target_unit_del_sync_req_comp_pending) );
ms00f80 pci_target_unit_del_sync_req_comp_pending_sample_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_sync_req_comp_pending), .o(pci_target_unit_del_sync_req_comp_pending_sample_reg_Q) );
in01s01 pci_target_unit_del_sync_req_comp_pending_sample_reg_u1 ( .a(pci_target_unit_del_sync_req_comp_pending_sample_reg_Q), .o(pci_target_unit_del_sync_req_comp_pending_sample) );
ms00f80 pci_target_unit_del_sync_req_done_reg_reg_u0 ( .ck(ispd_clk), .d(n_4532), .o(pci_target_unit_del_sync_req_done_reg) );
ms00f80 pci_target_unit_del_sync_req_req_pending_reg_u0 ( .ck(ispd_clk), .d(n_2445), .o(pci_target_unit_pcit_if_req_req_pending_in) );
ms00f80 pci_target_unit_del_sync_req_rty_exp_clr_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_req_rty_exp_reg), .o(pci_target_unit_del_sync_req_rty_exp_clr_reg_Q) );
in01s01 pci_target_unit_del_sync_req_rty_exp_clr_reg_u1 ( .a(pci_target_unit_del_sync_req_rty_exp_clr_reg_Q), .o(pci_target_unit_del_sync_req_rty_exp_clr) );
ms00f80 pci_target_unit_del_sync_req_rty_exp_reg_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_sync_req_rty_exp), .o(pci_target_unit_del_sync_req_rty_exp_reg) );
ms00f80 pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_pcit_if_req_req_pending_in), .o(pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__Q) );
in01s01 pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__u1 ( .a(pci_target_unit_del_sync_req_sync_sync_data_out_reg_0__Q), .o(pci_target_unit_del_sync_sync_comp_req_pending) );
ms00f80 pci_target_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_738), .o(pci_target_unit_del_sync_sync_comp_rty_exp_clr) );
ms00f80 pci_target_unit_del_sync_rty_exp_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_del_sync_comp_rty_exp_reg), .o(pci_target_unit_del_sync_sync_req_rty_exp) );
ms00f80 pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_42), .o(pci_target_unit_fifos_wb_clk_sync_inGreyCount) );
ms00f80 pci_target_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_inGreyCount_reg_1__Q), .o(pci_target_unit_fifos_wb_clk_sync_inGreyCount_36) );
ms00f80 pci_target_unit_fifos_inGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(n_5547), .o(pci_target_unit_fifos_inGreyCount_reg_0__Q) );
in01s01 pci_target_unit_fifos_inGreyCount_reg_0__u1 ( .a(pci_target_unit_fifos_inGreyCount_reg_0__Q), .o(pci_target_unit_fifos_inGreyCount_0_) );
ms00f80 pci_target_unit_fifos_inGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(n_4798), .o(pci_target_unit_fifos_inGreyCount_reg_1__Q) );
ms00f80 pci_target_unit_fifos_outGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(n_13622), .o(pci_target_unit_fifos_outGreyCount_reg_0__Q) );
in01m20 pci_target_unit_fifos_outGreyCount_reg_0__u1 ( .a(pci_target_unit_fifos_outGreyCount_reg_0__Q), .o(pci_target_unit_fifos_outGreyCount_0_) );
ms00f80 pci_target_unit_fifos_outGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(n_13482), .o(pci_target_unit_fifos_outGreyCount_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23424), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23426), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_100) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_rgrey_addr_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23428), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_101) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_39) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_40) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__u0 ( .ck(ispd_clk), .d(n_9168), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_1__u0 ( .ck(ispd_clk), .d(n_8854), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__u0 ( .ck(ispd_clk), .d(n_8855), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__Q) );
in01f20 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_reg_2__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_plus_one_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__u0 ( .ck(ispd_clk), .d(n_8877), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__u0 ( .ck(ispd_clk), .d(n_8853), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__Q) );
in01m20 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_1__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__u0 ( .ck(ispd_clk), .d(n_8852), .o(pci_target_unit_fifos_pcir_fifo_ctrl_raddr_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__Q) );
in01f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_0__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_39), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__Q) );
in01f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_1__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_sync_wgrey_addr_40), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__Q) );
in01f80 pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__u1 ( .a(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_reg_2__Q), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rclk_wgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_8851), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_8850), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_8849), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_8848), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_8847), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_8846), .o(pci_target_unit_fifos_pcir_fifo_ctrl_rgrey_next_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg_0__u0 ( .ck(ispd_clk), .d(n_8501), .o(pci_target_unit_fifos_pcir_whole_waddr) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg_1__u0 ( .ck(ispd_clk), .d(n_8505), .o(pci_target_unit_fifos_pcir_whole_waddr_94) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_waddr_reg_2__u0 ( .ck(ispd_clk), .d(n_7836), .o(n_1117) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_100), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_sync_rgrey_addr_101), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wclk_rgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_7830), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_7833), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_7828), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_addr_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_8504), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_0_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_8502), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_1_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_7826), .o(pci_target_unit_fifos_pcir_fifo_ctrl_wgrey_next_2_) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_0__u0 ( .ck(ispd_clk), .d(n_12558), .o(pci_target_unit_pcit_if_pcir_fifo_data_in) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_10__u0 ( .ck(ispd_clk), .d(n_12557), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_775) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_11__u0 ( .ck(ispd_clk), .d(n_12556), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_776) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_12__u0 ( .ck(ispd_clk), .d(n_12555), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_777) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_13__u0 ( .ck(ispd_clk), .d(n_12554), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_778) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_14__u0 ( .ck(ispd_clk), .d(n_12553), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_779) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_15__u0 ( .ck(ispd_clk), .d(n_12771), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_780) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_16__u0 ( .ck(ispd_clk), .d(n_12552), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_781) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_17__u0 ( .ck(ispd_clk), .d(n_12551), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_782) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_18__u0 ( .ck(ispd_clk), .d(n_12550), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_783) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_19__u0 ( .ck(ispd_clk), .d(n_12549), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_784) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_1__u0 ( .ck(ispd_clk), .d(n_12548), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_766) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_20__u0 ( .ck(ispd_clk), .d(n_12547), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_785) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_21__u0 ( .ck(ispd_clk), .d(n_12546), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_786) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_22__u0 ( .ck(ispd_clk), .d(n_12545), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_787) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_23__u0 ( .ck(ispd_clk), .d(n_12544), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_788) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_24__u0 ( .ck(ispd_clk), .d(n_12543), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_789) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_25__u0 ( .ck(ispd_clk), .d(n_12770), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_790) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_26__u0 ( .ck(ispd_clk), .d(n_12542), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_791) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_27__u0 ( .ck(ispd_clk), .d(n_12541), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_792) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_28__u0 ( .ck(ispd_clk), .d(n_12540), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_793) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_29__u0 ( .ck(ispd_clk), .d(n_12539), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_794) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_2__u0 ( .ck(ispd_clk), .d(n_12538), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_767) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_30__u0 ( .ck(ispd_clk), .d(n_12537), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_795) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_31__u0 ( .ck(ispd_clk), .d(n_12536), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_796) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_37__u0 ( .ck(ispd_clk), .d(n_12535), .o(pci_target_unit_pcit_if_pcir_fifo_control_in_637) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_3__u0 ( .ck(ispd_clk), .d(n_12534), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_768) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_4__u0 ( .ck(ispd_clk), .d(n_12533), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_769) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_5__u0 ( .ck(ispd_clk), .d(n_12532), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_770) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_6__u0 ( .ck(ispd_clk), .d(n_12531), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_771) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_7__u0 ( .ck(ispd_clk), .d(n_12769), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_772) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_8__u0 ( .ck(ispd_clk), .d(n_12530), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_773) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_do_reg_b_reg_9__u0 ( .ck(ispd_clk), .d(n_12529), .o(pci_target_unit_pcit_if_pcir_fifo_data_in_774) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__u0 ( .ck(ispd_clk), .d(n_7915), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__u0 ( .ck(ispd_clk), .d(n_7913), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__u0 ( .ck(ispd_clk), .d(n_7911), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__u0 ( .ck(ispd_clk), .d(n_7909), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__u0 ( .ck(ispd_clk), .d(n_7907), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__u0 ( .ck(ispd_clk), .d(n_7905), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__u0 ( .ck(ispd_clk), .d(n_7903), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__u0 ( .ck(ispd_clk), .d(n_7901), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__u0 ( .ck(ispd_clk), .d(n_7899), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__u0 ( .ck(ispd_clk), .d(n_7897), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23430), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__u0 ( .ck(ispd_clk), .d(n_7893), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__u0 ( .ck(ispd_clk), .d(n_7891), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__u0 ( .ck(ispd_clk), .d(n_7889), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__u0 ( .ck(ispd_clk), .d(n_7887), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__u0 ( .ck(ispd_clk), .d(n_7885), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23432), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__u0 ( .ck(ispd_clk), .d(n_7881), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23434), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__u0 ( .ck(ispd_clk), .d(n_7877), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__u0 ( .ck(ispd_clk), .d(n_7875), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__u0 ( .ck(ispd_clk), .d(n_7873), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__u0 ( .ck(ispd_clk), .d(n_7871), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__u0 ( .ck(ispd_clk), .d(n_7869), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__u0 ( .ck(ispd_clk), .d(n_7867), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__u0 ( .ck(ispd_clk), .d(n_7865), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__u0 ( .ck(ispd_clk), .d(n_7863), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__u0 ( .ck(ispd_clk), .d(n_7861), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__u0 ( .ck(ispd_clk), .d(n_7859), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23436), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__u0 ( .ck(ispd_clk), .d(n_7855), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__u0 ( .ck(ispd_clk), .d(n_7853), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__u0 ( .ck(ispd_clk), .d(n_7851), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_0__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__u0 ( .ck(ispd_clk), .d(n_7849), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__u0 ( .ck(ispd_clk), .d(n_7847), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__u0 ( .ck(ispd_clk), .d(n_7844), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__u0 ( .ck(ispd_clk), .d(n_7842), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__u0 ( .ck(ispd_clk), .d(n_7840), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__u0 ( .ck(ispd_clk), .d(n_7838), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__u0 ( .ck(ispd_clk), .d(n_8123), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__u0 ( .ck(ispd_clk), .d(n_8121), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__u0 ( .ck(ispd_clk), .d(n_8118), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__u0 ( .ck(ispd_clk), .d(n_8116), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__u0 ( .ck(ispd_clk), .d(n_8114), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__u0 ( .ck(ispd_clk), .d(n_8111), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23438), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__u0 ( .ck(ispd_clk), .d(n_8107), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23440), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__u0 ( .ck(ispd_clk), .d(n_8102), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__u0 ( .ck(ispd_clk), .d(n_8100), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__u0 ( .ck(ispd_clk), .d(n_8097), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__u0 ( .ck(ispd_clk), .d(n_8094), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__u0 ( .ck(ispd_clk), .d(n_8092), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__u0 ( .ck(ispd_clk), .d(n_8089), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__u0 ( .ck(ispd_clk), .d(n_8087), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__u0 ( .ck(ispd_clk), .d(n_8084), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__u0 ( .ck(ispd_clk), .d(n_8082), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__u0 ( .ck(ispd_clk), .d(n_8079), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__u0 ( .ck(ispd_clk), .d(n_8076), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__u0 ( .ck(ispd_clk), .d(n_8073), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__u0 ( .ck(ispd_clk), .d(n_8071), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__u0 ( .ck(ispd_clk), .d(n_8068), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__u0 ( .ck(ispd_clk), .d(n_8066), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__u0 ( .ck(ispd_clk), .d(n_8064), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__u0 ( .ck(ispd_clk), .d(n_8062), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__u0 ( .ck(ispd_clk), .d(n_8059), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_1__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__u0 ( .ck(ispd_clk), .d(n_8056), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__u0 ( .ck(ispd_clk), .d(n_8054), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__u0 ( .ck(ispd_clk), .d(n_8052), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__u0 ( .ck(ispd_clk), .d(n_8049), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__u0 ( .ck(ispd_clk), .d(n_8047), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23442), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__u0 ( .ck(ispd_clk), .d(n_8041), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__u0 ( .ck(ispd_clk), .d(n_8039), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__u0 ( .ck(ispd_clk), .d(n_8036), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__u0 ( .ck(ispd_clk), .d(n_8034), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__u0 ( .ck(ispd_clk), .d(n_8032), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__u0 ( .ck(ispd_clk), .d(n_8030), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__u0 ( .ck(ispd_clk), .d(n_8027), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__u0 ( .ck(ispd_clk), .d(n_8024), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__u0 ( .ck(ispd_clk), .d(n_8021), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__u0 ( .ck(ispd_clk), .d(n_8019), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__u0 ( .ck(ispd_clk), .d(n_8017), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__u0 ( .ck(ispd_clk), .d(n_8014), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23444), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__u0 ( .ck(ispd_clk), .d(n_8009), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__u0 ( .ck(ispd_clk), .d(n_8007), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__u0 ( .ck(ispd_clk), .d(n_8005), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__u0 ( .ck(ispd_clk), .d(n_8003), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__u0 ( .ck(ispd_clk), .d(n_8001), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__u0 ( .ck(ispd_clk), .d(n_7999), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__u0 ( .ck(ispd_clk), .d(n_7997), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__u0 ( .ck(ispd_clk), .d(n_7995), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__u0 ( .ck(ispd_clk), .d(n_7993), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__u0 ( .ck(ispd_clk), .d(n_7991), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__u0 ( .ck(ispd_clk), .d(n_7989), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__u0 ( .ck(ispd_clk), .d(n_7987), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__u0 ( .ck(ispd_clk), .d(n_7985), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__u0 ( .ck(ispd_clk), .d(n_7983), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_2__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__u0 ( .ck(ispd_clk), .d(n_7981), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__u0 ( .ck(ispd_clk), .d(n_7979), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__u0 ( .ck(ispd_clk), .d(n_7977), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__u0 ( .ck(ispd_clk), .d(n_7975), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__u0 ( .ck(ispd_clk), .d(n_7973), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__u0 ( .ck(ispd_clk), .d(n_7971), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__u0 ( .ck(ispd_clk), .d(n_7969), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__u0 ( .ck(ispd_clk), .d(n_7967), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__u0 ( .ck(ispd_clk), .d(n_7965), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__u0 ( .ck(ispd_clk), .d(n_7963), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__u0 ( .ck(ispd_clk), .d(n_7961), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__u0 ( .ck(ispd_clk), .d(n_7959), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23446), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__u0 ( .ck(ispd_clk), .d(n_7955), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__u0 ( .ck(ispd_clk), .d(n_7953), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__u0 ( .ck(ispd_clk), .d(n_7951), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__u0 ( .ck(ispd_clk), .d(n_7949), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__u0 ( .ck(ispd_clk), .d(n_7947), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__u0 ( .ck(ispd_clk), .d(n_7945), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23448), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__u0 ( .ck(ispd_clk), .d(n_7941), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__u0 ( .ck(ispd_clk), .d(n_7939), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__u0 ( .ck(ispd_clk), .d(n_7937), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__u0 ( .ck(ispd_clk), .d(n_7935), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__u0 ( .ck(ispd_clk), .d(n_7933), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__u0 ( .ck(ispd_clk), .d(n_7931), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__u0 ( .ck(ispd_clk), .d(n_7929), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__u0 ( .ck(ispd_clk), .d(n_7927), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__u0 ( .ck(ispd_clk), .d(n_7925), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__u0 ( .ck(ispd_clk), .d(n_7923), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__u0 ( .ck(ispd_clk), .d(n_7921), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__u0 ( .ck(ispd_clk), .d(n_7919), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__u0 ( .ck(ispd_clk), .d(n_7917), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_3__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__u0 ( .ck(ispd_clk), .d(n_8430), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__u0 ( .ck(ispd_clk), .d(n_8428), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__u0 ( .ck(ispd_clk), .d(n_8426), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__u0 ( .ck(ispd_clk), .d(n_8423), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__u0 ( .ck(ispd_clk), .d(n_8421), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__u0 ( .ck(ispd_clk), .d(n_8419), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__u0 ( .ck(ispd_clk), .d(n_8417), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__u0 ( .ck(ispd_clk), .d(n_8415), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__u0 ( .ck(ispd_clk), .d(n_8413), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__u0 ( .ck(ispd_clk), .d(n_8411), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__u0 ( .ck(ispd_clk), .d(n_8409), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__u0 ( .ck(ispd_clk), .d(n_8406), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__u0 ( .ck(ispd_clk), .d(n_8404), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__u0 ( .ck(ispd_clk), .d(n_8402), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__u0 ( .ck(ispd_clk), .d(n_8400), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__u0 ( .ck(ispd_clk), .d(n_8397), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__u0 ( .ck(ispd_clk), .d(n_8395), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__u0 ( .ck(ispd_clk), .d(n_8393), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__u0 ( .ck(ispd_clk), .d(n_8391), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__u0 ( .ck(ispd_clk), .d(n_8389), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__u0 ( .ck(ispd_clk), .d(n_8387), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__u0 ( .ck(ispd_clk), .d(n_8384), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__u0 ( .ck(ispd_clk), .d(n_8382), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__u0 ( .ck(ispd_clk), .d(n_8379), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__u0 ( .ck(ispd_clk), .d(n_8376), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__u0 ( .ck(ispd_clk), .d(n_8373), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__u0 ( .ck(ispd_clk), .d(n_8371), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__u0 ( .ck(ispd_clk), .d(n_8368), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__u0 ( .ck(ispd_clk), .d(n_8366), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__u0 ( .ck(ispd_clk), .d(n_8364), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__u0 ( .ck(ispd_clk), .d(n_8362), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__u0 ( .ck(ispd_clk), .d(n_8360), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__u0 ( .ck(ispd_clk), .d(n_8358), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_4__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__u0 ( .ck(ispd_clk), .d(n_8355), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__u0 ( .ck(ispd_clk), .d(n_8353), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__u0 ( .ck(ispd_clk), .d(n_8351), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__u0 ( .ck(ispd_clk), .d(n_8349), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__u0 ( .ck(ispd_clk), .d(n_8346), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__u0 ( .ck(ispd_clk), .d(n_8344), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__u0 ( .ck(ispd_clk), .d(n_8341), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__u0 ( .ck(ispd_clk), .d(n_8339), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__u0 ( .ck(ispd_clk), .d(n_8337), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__u0 ( .ck(ispd_clk), .d(n_8335), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__u0 ( .ck(ispd_clk), .d(n_8333), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__u0 ( .ck(ispd_clk), .d(n_8331), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__u0 ( .ck(ispd_clk), .d(n_8329), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__u0 ( .ck(ispd_clk), .d(n_8327), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__u0 ( .ck(ispd_clk), .d(n_8325), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23450), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__u0 ( .ck(ispd_clk), .d(n_8321), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__u0 ( .ck(ispd_clk), .d(n_8319), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23452), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__u0 ( .ck(ispd_clk), .d(n_8313), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__u0 ( .ck(ispd_clk), .d(n_8311), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__u0 ( .ck(ispd_clk), .d(n_8309), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__u0 ( .ck(ispd_clk), .d(n_8307), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__u0 ( .ck(ispd_clk), .d(n_8304), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__u0 ( .ck(ispd_clk), .d(n_8302), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__u0 ( .ck(ispd_clk), .d(n_8299), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__u0 ( .ck(ispd_clk), .d(n_8297), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23454), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__u0 ( .ck(ispd_clk), .d(n_8293), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23456), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__u0 ( .ck(ispd_clk), .d(n_8288), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__u0 ( .ck(ispd_clk), .d(n_8285), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__u0 ( .ck(ispd_clk), .d(n_8283), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_5__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__u0 ( .ck(ispd_clk), .d(n_8281), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__u0 ( .ck(ispd_clk), .d(n_8279), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__u0 ( .ck(ispd_clk), .d(n_8277), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__u0 ( .ck(ispd_clk), .d(n_8274), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__u0 ( .ck(ispd_clk), .d(n_8271), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__u0 ( .ck(ispd_clk), .d(n_8269), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__u0 ( .ck(ispd_clk), .d(n_8267), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__u0 ( .ck(ispd_clk), .d(n_8264), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__u0 ( .ck(ispd_clk), .d(n_8262), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__u0 ( .ck(ispd_clk), .d(n_8260), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__u0 ( .ck(ispd_clk), .d(n_8258), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__u0 ( .ck(ispd_clk), .d(n_8255), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__u0 ( .ck(ispd_clk), .d(n_8253), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__u0 ( .ck(ispd_clk), .d(n_8251), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__u0 ( .ck(ispd_clk), .d(n_8248), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__u0 ( .ck(ispd_clk), .d(n_8246), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__u0 ( .ck(ispd_clk), .d(n_8244), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__u0 ( .ck(ispd_clk), .d(n_8241), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__u0 ( .ck(ispd_clk), .d(n_8239), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__u0 ( .ck(ispd_clk), .d(n_8236), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__u0 ( .ck(ispd_clk), .d(n_8234), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__u0 ( .ck(ispd_clk), .d(n_8231), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23458), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__u0 ( .ck(ispd_clk), .d(n_8226), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__u0 ( .ck(ispd_clk), .d(n_8223), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__u0 ( .ck(ispd_clk), .d(n_8220), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__u0 ( .ck(ispd_clk), .d(n_8218), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__u0 ( .ck(ispd_clk), .d(n_8215), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__u0 ( .ck(ispd_clk), .d(n_8213), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__u0 ( .ck(ispd_clk), .d(n_8210), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__u0 ( .ck(ispd_clk), .d(n_8208), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__u0 ( .ck(ispd_clk), .d(n_8205), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__u0 ( .ck(ispd_clk), .d(n_8203), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_6__9__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__u0 ( .ck(ispd_clk), .d(n_8200), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__0__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__u0 ( .ck(ispd_clk), .d(n_8198), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__10__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__u0 ( .ck(ispd_clk), .d(n_8196), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__11__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__u0 ( .ck(ispd_clk), .d(n_8193), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__12__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__u0 ( .ck(ispd_clk), .d(n_8191), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__13__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__u0 ( .ck(ispd_clk), .d(n_8189), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__14__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__u0 ( .ck(ispd_clk), .d(n_8186), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__15__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__u0 ( .ck(ispd_clk), .d(n_8184), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__16__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__u0 ( .ck(ispd_clk), .d(n_8182), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__17__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__u0 ( .ck(ispd_clk), .d(n_8180), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__18__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23460), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__19__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__u0 ( .ck(ispd_clk), .d(n_8175), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__1__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__u0 ( .ck(ispd_clk), .d(n_8173), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__20__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__u0 ( .ck(ispd_clk), .d(n_8171), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__21__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__u0 ( .ck(ispd_clk), .d(n_8168), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__22__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23462), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__23__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__u0 ( .ck(ispd_clk), .d(n_8163), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__24__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__u0 ( .ck(ispd_clk), .d(n_8161), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__25__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__u0 ( .ck(ispd_clk), .d(n_8159), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__26__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__u0 ( .ck(ispd_clk), .d(n_8157), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__27__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__u0 ( .ck(ispd_clk), .d(n_8154), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__28__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__u0 ( .ck(ispd_clk), .d(n_8152), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__29__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__u0 ( .ck(ispd_clk), .d(n_8150), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__2__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__u0 ( .ck(ispd_clk), .d(n_8147), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__30__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23464), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__31__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__u0 ( .ck(ispd_clk), .d(n_8142), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__37__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__u0 ( .ck(ispd_clk), .d(n_8139), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__3__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__u0 ( .ck(ispd_clk), .d(n_8137), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__4__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__u0 ( .ck(ispd_clk), .d(n_8135), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__5__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__u0 ( .ck(ispd_clk), .d(n_8132), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__6__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__u0 ( .ck(ispd_clk), .d(n_8130), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__7__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__u0 ( .ck(ispd_clk), .d(n_8128), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__8__Q) );
ms00f80 pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__u0 ( .ck(ispd_clk), .d(n_8125), .o(pci_target_unit_fifos_pcir_fifo_storage_mem_reg_7__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus2) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_94) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_rgrey_minus2_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_95) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23466), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23468), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_74) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23470), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_75) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__u0 ( .ck(ispd_clk), .d(n_13682), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__u0 ( .ck(ispd_clk), .d(n_13619), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__u0 ( .ck(ispd_clk), .d(n_13618), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_plus_one_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__u0 ( .ck(ispd_clk), .d(n_16970), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__u0 ( .ck(ispd_clk), .d(n_13479), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__u0 ( .ck(ispd_clk), .d(n_13475), .o(pci_target_unit_fifos_pciw_fifo_ctrl_raddr_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_74), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_sync_wgrey_addr_75), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rclk_wgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_13616), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_13614), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_13613), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23472), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__u0 ( .ck(ispd_clk), .d(n_13609), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__u0 ( .ck(ispd_clk), .d(n_13607), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus1_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__u0 ( .ck(ispd_clk), .d(n_13605), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__u0 ( .ck(ispd_clk), .d(n_13603), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__u0 ( .ck(ispd_clk), .d(n_13601), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_minus2_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_13599), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_13597), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_13595), .o(pci_target_unit_fifos_pciw_fifo_ctrl_rgrey_next_reg_2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg_0__u0 ( .ck(ispd_clk), .d(n_4616), .o(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg_1__u0 ( .ck(ispd_clk), .d(n_4639), .o(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_reg_2__u0 ( .ck(ispd_clk), .d(n_4130), .o(pci_target_unit_fifos_pciw_fifo_ctrl_waddr_plus1_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg_0__u0 ( .ck(ispd_clk), .d(n_4614), .o(pci_target_unit_fifos_pciw_whole_waddr) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg_1__u0 ( .ck(ispd_clk), .d(n_4634), .o(pci_target_unit_fifos_pciw_whole_waddr_47) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_waddr_reg_2__u0 ( .ck(ispd_clk), .d(n_4134), .o(n_1293) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus2), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_94), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_reg_2__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_sync_rgrey_minus_95), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wclk_rgrey_minus2_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_4115), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_4107), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_4114), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_addr_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg_0__u0 ( .ck(ispd_clk), .d(n_4113), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg_1__u0 ( .ck(ispd_clk), .d(n_4108), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_reg_2__u0 ( .ck(ispd_clk), .d(n_4112), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_minus1_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg_0__u0 ( .ck(ispd_clk), .d(n_4638), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg_1__u0 ( .ck(ispd_clk), .d(n_4138), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_reg_2__u0 ( .ck(ispd_clk), .d(n_4109), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_plus1_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_4636), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_0_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_4632), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_1_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_4111), .o(pci_target_unit_fifos_pciw_fifo_ctrl_wgrey_next_2_) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_0__u0 ( .ck(ispd_clk), .d(n_14613), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_10__u0 ( .ck(ispd_clk), .d(n_14614), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_59) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_11__u0 ( .ck(ispd_clk), .d(n_14612), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_60) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_12__u0 ( .ck(ispd_clk), .d(n_14611), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_61) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_13__u0 ( .ck(ispd_clk), .d(n_14610), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_62) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_14__u0 ( .ck(ispd_clk), .d(n_14609), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_63) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_15__u0 ( .ck(ispd_clk), .d(n_16247), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_64) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_16__u0 ( .ck(ispd_clk), .d(n_14608), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_65) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_17__u0 ( .ck(ispd_clk), .d(n_14607), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_66) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_18__u0 ( .ck(ispd_clk), .d(n_16254), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_67) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_19__u0 ( .ck(ispd_clk), .d(n_16224), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_68) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_1__u0 ( .ck(ispd_clk), .d(n_14605), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_50) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_20__u0 ( .ck(ispd_clk), .d(n_14604), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_69) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_21__u0 ( .ck(ispd_clk), .d(n_14603), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_70) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_22__u0 ( .ck(ispd_clk), .d(n_14602), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_71) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_23__u0 ( .ck(ispd_clk), .d(n_14601), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_72) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_24__u0 ( .ck(ispd_clk), .d(n_16231), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_73) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_25__u0 ( .ck(ispd_clk), .d(n_14599), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_74) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_26__u0 ( .ck(ispd_clk), .d(n_14598), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_75) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_27__u0 ( .ck(ispd_clk), .d(n_14597), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_76) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_28__u0 ( .ck(ispd_clk), .d(n_14596), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_77) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_29__u0 ( .ck(ispd_clk), .d(n_14595), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_78) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_2__u0 ( .ck(ispd_clk), .d(n_14594), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_51) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_30__u0 ( .ck(ispd_clk), .d(n_14593), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_79) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_31__u0 ( .ck(ispd_clk), .d(n_14592), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_80) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_32__u0 ( .ck(ispd_clk), .d(n_14591), .o(pci_target_unit_wbm_sm_pciw_fifo_cbe_in) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_33__u0 ( .ck(ispd_clk), .d(n_14590), .o(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_81) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_34__u0 ( .ck(ispd_clk), .d(n_14589), .o(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_82) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_35__u0 ( .ck(ispd_clk), .d(n_14588), .o(pci_target_unit_wbm_sm_pciw_fifo_cbe_in_83) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_36__u0 ( .ck(ispd_clk), .d(n_16213), .o(pci_target_unit_wbm_sm_pciw_fifo_control_in) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__u0 ( .ck(ispd_clk), .d(n_14585), .o(pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__Q) );
in01f10 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_37__Q), .o(pci_target_unit_wbm_sm_pciw_fifo_control_in_84) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_38__u0 ( .ck(ispd_clk), .d(n_16173), .o(pci_target_unit_wbm_sm_pciw_fifo_control_in_85) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_39__u0 ( .ck(ispd_clk), .d(n_14583), .o(pci_target_unit_wbm_sm_pciw_fifo_control_in_86) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_3__u0 ( .ck(ispd_clk), .d(n_14582), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_52) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_4__u0 ( .ck(ispd_clk), .d(n_16240), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_53) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_5__u0 ( .ck(ispd_clk), .d(n_14580), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_54) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_6__u0 ( .ck(ispd_clk), .d(n_14579), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_55) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_7__u0 ( .ck(ispd_clk), .d(n_16261), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_56) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_8__u0 ( .ck(ispd_clk), .d(n_14578), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_57) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_do_reg_b_reg_9__u0 ( .ck(ispd_clk), .d(n_14577), .o(pci_target_unit_wbm_sm_pciw_fifo_addr_data_in_58) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__u0 ( .ck(ispd_clk), .d(n_6963), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__u0 ( .ck(ispd_clk), .d(n_5225), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__u0 ( .ck(ispd_clk), .d(n_5223), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__u0 ( .ck(ispd_clk), .d(n_5221), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__u0 ( .ck(ispd_clk), .d(n_5218), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__u0 ( .ck(ispd_clk), .d(n_5216), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__u0 ( .ck(ispd_clk), .d(n_5214), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__u0 ( .ck(ispd_clk), .d(n_5212), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__u0 ( .ck(ispd_clk), .d(n_5207), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__u0 ( .ck(ispd_clk), .d(n_5203), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__u0 ( .ck(ispd_clk), .d(n_5200), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__u0 ( .ck(ispd_clk), .d(n_6961), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__u0 ( .ck(ispd_clk), .d(n_5198), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__u0 ( .ck(ispd_clk), .d(n_5196), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__u0 ( .ck(ispd_clk), .d(n_5194), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__u0 ( .ck(ispd_clk), .d(n_5192), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__u0 ( .ck(ispd_clk), .d(n_5190), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__u0 ( .ck(ispd_clk), .d(n_5188), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__u0 ( .ck(ispd_clk), .d(n_5185), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__u0 ( .ck(ispd_clk), .d(n_5183), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__u0 ( .ck(ispd_clk), .d(n_5181), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__u0 ( .ck(ispd_clk), .d(n_5179), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__u0 ( .ck(ispd_clk), .d(n_4963), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__u0 ( .ck(ispd_clk), .d(n_5176), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__u0 ( .ck(ispd_clk), .d(n_5174), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__u0 ( .ck(ispd_clk), .d(n_7125), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__u0 ( .ck(ispd_clk), .d(n_5170), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__u0 ( .ck(ispd_clk), .d(n_5168), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__u0 ( .ck(ispd_clk), .d(n_5166), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__u0 ( .ck(ispd_clk), .d(n_7123), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__Q) );
in01m20 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__36__Q), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_0__153) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__u0 ( .ck(ispd_clk), .d(n_7681), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__u0 ( .ck(ispd_clk), .d(n_4926), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__u0 ( .ck(ispd_clk), .d(n_4605), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__u0 ( .ck(ispd_clk), .d(n_5163), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__u0 ( .ck(ispd_clk), .d(n_5161), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__u0 ( .ck(ispd_clk), .d(n_5158), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__u0 ( .ck(ispd_clk), .d(n_5156), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__u0 ( .ck(ispd_clk), .d(n_5153), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__u0 ( .ck(ispd_clk), .d(n_5151), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__u0 ( .ck(ispd_clk), .d(n_5146), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_0__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__u0 ( .ck(ispd_clk), .d(n_6956), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__u0 ( .ck(ispd_clk), .d(n_5140), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__u0 ( .ck(ispd_clk), .d(n_5138), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__u0 ( .ck(ispd_clk), .d(n_4978), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__u0 ( .ck(ispd_clk), .d(n_5136), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__u0 ( .ck(ispd_clk), .d(n_5134), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__u0 ( .ck(ispd_clk), .d(n_5132), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__u0 ( .ck(ispd_clk), .d(n_4959), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__u0 ( .ck(ispd_clk), .d(n_5130), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__u0 ( .ck(ispd_clk), .d(n_5128), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__u0 ( .ck(ispd_clk), .d(n_5126), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__u0 ( .ck(ispd_clk), .d(n_6953), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__u0 ( .ck(ispd_clk), .d(n_5124), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__u0 ( .ck(ispd_clk), .d(n_5120), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__u0 ( .ck(ispd_clk), .d(n_5118), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__u0 ( .ck(ispd_clk), .d(n_5116), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__u0 ( .ck(ispd_clk), .d(n_5114), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__u0 ( .ck(ispd_clk), .d(n_5112), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__u0 ( .ck(ispd_clk), .d(n_5110), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__u0 ( .ck(ispd_clk), .d(n_5108), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__u0 ( .ck(ispd_clk), .d(n_5106), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__u0 ( .ck(ispd_clk), .d(n_5104), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__u0 ( .ck(ispd_clk), .d(n_5102), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__u0 ( .ck(ispd_clk), .d(n_5100), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__u0 ( .ck(ispd_clk), .d(n_5098), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__u0 ( .ck(ispd_clk), .d(n_7121), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__u0 ( .ck(ispd_clk), .d(n_5096), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__u0 ( .ck(ispd_clk), .d(n_5094), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__u0 ( .ck(ispd_clk), .d(n_5092), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__u0 ( .ck(ispd_clk), .d(n_7119), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__Q) );
in01m20 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__36__Q), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_1__192) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__u0 ( .ck(ispd_clk), .d(n_7679), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__u0 ( .ck(ispd_clk), .d(n_4924), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__u0 ( .ck(ispd_clk), .d(n_4603), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__u0 ( .ck(ispd_clk), .d(n_5088), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__u0 ( .ck(ispd_clk), .d(n_5086), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__u0 ( .ck(ispd_clk), .d(n_5084), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__u0 ( .ck(ispd_clk), .d(n_5082), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__u0 ( .ck(ispd_clk), .d(n_5080), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__u0 ( .ck(ispd_clk), .d(n_5078), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__u0 ( .ck(ispd_clk), .d(n_5076), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_1__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__u0 ( .ck(ispd_clk), .d(n_6951), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__u0 ( .ck(ispd_clk), .d(n_5074), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__u0 ( .ck(ispd_clk), .d(n_5071), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__u0 ( .ck(ispd_clk), .d(n_5068), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__u0 ( .ck(ispd_clk), .d(n_5064), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__u0 ( .ck(ispd_clk), .d(n_5060), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__u0 ( .ck(ispd_clk), .d(n_5058), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__u0 ( .ck(ispd_clk), .d(n_5056), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__u0 ( .ck(ispd_clk), .d(n_5054), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__u0 ( .ck(ispd_clk), .d(n_5052), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__u0 ( .ck(ispd_clk), .d(n_5050), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__u0 ( .ck(ispd_clk), .d(n_6948), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__u0 ( .ck(ispd_clk), .d(n_5048), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__u0 ( .ck(ispd_clk), .d(n_5046), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__u0 ( .ck(ispd_clk), .d(n_5044), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__u0 ( .ck(ispd_clk), .d(n_5042), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__u0 ( .ck(ispd_clk), .d(n_5040), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__u0 ( .ck(ispd_clk), .d(n_5038), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__u0 ( .ck(ispd_clk), .d(n_5036), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__u0 ( .ck(ispd_clk), .d(n_5033), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__u0 ( .ck(ispd_clk), .d(n_5031), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__u0 ( .ck(ispd_clk), .d(n_5029), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__u0 ( .ck(ispd_clk), .d(n_5027), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__u0 ( .ck(ispd_clk), .d(n_5025), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__u0 ( .ck(ispd_clk), .d(n_5023), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__u0 ( .ck(ispd_clk), .d(n_7117), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__u0 ( .ck(ispd_clk), .d(n_5021), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__u0 ( .ck(ispd_clk), .d(n_5018), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__u0 ( .ck(ispd_clk), .d(n_5016), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__u0 ( .ck(ispd_clk), .d(n_7126), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__Q) );
in01m20 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__36__Q), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_2__231) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__u0 ( .ck(ispd_clk), .d(n_7683), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__u0 ( .ck(ispd_clk), .d(n_4922), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__u0 ( .ck(ispd_clk), .d(n_4607), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__u0 ( .ck(ispd_clk), .d(n_5066), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__u0 ( .ck(ispd_clk), .d(n_5205), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__u0 ( .ck(ispd_clk), .d(n_4957), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__u0 ( .ck(ispd_clk), .d(n_5014), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__u0 ( .ck(ispd_clk), .d(n_4961), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__u0 ( .ck(ispd_clk), .d(n_5012), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__u0 ( .ck(ispd_clk), .d(n_5062), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_2__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__u0 ( .ck(ispd_clk), .d(n_6946), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__u0 ( .ck(ispd_clk), .d(n_5009), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__u0 ( .ck(ispd_clk), .d(n_5149), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__u0 ( .ck(ispd_clk), .d(n_5090), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__u0 ( .ck(ispd_clk), .d(n_5006), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__u0 ( .ck(ispd_clk), .d(n_5003), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__u0 ( .ck(ispd_clk), .d(n_5122), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__u0 ( .ck(ispd_clk), .d(n_5001), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__u0 ( .ck(ispd_clk), .d(n_5143), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__u0 ( .ck(ispd_clk), .d(n_4999), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__u0 ( .ck(ispd_clk), .d(n_5172), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__u0 ( .ck(ispd_clk), .d(n_6958), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__u0 ( .ck(ispd_clk), .d(n_4996), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__u0 ( .ck(ispd_clk), .d(n_4993), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__u0 ( .ck(ispd_clk), .d(n_5210), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__u0 ( .ck(ispd_clk), .d(n_4991), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__u0 ( .ck(ispd_clk), .d(n_4988), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__u0 ( .ck(ispd_clk), .d(n_4986), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__u0 ( .ck(ispd_clk), .d(n_5227), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__u0 ( .ck(ispd_clk), .d(n_4984), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__u0 ( .ck(ispd_clk), .d(n_4941), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__u0 ( .ck(ispd_clk), .d(n_4982), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__u0 ( .ck(ispd_clk), .d(n_4943), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__u0 ( .ck(ispd_clk), .d(n_4980), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__u0 ( .ck(ispd_clk), .d(n_4945), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__u0 ( .ck(ispd_clk), .d(n_7112), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__u0 ( .ck(ispd_clk), .d(n_4949), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__u0 ( .ck(ispd_clk), .d(n_4955), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__u0 ( .ck(ispd_clk), .d(n_4953), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__u0 ( .ck(ispd_clk), .d(n_7122), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__Q) );
in01s01 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__u1 ( .a(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__36__Q), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_3__270) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__u0 ( .ck(ispd_clk), .d(n_7677), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__u0 ( .ck(ispd_clk), .d(n_4920), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__u0 ( .ck(ispd_clk), .d(n_4601), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__u0 ( .ck(ispd_clk), .d(n_4975), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__u0 ( .ck(ispd_clk), .d(n_4947), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__u0 ( .ck(ispd_clk), .d(n_4973), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__u0 ( .ck(ispd_clk), .d(n_4970), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__u0 ( .ck(ispd_clk), .d(n_4968), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__u0 ( .ck(ispd_clk), .d(n_4951), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__u0 ( .ck(ispd_clk), .d(n_4965), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_3__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__u0 ( .ck(ispd_clk), .d(n_6977), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__u0 ( .ck(ispd_clk), .d(n_5414), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__u0 ( .ck(ispd_clk), .d(n_5308), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__u0 ( .ck(ispd_clk), .d(n_5361), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__u0 ( .ck(ispd_clk), .d(n_5363), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__u0 ( .ck(ispd_clk), .d(n_5366), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__u0 ( .ck(ispd_clk), .d(n_5371), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__u0 ( .ck(ispd_clk), .d(n_5380), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__u0 ( .ck(ispd_clk), .d(n_5386), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__u0 ( .ck(ispd_clk), .d(n_5388), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__u0 ( .ck(ispd_clk), .d(n_5409), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__u0 ( .ck(ispd_clk), .d(n_6975), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__u0 ( .ck(ispd_clk), .d(n_5290), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__u0 ( .ck(ispd_clk), .d(n_5303), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__u0 ( .ck(ispd_clk), .d(n_5300), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__u0 ( .ck(ispd_clk), .d(n_5406), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__u0 ( .ck(ispd_clk), .d(n_5404), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__u0 ( .ck(ispd_clk), .d(n_5318), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__u0 ( .ck(ispd_clk), .d(n_5402), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__u0 ( .ck(ispd_clk), .d(n_5337), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__u0 ( .ck(ispd_clk), .d(n_5399), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__u0 ( .ck(ispd_clk), .d(n_5354), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__u0 ( .ck(ispd_clk), .d(n_5418), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__u0 ( .ck(ispd_clk), .d(n_5421), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__u0 ( .ck(ispd_clk), .d(n_5396), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__u0 ( .ck(ispd_clk), .d(n_7128), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__u0 ( .ck(ispd_clk), .d(n_5393), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__u0 ( .ck(ispd_clk), .d(n_5391), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__u0 ( .ck(ispd_clk), .d(n_5305), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__u0 ( .ck(ispd_clk), .d(n_6115), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__36__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__u0 ( .ck(ispd_clk), .d(n_7692), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__u0 ( .ck(ispd_clk), .d(n_4928), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__u0 ( .ck(ispd_clk), .d(n_4623), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__u0 ( .ck(ispd_clk), .d(n_5323), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__u0 ( .ck(ispd_clk), .d(n_5332), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__u0 ( .ck(ispd_clk), .d(n_5315), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__u0 ( .ck(ispd_clk), .d(n_5412), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__u0 ( .ck(ispd_clk), .d(n_5267), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__u0 ( .ck(ispd_clk), .d(n_5416), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__u0 ( .ck(ispd_clk), .d(n_5448), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_4__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__u0 ( .ck(ispd_clk), .d(n_6971), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__u0 ( .ck(ispd_clk), .d(n_5383), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__u0 ( .ck(ispd_clk), .d(n_5265), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__u0 ( .ck(ispd_clk), .d(n_5378), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__u0 ( .ck(ispd_clk), .d(n_5275), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__u0 ( .ck(ispd_clk), .d(n_5376), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__u0 ( .ck(ispd_clk), .d(n_5281), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__u0 ( .ck(ispd_clk), .d(n_5288), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__u0 ( .ck(ispd_clk), .d(n_5296), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__u0 ( .ck(ispd_clk), .d(n_5373), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__u0 ( .ck(ispd_clk), .d(n_5298), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__u0 ( .ck(ispd_clk), .d(n_6967), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__u0 ( .ck(ispd_clk), .d(n_5237), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__u0 ( .ck(ispd_clk), .d(n_5368), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__u0 ( .ck(ispd_clk), .d(n_5244), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__u0 ( .ck(ispd_clk), .d(n_5255), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__u0 ( .ck(ispd_clk), .d(n_5258), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__u0 ( .ck(ispd_clk), .d(n_5424), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__u0 ( .ck(ispd_clk), .d(n_5429), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__u0 ( .ck(ispd_clk), .d(n_5433), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__u0 ( .ck(ispd_clk), .d(n_5441), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__u0 ( .ck(ispd_clk), .d(n_5450), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__u0 ( .ck(ispd_clk), .d(n_5458), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__u0 ( .ck(ispd_clk), .d(n_5461), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__u0 ( .ck(ispd_clk), .d(n_5463), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__u0 ( .ck(ispd_clk), .d(n_7134), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__u0 ( .ck(ispd_clk), .d(n_5478), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__u0 ( .ck(ispd_clk), .d(n_5481), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__u0 ( .ck(ispd_clk), .d(n_5491), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__u0 ( .ck(ispd_clk), .d(n_6132), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__36__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__u0 ( .ck(ispd_clk), .d(n_7689), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__u0 ( .ck(ispd_clk), .d(n_4932), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__u0 ( .ck(ispd_clk), .d(n_4627), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__u0 ( .ck(ispd_clk), .d(n_5493), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__u0 ( .ck(ispd_clk), .d(n_5497), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__u0 ( .ck(ispd_clk), .d(n_5501), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__u0 ( .ck(ispd_clk), .d(n_5505), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__u0 ( .ck(ispd_clk), .d(n_5358), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__u0 ( .ck(ispd_clk), .d(n_5509), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__u0 ( .ck(ispd_clk), .d(n_5511), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_5__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__u0 ( .ck(ispd_clk), .d(n_6980), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__u0 ( .ck(ispd_clk), .d(n_5470), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__u0 ( .ck(ispd_clk), .d(n_5356), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__u0 ( .ck(ispd_clk), .d(n_5539), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__u0 ( .ck(ispd_clk), .d(n_5534), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__u0 ( .ck(ispd_clk), .d(n_5248), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__u0 ( .ck(ispd_clk), .d(n_5351), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__u0 ( .ck(ispd_clk), .d(n_5531), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__u0 ( .ck(ispd_clk), .d(n_5349), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__u0 ( .ck(ispd_clk), .d(n_5483), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__u0 ( .ck(ispd_clk), .d(n_5347), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__u0 ( .ck(ispd_clk), .d(n_5716), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__u0 ( .ck(ispd_clk), .d(n_5345), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__u0 ( .ck(ispd_clk), .d(n_5521), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__u0 ( .ck(ispd_clk), .d(n_5342), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__u0 ( .ck(ispd_clk), .d(n_5528), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__u0 ( .ck(ispd_clk), .d(n_5499), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__u0 ( .ck(ispd_clk), .d(n_5260), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__u0 ( .ck(ispd_clk), .d(n_5339), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__u0 ( .ck(ispd_clk), .d(n_5240), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__u0 ( .ck(ispd_clk), .d(n_5242), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__u0 ( .ck(ispd_clk), .d(n_5253), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__u0 ( .ck(ispd_clk), .d(n_5427), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__u0 ( .ck(ispd_clk), .d(n_5446), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__u0 ( .ck(ispd_clk), .d(n_5467), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__u0 ( .ck(ispd_clk), .d(n_7130), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__u0 ( .ck(ispd_clk), .d(n_5335), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__u0 ( .ck(ispd_clk), .d(n_5537), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__u0 ( .ck(ispd_clk), .d(n_5489), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__u0 ( .ck(ispd_clk), .d(n_6135), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__36__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__u0 ( .ck(ispd_clk), .d(n_7694), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__u0 ( .ck(ispd_clk), .d(n_4930), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__u0 ( .ck(ispd_clk), .d(n_4625), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__u0 ( .ck(ispd_clk), .d(n_5503), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__u0 ( .ck(ispd_clk), .d(n_5330), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__u0 ( .ck(ispd_clk), .d(n_5517), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__u0 ( .ck(ispd_clk), .d(n_5513), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__u0 ( .ck(ispd_clk), .d(n_5523), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__u0 ( .ck(ispd_clk), .d(n_5327), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__u0 ( .ck(ispd_clk), .d(n_5543), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_6__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__u0 ( .ck(ispd_clk), .d(n_6969), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__0__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__u0 ( .ck(ispd_clk), .d(n_5277), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__10__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__u0 ( .ck(ispd_clk), .d(n_5285), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__11__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__u0 ( .ck(ispd_clk), .d(n_5325), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__12__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__u0 ( .ck(ispd_clk), .d(n_5438), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__13__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__u0 ( .ck(ispd_clk), .d(n_5431), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__14__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__u0 ( .ck(ispd_clk), .d(n_5454), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__15__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__u0 ( .ck(ispd_clk), .d(n_5320), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__16__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__u0 ( .ck(ispd_clk), .d(n_5272), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__17__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__u0 ( .ck(ispd_clk), .d(n_5293), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__18__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__u0 ( .ck(ispd_clk), .d(n_5235), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__19__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__u0 ( .ck(ispd_clk), .d(n_6973), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__1__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__u0 ( .ck(ispd_clk), .d(n_5246), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__20__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__u0 ( .ck(ispd_clk), .d(n_5486), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__21__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__u0 ( .ck(ispd_clk), .d(n_5495), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__22__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__u0 ( .ck(ispd_clk), .d(n_5313), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__23__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__u0 ( .ck(ispd_clk), .d(n_5519), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__24__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__u0 ( .ck(ispd_clk), .d(n_5526), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__25__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__u0 ( .ck(ispd_clk), .d(n_5435), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__26__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__u0 ( .ck(ispd_clk), .d(n_5452), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__27__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__u0 ( .ck(ispd_clk), .d(n_5311), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__28__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__u0 ( .ck(ispd_clk), .d(n_5456), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__29__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__u0 ( .ck(ispd_clk), .d(n_5507), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__2__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__u0 ( .ck(ispd_clk), .d(n_5476), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__30__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__u0 ( .ck(ispd_clk), .d(n_5541), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__31__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__u0 ( .ck(ispd_clk), .d(n_7132), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__32__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__u0 ( .ck(ispd_clk), .d(n_5444), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__33__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__u0 ( .ck(ispd_clk), .d(n_5465), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__34__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__u0 ( .ck(ispd_clk), .d(n_5515), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__35__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__u0 ( .ck(ispd_clk), .d(n_6125), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__36__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__u0 ( .ck(ispd_clk), .d(n_7687), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__37__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__u0 ( .ck(ispd_clk), .d(n_4934), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__38__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23474), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__39__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__u0 ( .ck(ispd_clk), .d(n_5251), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__3__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__u0 ( .ck(ispd_clk), .d(n_5472), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__4__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__u0 ( .ck(ispd_clk), .d(n_5263), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__5__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__u0 ( .ck(ispd_clk), .d(n_5474), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__6__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__u0 ( .ck(ispd_clk), .d(n_5269), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__7__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__u0 ( .ck(ispd_clk), .d(n_5279), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__8__Q) );
ms00f80 pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__u0 ( .ck(ispd_clk), .d(n_5283), .o(pci_target_unit_fifos_pciw_fifo_storage_mem_reg_7__9__Q) );
ms00f80 pci_target_unit_fifos_pciw_inTransactionCount_reg_0__u0 ( .ck(ispd_clk), .d(n_4797), .o(pci_target_unit_fifos_pciw_inTransactionCount_0_) );
ms00f80 pci_target_unit_fifos_pciw_inTransactionCount_reg_1__u0 ( .ck(ispd_clk), .d(n_5548), .o(pci_target_unit_fifos_pciw_inTransactionCount_reg_1__Q) );
in01s02 pci_target_unit_fifos_pciw_inTransactionCount_reg_1__u1 ( .a(pci_target_unit_fifos_pciw_inTransactionCount_reg_1__Q), .o(pci_target_unit_fifos_pciw_inTransactionCount_1_) );
ms00f80 pci_target_unit_fifos_pciw_outTransactionCount_reg_0__u0 ( .ck(ispd_clk), .d(n_13483), .o(pci_target_unit_fifos_pciw_outTransactionCount_reg_0__Q) );
ms00f80 pci_target_unit_fifos_pciw_outTransactionCount_reg_1__u0 ( .ck(ispd_clk), .d(n_13623), .o(pci_target_unit_fifos_pciw_outTransactionCount_reg_1__Q) );
in01s20 pci_target_unit_fifos_pciw_outTransactionCount_reg_1__u1 ( .a(pci_target_unit_fifos_pciw_outTransactionCount_reg_1__Q), .o(pci_target_unit_fifos_pciw_outTransactionCount_1_) );
ms00f80 pci_target_unit_fifos_wb_clk_inGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_wb_clk_sync_inGreyCount), .o(pci_target_unit_fifos_wb_clk_inGreyCount_0_) );
ms00f80 pci_target_unit_fifos_wb_clk_inGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(pci_target_unit_fifos_wb_clk_sync_inGreyCount_36), .o(pci_target_unit_fifos_wb_clk_inGreyCount_1_) );
ms00f80 pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_u0 ( .ck(ispd_clk), .d(n_4667), .o(pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_Q) );
in01m80 pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_u1 ( .a(pci_target_unit_pci_target_if_async_reset_as_pcir_flush_async_reset_data_out_reg_Q), .o(pci_target_unit_fifos_pcir_flush_in) );
ms00f80 pci_target_unit_pci_target_if_keep_desconnect_wo_data_set_reg_u0 ( .ck(ispd_clk), .d(n_12170), .o(pci_target_unit_pci_target_if_keep_desconnect_wo_data_set) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_0__u0 ( .ck(ispd_clk), .d(n_2603), .o(pci_target_unit_pci_target_if_norm_address_reg_0__Q) );
in01s06 pci_target_unit_pci_target_if_norm_address_reg_0__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_0__Q), .o(pci_target_unit_del_sync_addr_in) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_10__u0 ( .ck(ispd_clk), .d(n_2592), .o(pci_target_unit_del_sync_addr_in_213) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_11__u0 ( .ck(ispd_clk), .d(n_2595), .o(pci_target_unit_del_sync_addr_in_214) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_12__u0 ( .ck(ispd_clk), .d(n_2576), .o(pci_target_unit_del_sync_addr_in_215) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_13__u0 ( .ck(ispd_clk), .d(n_2593), .o(pci_target_unit_del_sync_addr_in_216) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_14__u0 ( .ck(ispd_clk), .d(n_2573), .o(pci_target_unit_del_sync_addr_in_217) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_15__u0 ( .ck(ispd_clk), .d(n_2574), .o(pci_target_unit_del_sync_addr_in_218) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_16__u0 ( .ck(ispd_clk), .d(n_2577), .o(pci_target_unit_del_sync_addr_in_219) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_17__u0 ( .ck(ispd_clk), .d(n_2570), .o(pci_target_unit_del_sync_addr_in_220) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_18__u0 ( .ck(ispd_clk), .d(n_2594), .o(pci_target_unit_del_sync_addr_in_221) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_19__u0 ( .ck(ispd_clk), .d(n_2588), .o(pci_target_unit_del_sync_addr_in_222) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_1__u0 ( .ck(ispd_clk), .d(n_2794), .o(pci_target_unit_pci_target_if_norm_address_reg_1__Q) );
in01s06 pci_target_unit_pci_target_if_norm_address_reg_1__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_1__Q), .o(pci_target_unit_del_sync_addr_in_204) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_20__u0 ( .ck(ispd_clk), .d(n_2571), .o(pci_target_unit_del_sync_addr_in_223) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_21__u0 ( .ck(ispd_clk), .d(n_2581), .o(pci_target_unit_del_sync_addr_in_224) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_22__u0 ( .ck(ispd_clk), .d(n_2590), .o(pci_target_unit_del_sync_addr_in_225) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_23__u0 ( .ck(ispd_clk), .d(n_2482), .o(pci_target_unit_del_sync_addr_in_226) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_24__u0 ( .ck(ispd_clk), .d(n_2572), .o(pci_target_unit_del_sync_addr_in_227) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_25__u0 ( .ck(ispd_clk), .d(n_2582), .o(pci_target_unit_del_sync_addr_in_228) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_26__u0 ( .ck(ispd_clk), .d(n_2583), .o(pci_target_unit_del_sync_addr_in_229) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_27__u0 ( .ck(ispd_clk), .d(n_2584), .o(pci_target_unit_del_sync_addr_in_230) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_28__u0 ( .ck(ispd_clk), .d(n_2585), .o(pci_target_unit_del_sync_addr_in_231) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_29__u0 ( .ck(ispd_clk), .d(n_2569), .o(pci_target_unit_del_sync_addr_in_232) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_2__u0 ( .ck(ispd_clk), .d(n_2792), .o(pci_target_unit_pci_target_if_norm_address_reg_2__Q) );
in01m20 pci_target_unit_pci_target_if_norm_address_reg_2__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_2__Q), .o(pci_target_unit_del_sync_addr_in_205) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_30__u0 ( .ck(ispd_clk), .d(n_2587), .o(pci_target_unit_del_sync_addr_in_233) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_31__u0 ( .ck(ispd_clk), .d(n_2586), .o(pci_target_unit_del_sync_addr_in_234) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_3__u0 ( .ck(ispd_clk), .d(n_2789), .o(pci_target_unit_pci_target_if_norm_address_reg_3__Q) );
in01m03 pci_target_unit_pci_target_if_norm_address_reg_3__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_3__Q), .o(pci_target_unit_del_sync_addr_in_206) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_4__u0 ( .ck(ispd_clk), .d(n_2734), .o(pci_target_unit_pci_target_if_norm_address_reg_4__Q) );
in01m20 pci_target_unit_pci_target_if_norm_address_reg_4__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_4__Q), .o(pci_target_unit_del_sync_addr_in_207) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_5__u0 ( .ck(ispd_clk), .d(n_2605), .o(pci_target_unit_pci_target_if_norm_address_reg_5__Q) );
in01m03 pci_target_unit_pci_target_if_norm_address_reg_5__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_5__Q), .o(pci_target_unit_del_sync_addr_in_208) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_6__u0 ( .ck(ispd_clk), .d(n_2787), .o(pci_target_unit_pci_target_if_norm_address_reg_6__Q) );
in01m03 pci_target_unit_pci_target_if_norm_address_reg_6__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_6__Q), .o(pci_target_unit_del_sync_addr_in_209) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_7__u0 ( .ck(ispd_clk), .d(n_2608), .o(pci_target_unit_pci_target_if_norm_address_reg_7__Q) );
in01m20 pci_target_unit_pci_target_if_norm_address_reg_7__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_7__Q), .o(pci_target_unit_del_sync_addr_in_210) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_8__u0 ( .ck(ispd_clk), .d(n_2611), .o(pci_target_unit_pci_target_if_norm_address_reg_8__Q) );
in01m20 pci_target_unit_pci_target_if_norm_address_reg_8__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_8__Q), .o(pci_target_unit_del_sync_addr_in_211) );
ms00f80 pci_target_unit_pci_target_if_norm_address_reg_9__u0 ( .ck(ispd_clk), .d(n_2613), .o(pci_target_unit_pci_target_if_norm_address_reg_9__Q) );
in01m20 pci_target_unit_pci_target_if_norm_address_reg_9__u1 ( .a(pci_target_unit_pci_target_if_norm_address_reg_9__Q), .o(pci_target_unit_del_sync_addr_in_212) );
ms00f80 pci_target_unit_pci_target_if_norm_bc_reg_0__u0 ( .ck(ispd_clk), .d(n_3220), .o(pci_target_unit_del_sync_bc_in) );
ms00f80 pci_target_unit_pci_target_if_norm_bc_reg_1__u0 ( .ck(ispd_clk), .d(n_2793), .o(pci_target_unit_del_sync_bc_in_201) );
ms00f80 pci_target_unit_pci_target_if_norm_bc_reg_2__u0 ( .ck(ispd_clk), .d(n_2575), .o(pci_target_unit_del_sync_bc_in_202) );
ms00f80 pci_target_unit_pci_target_if_norm_bc_reg_3__u0 ( .ck(ispd_clk), .d(n_2579), .o(pci_target_unit_del_sync_bc_in_203) );
ms00f80 pci_target_unit_pci_target_if_norm_prf_en_reg_u0 ( .ck(ispd_clk), .d(n_8659), .o(pci_target_unit_pci_target_if_norm_prf_en) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_reg_1__u0 ( .ck(ispd_clk), .d(n_13146), .o(pci_target_unit_pci_target_if_pcir_fifo_ctrl_reg_77) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__u0 ( .ck(ispd_clk), .d(n_12980), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_0__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__u0 ( .ck(ispd_clk), .d(n_12978), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_10__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__u0 ( .ck(ispd_clk), .d(n_12976), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_11__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__u0 ( .ck(ispd_clk), .d(n_12974), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_12__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__u0 ( .ck(ispd_clk), .d(n_12972), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_13__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__u0 ( .ck(ispd_clk), .d(n_12970), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_14__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__u0 ( .ck(ispd_clk), .d(n_13097), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_15__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__u0 ( .ck(ispd_clk), .d(n_12968), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_16__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__u0 ( .ck(ispd_clk), .d(n_12966), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_17__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__u0 ( .ck(ispd_clk), .d(n_13095), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_18__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__u0 ( .ck(ispd_clk), .d(n_13094), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_19__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__u0 ( .ck(ispd_clk), .d(n_13093), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_1__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__u0 ( .ck(ispd_clk), .d(n_13091), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_20__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__u0 ( .ck(ispd_clk), .d(n_13090), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_21__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__u0 ( .ck(ispd_clk), .d(n_13089), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_22__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__u0 ( .ck(ispd_clk), .d(n_13088), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_23__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__u0 ( .ck(ispd_clk), .d(n_13087), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_24__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__u0 ( .ck(ispd_clk), .d(n_13125), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_25__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__u0 ( .ck(ispd_clk), .d(n_13086), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_26__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__u0 ( .ck(ispd_clk), .d(n_13085), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_27__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__u0 ( .ck(ispd_clk), .d(n_13084), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_28__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__u0 ( .ck(ispd_clk), .d(n_13083), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_29__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__u0 ( .ck(ispd_clk), .d(n_13082), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_2__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__u0 ( .ck(ispd_clk), .d(n_13081), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_30__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__u0 ( .ck(ispd_clk), .d(n_13080), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_31__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__u0 ( .ck(ispd_clk), .d(n_13079), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_3__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__u0 ( .ck(ispd_clk), .d(n_13078), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_4__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__u0 ( .ck(ispd_clk), .d(n_13077), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_5__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__u0 ( .ck(ispd_clk), .d(n_13076), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_6__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__u0 ( .ck(ispd_clk), .d(n_13123), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_7__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__u0 ( .ck(ispd_clk), .d(n_13075), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_8__Q) );
ms00f80 pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__u0 ( .ck(ispd_clk), .d(n_13074), .o(pci_target_unit_pci_target_if_pcir_fifo_data_reg_reg_9__Q) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_2776), .o(pci_target_unit_fifos_pciw_addr_data_in) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_10__u0 ( .ck(ispd_clk), .d(n_2519), .o(pci_target_unit_fifos_pciw_addr_data_in_130) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_11__u0 ( .ck(ispd_clk), .d(n_2517), .o(pci_target_unit_fifos_pciw_addr_data_in_131) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_12__u0 ( .ck(ispd_clk), .d(n_2546), .o(pci_target_unit_fifos_pciw_addr_data_in_132) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_13__u0 ( .ck(ispd_clk), .d(n_2534), .o(pci_target_unit_fifos_pciw_addr_data_in_133) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_14__u0 ( .ck(ispd_clk), .d(n_2496), .o(pci_target_unit_fifos_pciw_addr_data_in_134) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_15__u0 ( .ck(ispd_clk), .d(n_2498), .o(pci_target_unit_fifos_pciw_addr_data_in_135) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_16__u0 ( .ck(ispd_clk), .d(n_2537), .o(pci_target_unit_fifos_pciw_addr_data_in_136) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_17__u0 ( .ck(ispd_clk), .d(n_2536), .o(pci_target_unit_fifos_pciw_addr_data_in_137) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_18__u0 ( .ck(ispd_clk), .d(n_2530), .o(pci_target_unit_fifos_pciw_addr_data_in_138) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_19__u0 ( .ck(ispd_clk), .d(n_2528), .o(pci_target_unit_fifos_pciw_addr_data_in_139) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_1__u0 ( .ck(ispd_clk), .d(n_2973), .o(pci_target_unit_fifos_pciw_addr_data_in_121) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_20__u0 ( .ck(ispd_clk), .d(n_2540), .o(pci_target_unit_fifos_pciw_addr_data_in_140) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_21__u0 ( .ck(ispd_clk), .d(n_2531), .o(pci_target_unit_fifos_pciw_addr_data_in_141) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_22__u0 ( .ck(ispd_clk), .d(n_2514), .o(pci_target_unit_fifos_pciw_addr_data_in_142) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_23__u0 ( .ck(ispd_clk), .d(n_2539), .o(pci_target_unit_fifos_pciw_addr_data_in_143) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_24__u0 ( .ck(ispd_clk), .d(n_2502), .o(pci_target_unit_fifos_pciw_addr_data_in_144) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_25__u0 ( .ck(ispd_clk), .d(n_2522), .o(pci_target_unit_fifos_pciw_addr_data_in_145) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_26__u0 ( .ck(ispd_clk), .d(n_2533), .o(pci_target_unit_fifos_pciw_addr_data_in_146) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_27__u0 ( .ck(ispd_clk), .d(n_2543), .o(pci_target_unit_fifos_pciw_addr_data_in_147) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_28__u0 ( .ck(ispd_clk), .d(n_2518), .o(pci_target_unit_fifos_pciw_addr_data_in_148) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_29__u0 ( .ck(ispd_clk), .d(n_2505), .o(pci_target_unit_fifos_pciw_addr_data_in_149) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2516), .o(pci_target_unit_fifos_pciw_addr_data_in_122) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_30__u0 ( .ck(ispd_clk), .d(n_2510), .o(pci_target_unit_fifos_pciw_addr_data_in_150) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_31__u0 ( .ck(ispd_clk), .d(n_2497), .o(pci_target_unit_fifos_pciw_addr_data_in_151) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2500), .o(pci_target_unit_fifos_pciw_addr_data_in_123) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_4__u0 ( .ck(ispd_clk), .d(n_2527), .o(pci_target_unit_fifos_pciw_addr_data_in_124) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_5__u0 ( .ck(ispd_clk), .d(n_2545), .o(pci_target_unit_fifos_pciw_addr_data_in_125) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_6__u0 ( .ck(ispd_clk), .d(n_2513), .o(pci_target_unit_fifos_pciw_addr_data_in_126) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_7__u0 ( .ck(ispd_clk), .d(n_2542), .o(pci_target_unit_fifos_pciw_addr_data_in_127) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_8__u0 ( .ck(ispd_clk), .d(n_2508), .o(pci_target_unit_fifos_pciw_addr_data_in_128) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_addr_data_out_reg_9__u0 ( .ck(ispd_clk), .d(n_2504), .o(pci_target_unit_fifos_pciw_addr_data_in_129) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg_0__u0 ( .ck(ispd_clk), .d(n_3000), .o(pci_target_unit_fifos_pciw_cbe_in) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23476), .o(pci_target_unit_fifos_pciw_cbe_in_152) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg_2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23478), .o(pci_target_unit_fifos_pciw_cbe_in_153) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_cbe_out_reg_3__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23480), .o(pci_target_unit_fifos_pciw_cbe_in_154) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__u0 ( .ck(ispd_clk), .d(FE_OFN793_n_2547), .o(pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__Q) );
in01s03 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__u1 ( .a(pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_0__Q), .o(pci_target_unit_fifos_pciw_control_in) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_1__u0 ( .ck(ispd_clk), .d(n_4142), .o(pci_target_unit_fifos_pciw_control_in_155) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_2__u0 ( .ck(ispd_clk), .d(n_2729), .o(pci_target_unit_fifos_pciw_control_in_156) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_control_out_reg_3__u0 ( .ck(ispd_clk), .d(n_2031), .o(pci_target_unit_fifos_pciw_control_in_157) );
ms00f80 pci_target_unit_pci_target_if_pciw_fifo_wenable_out_reg_u0 ( .ck(ispd_clk), .d(n_8566), .o(pci_target_unit_fifos_pciw_wenable_in) );
ms00f80 pci_target_unit_pci_target_if_same_read_reg_reg_u0 ( .ck(ispd_clk), .d(n_5640), .o(pci_target_unit_pci_target_if_same_read_reg) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_0__u0 ( .ck(ispd_clk), .d(n_2602), .o(conf_w_addr_in) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_1__u0 ( .ck(ispd_clk), .d(n_2780), .o(conf_w_addr_in_931) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_2__u0 ( .ck(ispd_clk), .d(n_4214), .o(conf_w_addr_in_932) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_3__u0 ( .ck(ispd_clk), .d(n_3216), .o(conf_w_addr_in_933) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_4__u0 ( .ck(ispd_clk), .d(n_2781), .o(n_2078) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_5__u0 ( .ck(ispd_clk), .d(n_2782), .o(conf_w_addr_in_935) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_6__u0 ( .ck(ispd_clk), .d(n_2784), .o(n_15998) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_7__u0 ( .ck(ispd_clk), .d(n_2745), .o(conf_w_addr_in_937) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_8__u0 ( .ck(ispd_clk), .d(n_2786), .o(conf_w_addr_in_938) );
ms00f80 pci_target_unit_pci_target_if_strd_address_reg_9__u0 ( .ck(ispd_clk), .d(n_2785), .o(conf_w_addr_in_939) );
ms00f80 pci_target_unit_pci_target_if_target_rd_reg_u0 ( .ck(ispd_clk), .d(n_3380), .o(pci_target_unit_pci_target_if_target_rd_completed) );
ms00f80 pci_target_unit_pci_target_sm_backoff_reg_u0 ( .ck(ispd_clk), .d(n_14630), .o(pci_target_unit_pci_target_sm_backoff) );
ms00f80 pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_u0 ( .ck(ispd_clk), .d(output_backup_trdy_out_reg_Q), .o(pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_Q) );
in01f80 pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_u1 ( .a(pci_target_unit_pci_target_sm_bckp_trdy_reg_reg_Q), .o(n_2597) );
ms00f80 pci_target_unit_pci_target_sm_c_state_reg_0__u0 ( .ck(ispd_clk), .d(n_9180), .o(n_1628) );
ms00f80 pci_target_unit_pci_target_sm_c_state_reg_1__u0 ( .ck(ispd_clk), .d(n_9179), .o(pci_target_unit_pci_target_sm_n_2) );
ms00f80 pci_target_unit_pci_target_sm_c_state_reg_2__u0 ( .ck(ispd_clk), .d(n_9176), .o(pci_target_unit_pci_target_sm_n_3) );
ms00f80 pci_target_unit_pci_target_sm_cnf_progress_reg_u0 ( .ck(ispd_clk), .d(n_2946), .o(pci_target_unit_pci_target_sm_cnf_progress) );
ms00f80 pci_target_unit_pci_target_sm_master_will_request_read_reg_u0 ( .ck(ispd_clk), .d(n_8528), .o(pci_target_unit_pci_target_sm_master_will_request_read) );
ms00f80 pci_target_unit_pci_target_sm_norm_access_to_conf_reg_reg_u0 ( .ck(ispd_clk), .d(n_8574), .o(n_2314) );
ms00f80 pci_target_unit_pci_target_sm_previous_frame_reg_u0 ( .ck(ispd_clk), .d(n_15302), .o(pci_target_unit_pci_target_sm_previous_frame) );
ms00f80 pci_target_unit_pci_target_sm_rd_from_fifo_reg_u0 ( .ck(ispd_clk), .d(n_3364), .o(pci_target_unit_pci_target_sm_rd_from_fifo) );
ms00f80 pci_target_unit_pci_target_sm_rd_progress_reg_u0 ( .ck(ispd_clk), .d(n_8688), .o(pci_target_unit_pci_target_sm_rd_progress) );
ms00f80 pci_target_unit_pci_target_sm_rd_request_reg_u0 ( .ck(ispd_clk), .d(n_8687), .o(pci_target_unit_pci_target_sm_rd_request_reg_Q) );
in01s01 pci_target_unit_pci_target_sm_rd_request_reg_u1 ( .a(pci_target_unit_pci_target_sm_rd_request_reg_Q), .o(pci_target_unit_pci_target_sm_rd_request) );
ms00f80 pci_target_unit_pci_target_sm_read_completed_reg_reg_u0 ( .ck(ispd_clk), .d(n_2337), .o(pci_target_unit_pci_target_sm_read_completed_reg_reg_Q) );
in01f40 pci_target_unit_pci_target_sm_read_completed_reg_reg_u1 ( .a(pci_target_unit_pci_target_sm_read_completed_reg_reg_Q), .o(pci_target_unit_pci_target_sm_read_completed_reg) );
ms00f80 pci_target_unit_pci_target_sm_rw_cbe0_reg_u0 ( .ck(ispd_clk), .d(n_3219), .o(n_978) );
ms00f80 pci_target_unit_pci_target_sm_same_read_reg_reg_u0 ( .ck(ispd_clk), .d(n_4895), .o(pci_target_unit_pci_target_sm_same_read_reg) );
ms00f80 pci_target_unit_pci_target_sm_state_backoff_reg_reg_u0 ( .ck(ispd_clk), .d(n_2140), .o(pci_target_unit_pci_target_sm_state_backoff_reg_reg_Q) );
ms00f80 pci_target_unit_pci_target_sm_state_transfere_reg_reg_u0 ( .ck(ispd_clk), .d(n_13817), .o(pci_target_unit_pci_target_sm_state_transfere_reg_reg_Q) );
in01f80 pci_target_unit_pci_target_sm_state_transfere_reg_reg_u1 ( .a(pci_target_unit_pci_target_sm_state_transfere_reg_reg_Q), .o(pci_target_unit_pci_target_sm_state_transfere_reg) );
ms00f80 pci_target_unit_pci_target_sm_wr_progress_reg_u0 ( .ck(ispd_clk), .d(n_8573), .o(pci_target_unit_pci_target_sm_wr_progress) );
ms00f80 pci_target_unit_pci_target_sm_wr_to_fifo_reg_u0 ( .ck(ispd_clk), .d(n_3499), .o(pci_target_unit_pci_target_sm_wr_to_fifo) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_0__u0 ( .ck(ispd_clk), .d(n_14804), .o(wbm_adr_o_0_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_10__u0 ( .ck(ispd_clk), .d(n_14813), .o(wbm_adr_o_10_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_11__u0 ( .ck(ispd_clk), .d(n_14812), .o(wbm_adr_o_11_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_12__u0 ( .ck(ispd_clk), .d(n_14811), .o(wbm_adr_o_12_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_13__u0 ( .ck(ispd_clk), .d(n_14810), .o(wbm_adr_o_13_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_14__u0 ( .ck(ispd_clk), .d(n_14847), .o(wbm_adr_o_14_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_15__u0 ( .ck(ispd_clk), .d(n_14808), .o(wbm_adr_o_15_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_16__u0 ( .ck(ispd_clk), .d(n_14848), .o(wbm_adr_o_16_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_17__u0 ( .ck(ispd_clk), .d(n_14828), .o(wbm_adr_o_17_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_18__u0 ( .ck(ispd_clk), .d(n_14803), .o(wbm_adr_o_18_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_19__u0 ( .ck(ispd_clk), .d(n_14826), .o(wbm_adr_o_19_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_1__u0 ( .ck(ispd_clk), .d(n_14805), .o(wbm_adr_o_1_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_20__u0 ( .ck(ispd_clk), .d(n_14825), .o(wbm_adr_o_20_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_21__u0 ( .ck(ispd_clk), .d(n_14818), .o(wbm_adr_o_21_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_22__u0 ( .ck(ispd_clk), .d(n_14824), .o(wbm_adr_o_22_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_23__u0 ( .ck(ispd_clk), .d(n_14846), .o(wbm_adr_o_23_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_24__u0 ( .ck(ispd_clk), .d(n_14822), .o(wbm_adr_o_24_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_25__u0 ( .ck(ispd_clk), .d(n_14821), .o(wbm_adr_o_25_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_26__u0 ( .ck(ispd_clk), .d(n_14845), .o(wbm_adr_o_26_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_27__u0 ( .ck(ispd_clk), .d(n_14819), .o(wbm_adr_o_27_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_28__u0 ( .ck(ispd_clk), .d(n_14815), .o(wbm_adr_o_28_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_29__u0 ( .ck(ispd_clk), .d(n_14817), .o(wbm_adr_o_29_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_2__u0 ( .ck(ispd_clk), .d(n_14844), .o(wbm_adr_o_2_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_30__u0 ( .ck(ispd_clk), .d(n_14816), .o(wbm_adr_o_30_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_31__u0 ( .ck(ispd_clk), .d(n_14814), .o(wbm_adr_o_31_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_3__u0 ( .ck(ispd_clk), .d(n_14842), .o(wbm_adr_o_3_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_4__u0 ( .ck(ispd_clk), .d(n_14841), .o(wbm_adr_o_4_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_5__u0 ( .ck(ispd_clk), .d(n_14840), .o(wbm_adr_o_5_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_6__u0 ( .ck(ispd_clk), .d(n_14838), .o(wbm_adr_o_6_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_7__u0 ( .ck(ispd_clk), .d(n_14807), .o(wbm_adr_o_7_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_8__u0 ( .ck(ispd_clk), .d(n_14836), .o(wbm_adr_o_8_) );
ms00f80 pci_target_unit_wishbone_master_addr_cnt_out_reg_9__u0 ( .ck(ispd_clk), .d(n_14834), .o(wbm_adr_o_9_) );
ms00f80 pci_target_unit_wishbone_master_addr_into_cnt_reg_reg_u0 ( .ck(ispd_clk), .d(n_8757), .o(pci_target_unit_wishbone_master_addr_into_cnt_reg) );
ms00f80 pci_target_unit_wishbone_master_bc_register_reg_0__u0 ( .ck(ispd_clk), .d(n_14687), .o(pci_target_unit_wishbone_master_bc_register_reg_0__Q) );
ms00f80 pci_target_unit_wishbone_master_bc_register_reg_1__u0 ( .ck(ispd_clk), .d(n_14686), .o(pci_target_unit_wishbone_master_bc_register_reg_1__Q) );
ms00f80 pci_target_unit_wishbone_master_bc_register_reg_2__u0 ( .ck(ispd_clk), .d(n_14685), .o(pci_target_unit_wishbone_master_bc_register_reg_2__Q) );
ms00f80 pci_target_unit_wishbone_master_bc_register_reg_3__u0 ( .ck(ispd_clk), .d(n_14683), .o(pci_target_unit_wishbone_master_bc_register_reg_3__Q) );
ms00f80 pci_target_unit_wishbone_master_burst_chopped_delayed_reg_u0 ( .ck(ispd_clk), .d(pci_target_unit_wishbone_master_burst_chopped), .o(pci_target_unit_wishbone_master_burst_chopped_delayed_reg_Q) );
in01f40 pci_target_unit_wishbone_master_burst_chopped_delayed_reg_u1 ( .a(pci_target_unit_wishbone_master_burst_chopped_delayed_reg_Q), .o(pci_target_unit_wishbone_master_burst_chopped_delayed) );
ms00f80 pci_target_unit_wishbone_master_burst_chopped_reg_u0 ( .ck(ispd_clk), .d(n_14694), .o(pci_target_unit_wishbone_master_burst_chopped) );
ms00f80 pci_target_unit_wishbone_master_c_state_reg_0__u0 ( .ck(ispd_clk), .d(n_16167), .o(pci_target_unit_wishbone_master_c_state_0_) );
ms00f80 pci_target_unit_wishbone_master_c_state_reg_1__u0 ( .ck(ispd_clk), .d(n_8452), .o(pci_target_unit_wishbone_master_c_state_1_) );
ms00f80 pci_target_unit_wishbone_master_c_state_reg_2__u0 ( .ck(ispd_clk), .d(n_15188), .o(pci_target_unit_wishbone_master_c_state_2_) );
ms00f80 pci_target_unit_wishbone_master_first_data_is_burst_reg_reg_u0 ( .ck(ispd_clk), .d(n_10787), .o(pci_target_unit_wishbone_master_first_data_is_burst_reg) );
ms00f80 pci_target_unit_wishbone_master_first_wb_data_access_reg_u0 ( .ck(ispd_clk), .d(n_13789), .o(pci_target_unit_wishbone_master_first_wb_data_access) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_control_out_reg_1__u0 ( .ck(ispd_clk), .d(n_3223), .o(pci_target_unit_fifos_pcir_control_in_192) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23482), .o(pci_target_unit_fifos_pcir_data_in) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_10__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23484), .o(pci_target_unit_fifos_pcir_data_in_167) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_11__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23486), .o(pci_target_unit_fifos_pcir_data_in_168) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_12__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23488), .o(pci_target_unit_fifos_pcir_data_in_169) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_13__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23490), .o(TIMEBOOST_net_21127) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_14__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23492), .o(pci_target_unit_fifos_pcir_data_in_171) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_15__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23494), .o(pci_target_unit_fifos_pcir_data_in_172) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_16__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23496), .o(pci_target_unit_fifos_pcir_data_in_173) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_17__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23498), .o(pci_target_unit_fifos_pcir_data_in_174) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_18__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23500), .o(pci_target_unit_fifos_pcir_data_in_175) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_19__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23502), .o(pci_target_unit_fifos_pcir_data_in_176) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23504), .o(pci_target_unit_fifos_pcir_data_in_158) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_20__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23506), .o(pci_target_unit_fifos_pcir_data_in_177) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_21__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23508), .o(pci_target_unit_fifos_pcir_data_in_178) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_22__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23510), .o(pci_target_unit_fifos_pcir_data_in_179) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_23__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23512), .o(pci_target_unit_fifos_pcir_data_in_180) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_24__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23514), .o(pci_target_unit_fifos_pcir_data_in_181) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_25__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23516), .o(TIMEBOOST_net_21207) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_26__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23518), .o(pci_target_unit_fifos_pcir_data_in_183) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_27__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23520), .o(pci_target_unit_fifos_pcir_data_in_184) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_28__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23522), .o(pci_target_unit_fifos_pcir_data_in_185) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_29__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23524), .o(TIMEBOOST_net_21119) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23526), .o(pci_target_unit_fifos_pcir_data_in_159) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_30__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23528), .o(pci_target_unit_fifos_pcir_data_in_187) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_31__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23530), .o(pci_target_unit_fifos_pcir_data_in_188) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_3__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23532), .o(pci_target_unit_fifos_pcir_data_in_160) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_4__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23534), .o(pci_target_unit_fifos_pcir_data_in_161) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_5__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23536), .o(TIMEBOOST_net_21161) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_6__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23538), .o(pci_target_unit_fifos_pcir_data_in_163) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_7__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23540), .o(pci_target_unit_fifos_pcir_data_in_164) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_8__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23542), .o(pci_target_unit_fifos_pcir_data_in_165) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_data_out_reg_9__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23544), .o(pci_target_unit_fifos_pcir_data_in_166) );
ms00f80 pci_target_unit_wishbone_master_pcir_fifo_wenable_out_reg_u0 ( .ck(ispd_clk), .d(n_3224), .o(pci_target_unit_fifos_pcir_wenable_in) );
ms00f80 pci_target_unit_wishbone_master_read_bound_reg_u0 ( .ck(ispd_clk), .d(n_7401), .o(pci_target_unit_wishbone_master_read_bound) );
ms00f80 pci_target_unit_wishbone_master_read_count_reg_0__u0 ( .ck(ispd_clk), .d(n_7575), .o(pci_target_unit_wishbone_master_read_count_0_) );
ms00f80 pci_target_unit_wishbone_master_read_count_reg_1__u0 ( .ck(ispd_clk), .d(n_7609), .o(pci_target_unit_wishbone_master_read_count_1_) );
ms00f80 pci_target_unit_wishbone_master_read_count_reg_2__u0 ( .ck(ispd_clk), .d(n_7791), .o(pci_target_unit_wishbone_master_read_count_reg_2__Q) );
ms00f80 pci_target_unit_wishbone_master_reset_rty_cnt_reg_u0 ( .ck(ispd_clk), .d(n_8494), .o(pci_target_unit_wishbone_master_reset_rty_cnt_reg_Q) );
in01s10 pci_target_unit_wishbone_master_reset_rty_cnt_reg_u1 ( .a(pci_target_unit_wishbone_master_reset_rty_cnt_reg_Q), .o(pci_target_unit_wishbone_master_reset_rty_cnt) );
ms00f80 pci_target_unit_wishbone_master_retried_reg_u0 ( .ck(ispd_clk), .d(n_3268), .o(pci_target_unit_wishbone_master_retried) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_0__u0 ( .ck(ispd_clk), .d(n_8818), .o(pci_target_unit_wishbone_master_rty_counter_0_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_1__u0 ( .ck(ispd_clk), .d(n_8721), .o(pci_target_unit_wishbone_master_rty_counter_1_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_2__u0 ( .ck(ispd_clk), .d(n_8726), .o(n_1263) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_3__u0 ( .ck(ispd_clk), .d(n_8725), .o(pci_target_unit_wishbone_master_rty_counter_3_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_4__u0 ( .ck(ispd_clk), .d(n_8724), .o(pci_target_unit_wishbone_master_rty_counter_4_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_5__u0 ( .ck(ispd_clk), .d(n_8734), .o(pci_target_unit_wishbone_master_rty_counter_5_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_6__u0 ( .ck(ispd_clk), .d(n_8733), .o(pci_target_unit_wishbone_master_rty_counter_6_) );
ms00f80 pci_target_unit_wishbone_master_rty_counter_reg_7__u0 ( .ck(ispd_clk), .d(n_8731), .o(pci_target_unit_wishbone_master_rty_counter_7_) );
ms00f80 pci_target_unit_wishbone_master_w_attempt_reg_u0 ( .ck(ispd_clk), .d(n_8565), .o(n_16501) );
ms00f80 pci_target_unit_wishbone_master_wb_cti_o_reg_0__u0 ( .ck(ispd_clk), .d(n_14904), .o(wbm_cti_o_0_) );
ms00f80 pci_target_unit_wishbone_master_wb_cti_o_reg_1__u0 ( .ck(ispd_clk), .d(n_14629), .o(wbm_cti_o_1_) );
ms00f80 pci_target_unit_wishbone_master_wb_cti_o_reg_2__u0 ( .ck(ispd_clk), .d(n_14903), .o(wbm_cti_o_2_) );
ms00f80 pci_target_unit_wishbone_master_wb_cyc_o_reg_u0 ( .ck(ispd_clk), .d(n_13624), .o(pci_target_unit_wishbone_master_wb_cyc_o_reg_Q) );
in01f20 pci_target_unit_wishbone_master_wb_cyc_o_reg_u1 ( .a(pci_target_unit_wishbone_master_wb_cyc_o_reg_Q), .o(wbm_cyc_o_1378) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_0__u0 ( .ck(ispd_clk), .d(n_14887), .o(wbm_dat_o_0_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_10__u0 ( .ck(ispd_clk), .d(n_15197), .o(wbm_dat_o_10_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_11__u0 ( .ck(ispd_clk), .d(n_14885), .o(wbm_dat_o_11_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_12__u0 ( .ck(ispd_clk), .d(n_14884), .o(wbm_dat_o_12_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_13__u0 ( .ck(ispd_clk), .d(n_14883), .o(wbm_dat_o_13_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_14__u0 ( .ck(ispd_clk), .d(n_14881), .o(wbm_dat_o_14_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_15__u0 ( .ck(ispd_clk), .d(n_14851), .o(wbm_dat_o_15_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_16__u0 ( .ck(ispd_clk), .d(n_14879), .o(wbm_dat_o_16_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_17__u0 ( .ck(ispd_clk), .d(n_14880), .o(wbm_dat_o_17_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_18__u0 ( .ck(ispd_clk), .d(n_14850), .o(wbm_dat_o_18_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_19__u0 ( .ck(ispd_clk), .d(n_14877), .o(wbm_dat_o_19_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_1__u0 ( .ck(ispd_clk), .d(n_14875), .o(wbm_dat_o_1_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_20__u0 ( .ck(ispd_clk), .d(n_14873), .o(wbm_dat_o_20_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_21__u0 ( .ck(ispd_clk), .d(n_14871), .o(wbm_dat_o_21_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_22__u0 ( .ck(ispd_clk), .d(n_16304), .o(wbm_dat_o_22_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_23__u0 ( .ck(ispd_clk), .d(n_14869), .o(wbm_dat_o_23_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_24__u0 ( .ck(ispd_clk), .d(n_14867), .o(wbm_dat_o_24_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_25__u0 ( .ck(ispd_clk), .d(n_14866), .o(wbm_dat_o_25_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_26__u0 ( .ck(ispd_clk), .d(n_14865), .o(wbm_dat_o_26_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_27__u0 ( .ck(ispd_clk), .d(n_14863), .o(wbm_dat_o_27_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_28__u0 ( .ck(ispd_clk), .d(n_14864), .o(wbm_dat_o_28_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_29__u0 ( .ck(ispd_clk), .d(n_14862), .o(wbm_dat_o_29_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_2__u0 ( .ck(ispd_clk), .d(n_14861), .o(wbm_dat_o_2_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_30__u0 ( .ck(ispd_clk), .d(n_14860), .o(wbm_dat_o_30_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_31__u0 ( .ck(ispd_clk), .d(n_14856), .o(wbm_dat_o_31_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_3__u0 ( .ck(ispd_clk), .d(n_14859), .o(wbm_dat_o_3_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_4__u0 ( .ck(ispd_clk), .d(n_14858), .o(wbm_dat_o_4_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_5__u0 ( .ck(ispd_clk), .d(n_14855), .o(wbm_dat_o_5_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_6__u0 ( .ck(ispd_clk), .d(n_14854), .o(wbm_dat_o_6_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_7__u0 ( .ck(ispd_clk), .d(n_14849), .o(wbm_dat_o_7_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_8__u0 ( .ck(ispd_clk), .d(n_14853), .o(wbm_dat_o_8_) );
ms00f80 pci_target_unit_wishbone_master_wb_dat_o_reg_9__u0 ( .ck(ispd_clk), .d(n_14852), .o(wbm_dat_o_9_) );
ms00f80 pci_target_unit_wishbone_master_wb_read_done_out_reg_u0 ( .ck(ispd_clk), .d(n_4896), .o(pci_target_unit_del_sync_comp_in) );
ms00f80 pci_target_unit_wishbone_master_wb_sel_o_reg_0__u0 ( .ck(ispd_clk), .d(n_14897), .o(wbm_sel_o_0_) );
ms00f80 pci_target_unit_wishbone_master_wb_sel_o_reg_1__u0 ( .ck(ispd_clk), .d(n_14894), .o(wbm_sel_o_1_) );
ms00f80 pci_target_unit_wishbone_master_wb_sel_o_reg_2__u0 ( .ck(ispd_clk), .d(n_14896), .o(wbm_sel_o_2_) );
ms00f80 pci_target_unit_wishbone_master_wb_sel_o_reg_3__u0 ( .ck(ispd_clk), .d(n_14893), .o(wbm_sel_o_3_) );
ms00f80 pci_target_unit_wishbone_master_wb_stb_o_reg_u0 ( .ck(ispd_clk), .d(n_13624), .o(wbm_stb_o) );
ms00f80 pci_target_unit_wishbone_master_wb_we_o_reg_u0 ( .ck(ispd_clk), .d(n_13481), .o(wbm_we_o) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_0__u0 ( .ck(ispd_clk), .d(n_9402), .o(wishbone_slave_unit_del_sync_addr_out_reg_0__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_10__u0 ( .ck(ispd_clk), .d(n_9400), .o(wishbone_slave_unit_del_sync_addr_out_reg_10__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_11__u0 ( .ck(ispd_clk), .d(n_9398), .o(wishbone_slave_unit_del_sync_addr_out_reg_11__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_12__u0 ( .ck(ispd_clk), .d(n_8989), .o(wishbone_slave_unit_del_sync_addr_out_reg_12__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_13__u0 ( .ck(ispd_clk), .d(n_9396), .o(wishbone_slave_unit_del_sync_addr_out_reg_13__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_14__u0 ( .ck(ispd_clk), .d(n_8986), .o(wishbone_slave_unit_del_sync_addr_out_reg_14__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_15__u0 ( .ck(ispd_clk), .d(n_9393), .o(wishbone_slave_unit_del_sync_addr_out_reg_15__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_16__u0 ( .ck(ispd_clk), .d(n_9391), .o(wishbone_slave_unit_del_sync_addr_out_reg_16__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_17__u0 ( .ck(ispd_clk), .d(n_9389), .o(wishbone_slave_unit_del_sync_addr_out_reg_17__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_18__u0 ( .ck(ispd_clk), .d(n_9387), .o(wishbone_slave_unit_del_sync_addr_out_reg_18__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_19__u0 ( .ck(ispd_clk), .d(n_9385), .o(wishbone_slave_unit_del_sync_addr_out_reg_19__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_1__u0 ( .ck(ispd_clk), .d(n_9383), .o(wishbone_slave_unit_del_sync_addr_out_reg_1__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_20__u0 ( .ck(ispd_clk), .d(n_9381), .o(wishbone_slave_unit_del_sync_addr_out_reg_20__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_21__u0 ( .ck(ispd_clk), .d(n_9379), .o(wishbone_slave_unit_del_sync_addr_out_reg_21__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_22__u0 ( .ck(ispd_clk), .d(n_8983), .o(wishbone_slave_unit_del_sync_addr_out_reg_22__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_23__u0 ( .ck(ispd_clk), .d(n_9377), .o(wishbone_slave_unit_del_sync_addr_out_reg_23__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_24__u0 ( .ck(ispd_clk), .d(n_9374), .o(wishbone_slave_unit_del_sync_addr_out_reg_24__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_25__u0 ( .ck(ispd_clk), .d(n_8981), .o(wishbone_slave_unit_del_sync_addr_out_reg_25__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_26__u0 ( .ck(ispd_clk), .d(n_9371), .o(wishbone_slave_unit_del_sync_addr_out_reg_26__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_27__u0 ( .ck(ispd_clk), .d(n_9368), .o(wishbone_slave_unit_del_sync_addr_out_reg_27__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_28__u0 ( .ck(ispd_clk), .d(n_9366), .o(wishbone_slave_unit_del_sync_addr_out_reg_28__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_29__u0 ( .ck(ispd_clk), .d(n_9363), .o(wishbone_slave_unit_del_sync_addr_out_reg_29__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_2__u0 ( .ck(ispd_clk), .d(n_8979), .o(wishbone_slave_unit_del_sync_addr_out_reg_2__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_30__u0 ( .ck(ispd_clk), .d(n_9361), .o(wishbone_slave_unit_del_sync_addr_out_reg_30__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_31__u0 ( .ck(ispd_clk), .d(n_9358), .o(wishbone_slave_unit_del_sync_addr_out_reg_31__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_3__u0 ( .ck(ispd_clk), .d(n_9355), .o(wishbone_slave_unit_del_sync_addr_out_reg_3__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_4__u0 ( .ck(ispd_clk), .d(n_8977), .o(wishbone_slave_unit_del_sync_addr_out_reg_4__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_5__u0 ( .ck(ispd_clk), .d(n_8975), .o(wishbone_slave_unit_del_sync_addr_out_reg_5__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_6__u0 ( .ck(ispd_clk), .d(n_8973), .o(wishbone_slave_unit_del_sync_addr_out_reg_6__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_7__u0 ( .ck(ispd_clk), .d(n_9353), .o(wishbone_slave_unit_del_sync_addr_out_reg_7__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_8__u0 ( .ck(ispd_clk), .d(n_9350), .o(wishbone_slave_unit_del_sync_addr_out_reg_8__Q) );
ms00f80 wishbone_slave_unit_del_sync_addr_out_reg_9__u0 ( .ck(ispd_clk), .d(n_9348), .o(wishbone_slave_unit_del_sync_addr_out_reg_9__Q) );
ms00f80 wishbone_slave_unit_del_sync_bc_out_reg_0__u0 ( .ck(ispd_clk), .d(n_8598), .o(wishbone_slave_unit_del_sync_bc_out_reg_0__Q) );
in01f03 wishbone_slave_unit_del_sync_bc_out_reg_0__u1 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_0__Q), .o(wishbone_slave_unit_pcim_if_del_bc_in) );
ms00f80 wishbone_slave_unit_del_sync_bc_out_reg_1__u0 ( .ck(ispd_clk), .d(n_8677), .o(wishbone_slave_unit_del_sync_bc_out_reg_1__Q) );
ms00f80 wishbone_slave_unit_del_sync_bc_out_reg_2__u0 ( .ck(ispd_clk), .d(n_8723), .o(wishbone_slave_unit_del_sync_bc_out_reg_2__Q) );
in01m20 wishbone_slave_unit_del_sync_bc_out_reg_2__u1 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_2__Q), .o(wishbone_slave_unit_pcim_if_del_bc_in_382) );
ms00f80 wishbone_slave_unit_del_sync_bc_out_reg_3__u0 ( .ck(ispd_clk), .d(n_8796), .o(wishbone_slave_unit_del_sync_bc_out_reg_3__Q) );
in01s20 wishbone_slave_unit_del_sync_bc_out_reg_3__u1 ( .a(wishbone_slave_unit_del_sync_bc_out_reg_3__Q), .o(wishbone_slave_unit_pcim_if_del_bc_in_383) );
ms00f80 wishbone_slave_unit_del_sync_be_out_reg_0__u0 ( .ck(ispd_clk), .d(n_8676), .o(wishbone_slave_unit_fifos_wbr_be_in) );
ms00f80 wishbone_slave_unit_del_sync_be_out_reg_1__u0 ( .ck(ispd_clk), .d(n_8675), .o(wishbone_slave_unit_fifos_wbr_be_in_264) );
ms00f80 wishbone_slave_unit_del_sync_be_out_reg_2__u0 ( .ck(ispd_clk), .d(n_8674), .o(wishbone_slave_unit_fifos_wbr_be_in_265) );
ms00f80 wishbone_slave_unit_del_sync_be_out_reg_3__u0 ( .ck(ispd_clk), .d(n_8673), .o(wishbone_slave_unit_fifos_wbr_be_in_266) );
ms00f80 wishbone_slave_unit_del_sync_burst_out_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23546), .o(wishbone_slave_unit_pcim_if_del_burst_in) );
ms00f80 wishbone_slave_unit_del_sync_comp_comp_pending_reg_u0 ( .ck(ispd_clk), .d(n_8496), .o(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_0__u0 ( .ck(ispd_clk), .d(n_8652), .o(wishbone_slave_unit_del_sync_comp_cycle_count_0_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__u0 ( .ck(ispd_clk), .d(n_8656), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__Q) );
in01f40 wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_10__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_10_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__u0 ( .ck(ispd_clk), .d(n_8651), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__Q) );
in01f40 wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_11__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_11_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__u0 ( .ck(ispd_clk), .d(n_8662), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__Q) );
in01m20 wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_12__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_12_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__u0 ( .ck(ispd_clk), .d(n_8650), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_13__Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__u0 ( .ck(ispd_clk), .d(n_8649), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_14__Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__u0 ( .ck(ispd_clk), .d(n_8648), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_15__Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__u0 ( .ck(ispd_clk), .d(n_8579), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_1__u0 ( .ck(ispd_clk), .d(n_8658), .o(wishbone_slave_unit_del_sync_comp_cycle_count_1_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_2__u0 ( .ck(ispd_clk), .d(n_8647), .o(wishbone_slave_unit_del_sync_comp_cycle_count_2_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_3__u0 ( .ck(ispd_clk), .d(n_8646), .o(wishbone_slave_unit_del_sync_comp_cycle_count_3_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_4__u0 ( .ck(ispd_clk), .d(n_8645), .o(wishbone_slave_unit_del_sync_comp_cycle_count_4_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_5__u0 ( .ck(ispd_clk), .d(n_8644), .o(wishbone_slave_unit_del_sync_comp_cycle_count_5_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_6__u0 ( .ck(ispd_clk), .d(n_8643), .o(wishbone_slave_unit_del_sync_comp_cycle_count_6_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_7__u0 ( .ck(ispd_clk), .d(n_8642), .o(wishbone_slave_unit_del_sync_comp_cycle_count_7_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__u0 ( .ck(ispd_clk), .d(n_8661), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__Q) );
in01f40 wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_8__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_8_) );
ms00f80 wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__u0 ( .ck(ispd_clk), .d(n_8655), .o(wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__Q) );
in01f40 wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__u1 ( .a(wishbone_slave_unit_del_sync_comp_cycle_count_reg_9__Q), .o(wishbone_slave_unit_del_sync_comp_cycle_count_9_) );
ms00f80 wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_comp_done_reg_main), .o(TIMEBOOST_net_20757) );
in01s01 wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_u1 ( .a(wishbone_slave_unit_del_sync_comp_done_reg_clr_reg_Q), .o(wishbone_slave_unit_del_sync_comp_done_reg_clr) );
ms00f80 wishbone_slave_unit_del_sync_comp_done_reg_main_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_sync_comp_done), .o(wishbone_slave_unit_del_sync_comp_done_reg_main) );
ms00f80 wishbone_slave_unit_del_sync_comp_flush_out_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_comp_cycle_count_reg_16__Q), .o(wishbone_slave_unit_del_sync_comp_flush_out) );
ms00f80 wishbone_slave_unit_del_sync_comp_req_pending_reg_u0 ( .ck(ispd_clk), .d(n_7716), .o(wishbone_slave_unit_del_sync_comp_req_pending_reg_Q) );
in01f20 wishbone_slave_unit_del_sync_comp_req_pending_reg_u1 ( .a(wishbone_slave_unit_del_sync_comp_req_pending_reg_Q), .o(wishbone_slave_unit_pcim_if_del_req_in) );
ms00f80 wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_sync_comp_rty_exp_clr), .o(wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_Q) );
in01s01 wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_u1 ( .a(wishbone_slave_unit_del_sync_comp_rty_exp_clr_reg_Q), .o(wishbone_slave_unit_del_sync_comp_rty_exp_clr) );
ms00f80 wishbone_slave_unit_del_sync_comp_rty_exp_reg_reg_u0 ( .ck(ispd_clk), .d(n_4140), .o(wishbone_slave_unit_del_sync_comp_rty_exp_reg) );
ms00f80 wishbone_slave_unit_del_sync_comp_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_comp_comp_pending_reg_Q), .o(TIMEBOOST_net_21117) );
ms00f80 wishbone_slave_unit_del_sync_done_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_325), .o(wishbone_slave_unit_del_sync_sync_comp_done) );
ms00f80 wishbone_slave_unit_del_sync_req_comp_pending_reg_u0 ( .ck(ispd_clk), .d(n_14621), .o(wishbone_slave_unit_del_sync_req_comp_pending) );
ms00f80 wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_sync_req_comp_pending), .o(wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_Q) );
in01s01 wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_u1 ( .a(wishbone_slave_unit_del_sync_req_comp_pending_sample_reg_Q), .o(wishbone_slave_unit_del_sync_req_comp_pending_sample) );
ms00f80 wishbone_slave_unit_del_sync_req_done_reg_reg_u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23548), .o(wishbone_slave_unit_del_sync_req_done_reg_reg_Q) );
in01m08 wishbone_slave_unit_del_sync_req_done_reg_reg_u1 ( .a(wishbone_slave_unit_del_sync_req_done_reg_reg_Q), .o(wishbone_slave_unit_del_sync_req_done_reg) );
ms00f80 wishbone_slave_unit_del_sync_req_req_pending_reg_u0 ( .ck(ispd_clk), .d(n_8495), .o(wishbone_slave_unit_wbs_sm_del_req_pending_in) );
ms00f80 wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_req_rty_exp_reg), .o(wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_Q) );
in01s01 wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_u1 ( .a(wishbone_slave_unit_del_sync_req_rty_exp_clr_reg_Q), .o(wishbone_slave_unit_del_sync_req_rty_exp_clr) );
ms00f80 wishbone_slave_unit_del_sync_req_rty_exp_reg_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_sync_req_rty_exp), .o(wishbone_slave_unit_del_sync_req_rty_exp_reg) );
ms00f80 wishbone_slave_unit_del_sync_req_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_wbs_sm_del_req_pending_in), .o(wishbone_slave_unit_del_sync_sync_comp_req_pending) );
ms00f80 wishbone_slave_unit_del_sync_rty_exp_back_prop_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_2386), .o(wishbone_slave_unit_del_sync_sync_comp_rty_exp_clr) );
ms00f80 wishbone_slave_unit_del_sync_rty_exp_sync_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_del_sync_comp_rty_exp_reg), .o(wishbone_slave_unit_del_sync_sync_req_rty_exp) );
ms00f80 wishbone_slave_unit_del_sync_we_out_reg_u0 ( .ck(ispd_clk), .d(n_8672), .o(wishbone_slave_unit_del_sync_we_out_reg_Q) );
in01f40 wishbone_slave_unit_del_sync_we_out_reg_u1 ( .a(wishbone_slave_unit_del_sync_we_out_reg_Q), .o(wishbone_slave_unit_pcim_if_del_we_in) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_70), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_70) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_10__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_80), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_80) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_11__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_81), .o(TIMEBOOST_net_13959) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_12__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_82), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_82) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_13__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_83), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_83) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_14__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_84), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_84) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_15__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_85), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_85) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_16__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_86), .o(TIMEBOOST_net_13957) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_17__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_87), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_87) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_18__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_88), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_88) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_19__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_89), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_89) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_71), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_71) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_20__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_90), .o(TIMEBOOST_net_21155) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_21__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_91), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_91) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_22__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_92), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_92) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_23__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_93), .o(TIMEBOOST_net_23386) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_24__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_94), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_94) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_25__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_95), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_95) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_26__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_96), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_96) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_27__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_97), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_97) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_28__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_98), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_98) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_29__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_99), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_99) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_72), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_72) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_30__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_100), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_100) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_31__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_101), .o(TIMEBOOST_net_13961) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_73), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_73) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_4__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_74), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_74) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_5__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_75), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_75) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_6__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_76), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_76) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_7__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_77), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_77) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_8__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_78), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_78) );
ms00f80 wishbone_slave_unit_delayed_write_data_comp_wdata_out_reg_9__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_delayed_write_data_comp_wdata_out_79), .o(wishbone_slave_unit_delayed_write_data_comp_wdata_out_79) );
ms00f80 wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_22), .o(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount) );
ms00f80 wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_inGreyCount_reg_1__Q), .o(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_49) );
ms00f80 wishbone_slave_unit_fifos_i_synchronizer_reg_inGreyCount_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_inGreyCount_reg_2__Q), .o(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_50) );
ms00f80 wishbone_slave_unit_fifos_inGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(n_9145), .o(wishbone_slave_unit_fifos_inGreyCount_reg_0__Q) );
in01s01 wishbone_slave_unit_fifos_inGreyCount_reg_0__u1 ( .a(wishbone_slave_unit_fifos_inGreyCount_reg_0__Q), .o(wishbone_slave_unit_fifos_inGreyCount_0_) );
ms00f80 wishbone_slave_unit_fifos_inGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(n_8920), .o(wishbone_slave_unit_fifos_inGreyCount_reg_1__Q) );
ms00f80 wishbone_slave_unit_fifos_inGreyCount_reg_2__u0 ( .ck(ispd_clk), .d(n_8919), .o(wishbone_slave_unit_fifos_inGreyCount_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_outGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(n_8717), .o(wishbone_slave_unit_fifos_outGreyCount_0_) );
ms00f80 wishbone_slave_unit_fifos_outGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(n_8589), .o(wishbone_slave_unit_fifos_outGreyCount_1_) );
ms00f80 wishbone_slave_unit_fifos_outGreyCount_reg_2__u0 ( .ck(ispd_clk), .d(n_8585), .o(wishbone_slave_unit_fifos_outGreyCount_2_) );
ms00f80 wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount), .o(wishbone_slave_unit_fifos_pci_clk_inGreyCount_0_) );
ms00f80 wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_49), .o(wishbone_slave_unit_fifos_pci_clk_inGreyCount_1_) );
ms00f80 wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_pci_clk_sync_inGreyCount_50), .o(wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__Q) );
in01f80 wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__u1 ( .a(wishbone_slave_unit_fifos_pci_clk_inGreyCount_reg_2__Q), .o(wishbone_slave_unit_fifos_pci_clk_inGreyCount_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_276), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_45) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_46) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_i_synchronizer_reg_wgrey_addr_sync_data_out_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_47) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__u0 ( .ck(ispd_clk), .d(n_9942), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__u0 ( .ck(ispd_clk), .d(n_9238), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_1__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_1_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__u0 ( .ck(ispd_clk), .d(n_9239), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__u0 ( .ck(ispd_clk), .d(n_9241), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_reg_3__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_plus_one_3_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__u0 ( .ck(ispd_clk), .d(n_9947), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__u0 ( .ck(ispd_clk), .d(n_9932), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_1__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__u0 ( .ck(ispd_clk), .d(n_9931), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__Q) );
in01f40 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__u0 ( .ck(ispd_clk), .d(n_9154), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_raddr_reg_3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__Q) );
in01f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_45), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__Q) );
in01f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_1__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_46), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__Q) );
in01f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_sync_wgrey_addr_47), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__Q) );
in01f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_reg_3__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rclk_wgrey_addr_3_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_9237), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_9236), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_9235), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_9234), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_rgrey_addr_3_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg_0__u0 ( .ck(ispd_clk), .d(n_6112), .o(wishbone_slave_unit_fifos_wbr_whole_waddr) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg_1__u0 ( .ck(ispd_clk), .d(n_7393), .o(wishbone_slave_unit_fifos_wbr_whole_waddr_104) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg_2__u0 ( .ck(ispd_clk), .d(n_5770), .o(wishbone_slave_unit_fifos_wbr_whole_waddr_105) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_waddr_reg_3__u0 ( .ck(ispd_clk), .d(n_6138), .o(wishbone_slave_unit_fifos_wbr_whole_waddr_106) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_7137), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__Q) );
in01s06 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_6937), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_5768), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_5766), .o(wishbone_slave_unit_fifos_wbr_fifo_ctrl_wgrey_addr_reg_3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_0__u0 ( .ck(ispd_clk), .d(n_13131), .o(wbs_wbb3_2_wbb2_dat_o_i) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_10__u0 ( .ck(ispd_clk), .d(n_13401), .o(wbs_wbb3_2_wbb2_dat_o_i_109) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_11__u0 ( .ck(ispd_clk), .d(n_13400), .o(wbs_wbb3_2_wbb2_dat_o_i_110) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_12__u0 ( .ck(ispd_clk), .d(n_13130), .o(wbs_wbb3_2_wbb2_dat_o_i_111) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_13__u0 ( .ck(ispd_clk), .d(n_13129), .o(wbs_wbb3_2_wbb2_dat_o_i_112) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_14__u0 ( .ck(ispd_clk), .d(n_13128), .o(wbs_wbb3_2_wbb2_dat_o_i_113) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_15__u0 ( .ck(ispd_clk), .d(n_13318), .o(wbs_wbb3_2_wbb2_dat_o_i_114) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_16__u0 ( .ck(ispd_clk), .d(n_13399), .o(wbs_wbb3_2_wbb2_dat_o_i_115) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_17__u0 ( .ck(ispd_clk), .d(n_13144), .o(wbs_wbb3_2_wbb2_dat_o_i_116) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_18__u0 ( .ck(ispd_clk), .d(n_13409), .o(wbs_wbb3_2_wbb2_dat_o_i_117) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_19__u0 ( .ck(ispd_clk), .d(n_13408), .o(wbs_wbb3_2_wbb2_dat_o_i_118) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_1__u0 ( .ck(ispd_clk), .d(n_13407), .o(wbs_wbb3_2_wbb2_dat_o_i_100) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_20__u0 ( .ck(ispd_clk), .d(n_13143), .o(wbs_wbb3_2_wbb2_dat_o_i_119) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_21__u0 ( .ck(ispd_clk), .d(n_13406), .o(wbs_wbb3_2_wbb2_dat_o_i_120) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_22__u0 ( .ck(ispd_clk), .d(n_13405), .o(wbs_wbb3_2_wbb2_dat_o_i_121) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_23__u0 ( .ck(ispd_clk), .d(n_13142), .o(wbs_wbb3_2_wbb2_dat_o_i_122) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_24__u0 ( .ck(ispd_clk), .d(n_13323), .o(wbs_wbb3_2_wbb2_dat_o_i_123) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_25__u0 ( .ck(ispd_clk), .d(n_15942), .o(wbs_wbb3_2_wbb2_dat_o_i_124) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_26__u0 ( .ck(ispd_clk), .d(n_13141), .o(wbs_wbb3_2_wbb2_dat_o_i_125) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_27__u0 ( .ck(ispd_clk), .d(n_13321), .o(wbs_wbb3_2_wbb2_dat_o_i_126) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_28__u0 ( .ck(ispd_clk), .d(n_13140), .o(wbs_wbb3_2_wbb2_dat_o_i_127) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_29__u0 ( .ck(ispd_clk), .d(n_13139), .o(wbs_wbb3_2_wbb2_dat_o_i_128) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_2__u0 ( .ck(ispd_clk), .d(n_13320), .o(wbs_wbb3_2_wbb2_dat_o_i_101) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_30__u0 ( .ck(ispd_clk), .d(n_13404), .o(wbs_wbb3_2_wbb2_dat_o_i_129) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_31__u0 ( .ck(ispd_clk), .d(n_13138), .o(wbs_wbb3_2_wbb2_dat_o_i_130) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_36__u0 ( .ck(ispd_clk), .d(n_13319), .o(wishbone_slave_unit_wbs_sm_wbr_control_in) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_37__u0 ( .ck(ispd_clk), .d(n_13137), .o(wishbone_slave_unit_wbs_sm_wbr_control_in_190) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_3__u0 ( .ck(ispd_clk), .d(n_13136), .o(wbs_wbb3_2_wbb2_dat_o_i_102) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_4__u0 ( .ck(ispd_clk), .d(n_13135), .o(wbs_wbb3_2_wbb2_dat_o_i_103) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_5__u0 ( .ck(ispd_clk), .d(n_13403), .o(wbs_wbb3_2_wbb2_dat_o_i_104) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_6__u0 ( .ck(ispd_clk), .d(n_13402), .o(wbs_wbb3_2_wbb2_dat_o_i_105) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_7__u0 ( .ck(ispd_clk), .d(n_13134), .o(wbs_wbb3_2_wbb2_dat_o_i_106) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_8__u0 ( .ck(ispd_clk), .d(n_13133), .o(wbs_wbb3_2_wbb2_dat_o_i_107) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_do_reg_b_reg_9__u0 ( .ck(ispd_clk), .d(n_13132), .o(wbs_wbb3_2_wbb2_dat_o_i_108) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__u0 ( .ck(ispd_clk), .d(n_6926), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__u0 ( .ck(ispd_clk), .d(n_6924), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__u0 ( .ck(ispd_clk), .d(n_6922), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__u0 ( .ck(ispd_clk), .d(n_6920), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__12__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__51) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__u0 ( .ck(ispd_clk), .d(n_6919), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__u0 ( .ck(ispd_clk), .d(n_6917), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__u0 ( .ck(ispd_clk), .d(n_6915), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__u0 ( .ck(ispd_clk), .d(n_6913), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__u0 ( .ck(ispd_clk), .d(n_6911), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__17__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__56) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__u0 ( .ck(ispd_clk), .d(n_6910), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__u0 ( .ck(ispd_clk), .d(n_6908), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__u0 ( .ck(ispd_clk), .d(n_6905), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__u0 ( .ck(ispd_clk), .d(n_6903), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__20__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__59) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__u0 ( .ck(ispd_clk), .d(n_6902), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__u0 ( .ck(ispd_clk), .d(n_6900), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__u0 ( .ck(ispd_clk), .d(n_6898), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__23__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__62) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__u0 ( .ck(ispd_clk), .d(n_6897), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__u0 ( .ck(ispd_clk), .d(n_6895), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__u0 ( .ck(ispd_clk), .d(n_6892), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__u0 ( .ck(ispd_clk), .d(n_6889), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__u0 ( .ck(ispd_clk), .d(n_6887), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__28__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__67) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__u0 ( .ck(ispd_clk), .d(n_6885), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__u0 ( .ck(ispd_clk), .d(n_6883), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__u0 ( .ck(ispd_clk), .d(n_6878), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__u0 ( .ck(ispd_clk), .d(n_6876), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__31__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__70) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__u0 ( .ck(ispd_clk), .d(n_6097), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__u0 ( .ck(ispd_clk), .d(n_7392), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__u0 ( .ck(ispd_clk), .d(n_6875), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__u0 ( .ck(ispd_clk), .d(n_6872), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__4__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__43) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__u0 ( .ck(ispd_clk), .d(n_6140), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__u0 ( .ck(ispd_clk), .d(n_6871), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__u0 ( .ck(ispd_clk), .d(n_6869), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__Q) );
in01s02 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__7__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__46) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__u0 ( .ck(ispd_clk), .d(n_6868), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__8__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_0__47) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__u0 ( .ck(ispd_clk), .d(n_6867), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_0__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__u0 ( .ck(ispd_clk), .d(n_6865), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__u0 ( .ck(ispd_clk), .d(n_6932), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__u0 ( .ck(ispd_clk), .d(n_6863), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__u0 ( .ck(ispd_clk), .d(n_6861), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__u0 ( .ck(ispd_clk), .d(n_6859), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__u0 ( .ck(ispd_clk), .d(n_6857), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__u0 ( .ck(ispd_clk), .d(n_6855), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__u0 ( .ck(ispd_clk), .d(n_6853), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__u0 ( .ck(ispd_clk), .d(n_6851), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__u0 ( .ck(ispd_clk), .d(n_6934), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__u0 ( .ck(ispd_clk), .d(n_6849), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__u0 ( .ck(ispd_clk), .d(n_6847), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__u0 ( .ck(ispd_clk), .d(n_6845), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__u0 ( .ck(ispd_clk), .d(n_6709), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__u0 ( .ck(ispd_clk), .d(n_6842), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__u0 ( .ck(ispd_clk), .d(n_6840), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__u0 ( .ck(ispd_clk), .d(n_6837), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__u0 ( .ck(ispd_clk), .d(n_6835), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__u0 ( .ck(ispd_clk), .d(n_6833), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__u0 ( .ck(ispd_clk), .d(n_6747), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__u0 ( .ck(ispd_clk), .d(n_6830), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__u0 ( .ck(ispd_clk), .d(n_6828), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__u0 ( .ck(ispd_clk), .d(n_6826), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__u0 ( .ck(ispd_clk), .d(n_6824), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__u0 ( .ck(ispd_clk), .d(n_6821), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__u0 ( .ck(ispd_clk), .d(n_6129), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__u0 ( .ck(ispd_clk), .d(n_7390), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__u0 ( .ck(ispd_clk), .d(n_6819), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__u0 ( .ck(ispd_clk), .d(n_6816), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__u0 ( .ck(ispd_clk), .d(n_6880), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__u0 ( .ck(ispd_clk), .d(n_6814), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__u0 ( .ck(ispd_clk), .d(n_6812), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__u0 ( .ck(ispd_clk), .d(n_6809), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__u0 ( .ck(ispd_clk), .d(n_6150), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_10__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__u0 ( .ck(ispd_clk), .d(n_6095), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__u0 ( .ck(ispd_clk), .d(n_5812), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__u0 ( .ck(ispd_clk), .d(n_6093), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__u0 ( .ck(ispd_clk), .d(n_6091), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__u0 ( .ck(ispd_clk), .d(n_5816), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__u0 ( .ck(ispd_clk), .d(n_6089), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__u0 ( .ck(ispd_clk), .d(n_6099), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__u0 ( .ck(ispd_clk), .d(n_6087), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__u0 ( .ck(ispd_clk), .d(n_6085), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__u0 ( .ck(ispd_clk), .d(n_6103), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__u0 ( .ck(ispd_clk), .d(n_6083), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__u0 ( .ck(ispd_clk), .d(n_6107), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__u0 ( .ck(ispd_clk), .d(n_6081), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__u0 ( .ck(ispd_clk), .d(n_5840), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__u0 ( .ck(ispd_clk), .d(n_5848), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__u0 ( .ck(ispd_clk), .d(n_6079), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__u0 ( .ck(ispd_clk), .d(n_6077), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__u0 ( .ck(ispd_clk), .d(n_6111), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__u0 ( .ck(ispd_clk), .d(n_6075), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__u0 ( .ck(ispd_clk), .d(n_5810), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__u0 ( .ck(ispd_clk), .d(n_5806), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__u0 ( .ck(ispd_clk), .d(n_5822), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__u0 ( .ck(ispd_clk), .d(n_6073), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__u0 ( .ck(ispd_clk), .d(n_5792), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__u0 ( .ck(ispd_clk), .d(n_6071), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23550), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__u0 ( .ck(ispd_clk), .d(n_7388), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__Q) );
in01m06 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_11__466) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__u0 ( .ck(ispd_clk), .d(n_5981), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__u0 ( .ck(ispd_clk), .d(n_6069), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__u0 ( .ck(ispd_clk), .d(n_6109), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__u0 ( .ck(ispd_clk), .d(n_6067), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__u0 ( .ck(ispd_clk), .d(n_6065), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__u0 ( .ck(ispd_clk), .d(n_6063), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__u0 ( .ck(ispd_clk), .d(n_6101), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_11__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__u0 ( .ck(ispd_clk), .d(n_6806), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__u0 ( .ck(ispd_clk), .d(n_6804), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__u0 ( .ck(ispd_clk), .d(n_6801), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__u0 ( .ck(ispd_clk), .d(n_6799), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__u0 ( .ck(ispd_clk), .d(n_6797), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__u0 ( .ck(ispd_clk), .d(n_6795), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__u0 ( .ck(ispd_clk), .d(n_6156), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__u0 ( .ck(ispd_clk), .d(n_6793), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__16__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__484) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__u0 ( .ck(ispd_clk), .d(n_6158), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__u0 ( .ck(ispd_clk), .d(n_6791), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__u0 ( .ck(ispd_clk), .d(n_6789), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__19__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_12__487) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__u0 ( .ck(ispd_clk), .d(n_6788), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__u0 ( .ck(ispd_clk), .d(n_6785), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__u0 ( .ck(ispd_clk), .d(n_6783), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__u0 ( .ck(ispd_clk), .d(n_6781), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__u0 ( .ck(ispd_clk), .d(n_6778), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__u0 ( .ck(ispd_clk), .d(n_6776), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__u0 ( .ck(ispd_clk), .d(n_6774), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__u0 ( .ck(ispd_clk), .d(n_6929), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__u0 ( .ck(ispd_clk), .d(n_6772), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__u0 ( .ck(ispd_clk), .d(n_6770), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__u0 ( .ck(ispd_clk), .d(n_6768), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__u0 ( .ck(ispd_clk), .d(n_6766), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__u0 ( .ck(ispd_clk), .d(n_6763), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__u0 ( .ck(ispd_clk), .d(n_6761), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__u0 ( .ck(ispd_clk), .d(n_6127), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__u0 ( .ck(ispd_clk), .d(n_7366), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__u0 ( .ck(ispd_clk), .d(n_6759), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__u0 ( .ck(ispd_clk), .d(n_6757), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__u0 ( .ck(ispd_clk), .d(n_6754), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__u0 ( .ck(ispd_clk), .d(n_6514), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__u0 ( .ck(ispd_clk), .d(n_6752), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__u0 ( .ck(ispd_clk), .d(n_6745), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__u0 ( .ck(ispd_clk), .d(n_6749), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_12__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__u0 ( .ck(ispd_clk), .d(n_6061), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__0__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13_) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__u0 ( .ck(ispd_clk), .d(n_6060), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__u0 ( .ck(ispd_clk), .d(n_6058), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__u0 ( .ck(ispd_clk), .d(n_6056), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__u0 ( .ck(ispd_clk), .d(n_5772), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__u0 ( .ck(ispd_clk), .d(n_5774), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__u0 ( .ck(ispd_clk), .d(n_6054), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__15__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__522) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__u0 ( .ck(ispd_clk), .d(n_5804), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__u0 ( .ck(ispd_clk), .d(n_6053), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__u0 ( .ck(ispd_clk), .d(n_5838), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__u0 ( .ck(ispd_clk), .d(n_6051), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__u0 ( .ck(ispd_clk), .d(n_5844), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__u0 ( .ck(ispd_clk), .d(n_6049), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__u0 ( .ck(ispd_clk), .d(n_6047), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__u0 ( .ck(ispd_clk), .d(n_5854), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__u0 ( .ck(ispd_clk), .d(n_5858), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__u0 ( .ck(ispd_clk), .d(n_5967), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__24__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__531) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__u0 ( .ck(ispd_clk), .d(n_5850), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__25__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__532) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__u0 ( .ck(ispd_clk), .d(n_6045), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__u0 ( .ck(ispd_clk), .d(n_5794), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__u0 ( .ck(ispd_clk), .d(n_6043), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__u0 ( .ck(ispd_clk), .d(n_6041), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__29__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__536) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__u0 ( .ck(ispd_clk), .d(n_6040), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__509) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__u0 ( .ck(ispd_clk), .d(n_5936), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__u0 ( .ck(ispd_clk), .d(n_6039), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__u0 ( .ck(ispd_clk), .d(n_5800), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__u0 ( .ck(ispd_clk), .d(n_7387), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_13__544) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__u0 ( .ck(ispd_clk), .d(n_5870), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__u0 ( .ck(ispd_clk), .d(n_6037), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__u0 ( .ck(ispd_clk), .d(n_5776), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__u0 ( .ck(ispd_clk), .d(n_6035), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__u0 ( .ck(ispd_clk), .d(n_5814), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__u0 ( .ck(ispd_clk), .d(n_6033), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__u0 ( .ck(ispd_clk), .d(n_5833), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_13__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__u0 ( .ck(ispd_clk), .d(n_6031), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__u0 ( .ck(ispd_clk), .d(n_6029), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__u0 ( .ck(ispd_clk), .d(n_5862), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__u0 ( .ck(ispd_clk), .d(n_6027), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__u0 ( .ck(ispd_clk), .d(n_6025), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__u0 ( .ck(ispd_clk), .d(n_6023), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__u0 ( .ck(ispd_clk), .d(n_5796), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__u0 ( .ck(ispd_clk), .d(n_6021), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__u0 ( .ck(ispd_clk), .d(n_6019), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__u0 ( .ck(ispd_clk), .d(n_6017), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__u0 ( .ck(ispd_clk), .d(n_6015), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__u0 ( .ck(ispd_clk), .d(n_6013), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__u0 ( .ck(ispd_clk), .d(n_6105), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__u0 ( .ck(ispd_clk), .d(n_6011), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__u0 ( .ck(ispd_clk), .d(n_6009), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__u0 ( .ck(ispd_clk), .d(n_6007), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__u0 ( .ck(ispd_clk), .d(n_5830), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__u0 ( .ck(ispd_clk), .d(n_6005), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__u0 ( .ck(ispd_clk), .d(n_6003), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__u0 ( .ck(ispd_clk), .d(n_6001), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__u0 ( .ck(ispd_clk), .d(n_5798), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__u0 ( .ck(ispd_clk), .d(n_5999), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__u0 ( .ck(ispd_clk), .d(n_5997), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__u0 ( .ck(ispd_clk), .d(n_5995), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__u0 ( .ck(ispd_clk), .d(n_5993), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__u0 ( .ck(ispd_clk), .d(n_5991), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__u0 ( .ck(ispd_clk), .d(n_7364), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_14__583) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__u0 ( .ck(ispd_clk), .d(n_5989), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__u0 ( .ck(ispd_clk), .d(n_5987), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__u0 ( .ck(ispd_clk), .d(n_5985), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__u0 ( .ck(ispd_clk), .d(n_5827), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__u0 ( .ck(ispd_clk), .d(n_5983), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__u0 ( .ck(ispd_clk), .d(n_5868), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__u0 ( .ck(ispd_clk), .d(n_5979), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_14__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__u0 ( .ck(ispd_clk), .d(n_5856), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__u0 ( .ck(ispd_clk), .d(n_5842), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__u0 ( .ck(ispd_clk), .d(n_5977), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__u0 ( .ck(ispd_clk), .d(n_5975), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__u0 ( .ck(ispd_clk), .d(n_5973), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__u0 ( .ck(ispd_clk), .d(n_5864), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__u0 ( .ck(ispd_clk), .d(n_5971), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__u0 ( .ck(ispd_clk), .d(n_5824), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__u0 ( .ck(ispd_clk), .d(n_5969), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__u0 ( .ck(ispd_clk), .d(n_5866), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__u0 ( .ck(ispd_clk), .d(n_5966), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__u0 ( .ck(ispd_clk), .d(n_5964), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__u0 ( .ck(ispd_clk), .d(n_5962), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__u0 ( .ck(ispd_clk), .d(n_5782), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__u0 ( .ck(ispd_clk), .d(n_5960), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__u0 ( .ck(ispd_clk), .d(n_5784), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__u0 ( .ck(ispd_clk), .d(n_5958), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__u0 ( .ck(ispd_clk), .d(n_5786), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__u0 ( .ck(ispd_clk), .d(n_5956), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__u0 ( .ck(ispd_clk), .d(n_5954), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__u0 ( .ck(ispd_clk), .d(n_5952), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__u0 ( .ck(ispd_clk), .d(n_5788), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__u0 ( .ck(ispd_clk), .d(n_5950), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__u0 ( .ck(ispd_clk), .d(n_5802), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__u0 ( .ck(ispd_clk), .d(n_5948), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__u0 ( .ck(ispd_clk), .d(n_5808), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__u0 ( .ck(ispd_clk), .d(n_7386), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_15__622) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__u0 ( .ck(ispd_clk), .d(n_5819), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__u0 ( .ck(ispd_clk), .d(n_5946), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__u0 ( .ck(ispd_clk), .d(n_5860), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__u0 ( .ck(ispd_clk), .d(n_5780), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__u0 ( .ck(ispd_clk), .d(n_5778), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__u0 ( .ck(ispd_clk), .d(n_5944), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__u0 ( .ck(ispd_clk), .d(n_5942), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_15__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__u0 ( .ck(ispd_clk), .d(n_6743), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__u0 ( .ck(ispd_clk), .d(n_6741), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__u0 ( .ck(ispd_clk), .d(n_6738), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__u0 ( .ck(ispd_clk), .d(n_6735), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__u0 ( .ck(ispd_clk), .d(n_6733), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__u0 ( .ck(ispd_clk), .d(n_6731), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__u0 ( .ck(ispd_clk), .d(n_6729), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__u0 ( .ck(ispd_clk), .d(n_6726), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__u0 ( .ck(ispd_clk), .d(n_6724), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__u0 ( .ck(ispd_clk), .d(n_6162), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__u0 ( .ck(ispd_clk), .d(n_6722), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__u0 ( .ck(ispd_clk), .d(n_6720), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__u0 ( .ck(ispd_clk), .d(n_6718), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__u0 ( .ck(ispd_clk), .d(n_6716), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__u0 ( .ck(ispd_clk), .d(n_6142), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__u0 ( .ck(ispd_clk), .d(n_6714), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__u0 ( .ck(ispd_clk), .d(n_6152), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__u0 ( .ck(ispd_clk), .d(n_6712), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__u0 ( .ck(ispd_clk), .d(n_6154), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__u0 ( .ck(ispd_clk), .d(n_6707), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__u0 ( .ck(ispd_clk), .d(n_6705), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__u0 ( .ck(ispd_clk), .d(n_6144), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__u0 ( .ck(ispd_clk), .d(n_6146), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__u0 ( .ck(ispd_clk), .d(n_6703), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__u0 ( .ck(ispd_clk), .d(n_6148), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__u0 ( .ck(ispd_clk), .d(n_5836), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__u0 ( .ck(ispd_clk), .d(n_7385), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__u0 ( .ck(ispd_clk), .d(n_6701), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__u0 ( .ck(ispd_clk), .d(n_6699), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__u0 ( .ck(ispd_clk), .d(n_6171), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__u0 ( .ck(ispd_clk), .d(n_6697), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__u0 ( .ck(ispd_clk), .d(n_6695), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__u0 ( .ck(ispd_clk), .d(n_6693), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__u0 ( .ck(ispd_clk), .d(n_6691), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_1__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__u0 ( .ck(ispd_clk), .d(n_6689), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__u0 ( .ck(ispd_clk), .d(n_6686), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__u0 ( .ck(ispd_clk), .d(n_6684), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__u0 ( .ck(ispd_clk), .d(n_6682), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__u0 ( .ck(ispd_clk), .d(n_6680), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__u0 ( .ck(ispd_clk), .d(n_6678), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__u0 ( .ck(ispd_clk), .d(n_6676), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__u0 ( .ck(ispd_clk), .d(n_6674), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__u0 ( .ck(ispd_clk), .d(n_6672), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__u0 ( .ck(ispd_clk), .d(n_6670), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__u0 ( .ck(ispd_clk), .d(n_6668), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__u0 ( .ck(ispd_clk), .d(n_6665), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__u0 ( .ck(ispd_clk), .d(n_6662), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__u0 ( .ck(ispd_clk), .d(n_6659), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__u0 ( .ck(ispd_clk), .d(n_6657), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__u0 ( .ck(ispd_clk), .d(n_6654), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__u0 ( .ck(ispd_clk), .d(n_6651), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__u0 ( .ck(ispd_clk), .d(n_6649), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__u0 ( .ck(ispd_clk), .d(n_6647), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__u0 ( .ck(ispd_clk), .d(n_6644), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__u0 ( .ck(ispd_clk), .d(n_6641), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__u0 ( .ck(ispd_clk), .d(n_6639), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__u0 ( .ck(ispd_clk), .d(n_6636), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__u0 ( .ck(ispd_clk), .d(n_6634), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__u0 ( .ck(ispd_clk), .d(n_6631), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__u0 ( .ck(ispd_clk), .d(n_5940), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__u0 ( .ck(ispd_clk), .d(n_7383), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__u0 ( .ck(ispd_clk), .d(n_6629), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__u0 ( .ck(ispd_clk), .d(n_6626), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__u0 ( .ck(ispd_clk), .d(n_6623), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__u0 ( .ck(ispd_clk), .d(n_6621), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__6__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_2__6) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__u0 ( .ck(ispd_clk), .d(n_6620), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__u0 ( .ck(ispd_clk), .d(n_6617), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__u0 ( .ck(ispd_clk), .d(n_6615), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_2__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__u0 ( .ck(ispd_clk), .d(n_6613), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__u0 ( .ck(ispd_clk), .d(n_6610), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__u0 ( .ck(ispd_clk), .d(n_6607), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__u0 ( .ck(ispd_clk), .d(n_6605), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__u0 ( .ck(ispd_clk), .d(n_6603), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__u0 ( .ck(ispd_clk), .d(n_6601), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__u0 ( .ck(ispd_clk), .d(n_6598), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__u0 ( .ck(ispd_clk), .d(n_6596), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__u0 ( .ck(ispd_clk), .d(n_6594), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__u0 ( .ck(ispd_clk), .d(n_6592), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__u0 ( .ck(ispd_clk), .d(n_6589), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__u0 ( .ck(ispd_clk), .d(n_6587), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__u0 ( .ck(ispd_clk), .d(n_6585), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__u0 ( .ck(ispd_clk), .d(n_6582), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__21__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__177) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__u0 ( .ck(ispd_clk), .d(n_6580), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__22__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__178) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__u0 ( .ck(ispd_clk), .d(n_6578), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__u0 ( .ck(ispd_clk), .d(n_6575), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__u0 ( .ck(ispd_clk), .d(n_6572), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__u0 ( .ck(ispd_clk), .d(n_6569), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__u0 ( .ck(ispd_clk), .d(n_6567), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__Q) );
in01m01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__27__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_3__183) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__u0 ( .ck(ispd_clk), .d(n_6566), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__u0 ( .ck(ispd_clk), .d(n_6563), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__u0 ( .ck(ispd_clk), .d(n_6561), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__u0 ( .ck(ispd_clk), .d(n_6558), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__u0 ( .ck(ispd_clk), .d(n_6556), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__u0 ( .ck(ispd_clk), .d(n_6123), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__u0 ( .ck(ispd_clk), .d(n_7381), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__u0 ( .ck(ispd_clk), .d(n_6553), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__u0 ( .ck(ispd_clk), .d(n_6550), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__u0 ( .ck(ispd_clk), .d(n_6548), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__u0 ( .ck(ispd_clk), .d(n_6546), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__u0 ( .ck(ispd_clk), .d(n_6543), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__u0 ( .ck(ispd_clk), .d(n_6541), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__u0 ( .ck(ispd_clk), .d(n_6538), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_3__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__u0 ( .ck(ispd_clk), .d(n_6536), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__u0 ( .ck(ispd_clk), .d(n_6534), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__u0 ( .ck(ispd_clk), .d(n_6532), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__u0 ( .ck(ispd_clk), .d(n_6530), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__u0 ( .ck(ispd_clk), .d(n_6528), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__u0 ( .ck(ispd_clk), .d(n_6526), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__u0 ( .ck(ispd_clk), .d(n_6523), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__u0 ( .ck(ispd_clk), .d(n_6521), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__u0 ( .ck(ispd_clk), .d(n_6518), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__u0 ( .ck(ispd_clk), .d(n_6516), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__u0 ( .ck(ispd_clk), .d(n_6166), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__u0 ( .ck(ispd_clk), .d(n_6512), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__u0 ( .ck(ispd_clk), .d(n_6509), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__u0 ( .ck(ispd_clk), .d(n_6168), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__u0 ( .ck(ispd_clk), .d(n_6506), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__u0 ( .ck(ispd_clk), .d(n_6504), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__u0 ( .ck(ispd_clk), .d(n_6501), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__u0 ( .ck(ispd_clk), .d(n_6498), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__u0 ( .ck(ispd_clk), .d(n_6495), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__u0 ( .ck(ispd_clk), .d(n_6493), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__u0 ( .ck(ispd_clk), .d(n_6490), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__u0 ( .ck(ispd_clk), .d(n_6488), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__u0 ( .ck(ispd_clk), .d(n_6485), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__u0 ( .ck(ispd_clk), .d(n_6483), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__u0 ( .ck(ispd_clk), .d(n_6480), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__u0 ( .ck(ispd_clk), .d(n_5938), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__u0 ( .ck(ispd_clk), .d(n_7379), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__u0 ( .ck(ispd_clk), .d(n_6477), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__u0 ( .ck(ispd_clk), .d(n_6475), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__u0 ( .ck(ispd_clk), .d(n_6473), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__u0 ( .ck(ispd_clk), .d(n_6470), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__u0 ( .ck(ispd_clk), .d(n_6468), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__u0 ( .ck(ispd_clk), .d(n_6465), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__u0 ( .ck(ispd_clk), .d(n_6463), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_4__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__u0 ( .ck(ispd_clk), .d(n_6461), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__u0 ( .ck(ispd_clk), .d(n_6458), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__u0 ( .ck(ispd_clk), .d(n_6160), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__u0 ( .ck(ispd_clk), .d(n_6456), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__u0 ( .ck(ispd_clk), .d(n_6453), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__u0 ( .ck(ispd_clk), .d(n_6451), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__u0 ( .ck(ispd_clk), .d(n_6448), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__u0 ( .ck(ispd_clk), .d(n_6446), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__u0 ( .ck(ispd_clk), .d(n_6443), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__u0 ( .ck(ispd_clk), .d(n_6440), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__u0 ( .ck(ispd_clk), .d(n_6438), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__u0 ( .ck(ispd_clk), .d(n_6435), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__u0 ( .ck(ispd_clk), .d(n_6433), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__u0 ( .ck(ispd_clk), .d(n_6430), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__u0 ( .ck(ispd_clk), .d(n_6427), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__u0 ( .ck(ispd_clk), .d(n_6425), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__u0 ( .ck(ispd_clk), .d(n_6423), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__u0 ( .ck(ispd_clk), .d(n_6420), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__u0 ( .ck(ispd_clk), .d(n_6417), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__u0 ( .ck(ispd_clk), .d(n_6415), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__u0 ( .ck(ispd_clk), .d(n_6413), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__u0 ( .ck(ispd_clk), .d(n_6410), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__u0 ( .ck(ispd_clk), .d(n_6407), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__u0 ( .ck(ispd_clk), .d(n_6405), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__u0 ( .ck(ispd_clk), .d(n_6402), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__u0 ( .ck(ispd_clk), .d(n_6121), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__u0 ( .ck(ispd_clk), .d(n_7377), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__u0 ( .ck(ispd_clk), .d(n_6400), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__u0 ( .ck(ispd_clk), .d(n_6398), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__u0 ( .ck(ispd_clk), .d(n_6395), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__u0 ( .ck(ispd_clk), .d(n_6393), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__u0 ( .ck(ispd_clk), .d(n_6390), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__u0 ( .ck(ispd_clk), .d(n_6388), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__u0 ( .ck(ispd_clk), .d(n_6386), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_5__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__u0 ( .ck(ispd_clk), .d(n_6384), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__u0 ( .ck(ispd_clk), .d(n_6382), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__u0 ( .ck(ispd_clk), .d(n_6379), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__u0 ( .ck(ispd_clk), .d(n_6376), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__u0 ( .ck(ispd_clk), .d(n_6374), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__13__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__247) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__u0 ( .ck(ispd_clk), .d(n_6373), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__Q) );
in01s20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__14__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__248) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__u0 ( .ck(ispd_clk), .d(n_6372), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__15__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__249) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__u0 ( .ck(ispd_clk), .d(n_6371), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__u0 ( .ck(ispd_clk), .d(n_6369), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__u0 ( .ck(ispd_clk), .d(n_6366), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__u0 ( .ck(ispd_clk), .d(n_6364), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__u0 ( .ck(ispd_clk), .d(n_6361), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__u0 ( .ck(ispd_clk), .d(n_6358), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__u0 ( .ck(ispd_clk), .d(n_6355), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__u0 ( .ck(ispd_clk), .d(n_6353), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__u0 ( .ck(ispd_clk), .d(n_6350), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__u0 ( .ck(ispd_clk), .d(n_6348), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__24__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__258) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__u0 ( .ck(ispd_clk), .d(n_6347), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__u0 ( .ck(ispd_clk), .d(n_6345), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__26__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__260) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__u0 ( .ck(ispd_clk), .d(n_6344), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__u0 ( .ck(ispd_clk), .d(n_6342), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__u0 ( .ck(ispd_clk), .d(n_6340), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__u0 ( .ck(ispd_clk), .d(n_6338), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__2__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__236) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__u0 ( .ck(ispd_clk), .d(n_6337), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__u0 ( .ck(ispd_clk), .d(n_6335), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__31__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__265) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__u0 ( .ck(ispd_clk), .d(n_6119), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__u0 ( .ck(ispd_clk), .d(n_7375), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__Q) );
in01m03 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__271) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__u0 ( .ck(ispd_clk), .d(n_6334), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__Q) );
in01s01 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__3__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__237) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__u0 ( .ck(ispd_clk), .d(n_6333), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__4__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__238) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__u0 ( .ck(ispd_clk), .d(n_6331), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__u0 ( .ck(ispd_clk), .d(n_6329), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__u0 ( .ck(ispd_clk), .d(n_6327), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__u0 ( .ck(ispd_clk), .d(n_6325), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__u0 ( .ck(ispd_clk), .d(n_6323), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_6__9__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_6__243) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__u0 ( .ck(ispd_clk), .d(n_5846), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__u0 ( .ck(ispd_clk), .d(n_5934), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__u0 ( .ck(ispd_clk), .d(n_5932), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__u0 ( .ck(ispd_clk), .d(n_5930), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__u0 ( .ck(ispd_clk), .d(n_5928), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__u0 ( .ck(ispd_clk), .d(n_5926), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__u0 ( .ck(ispd_clk), .d(n_5924), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__u0 ( .ck(ispd_clk), .d(n_5922), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__u0 ( .ck(ispd_clk), .d(n_5920), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__u0 ( .ck(ispd_clk), .d(n_5918), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__u0 ( .ck(ispd_clk), .d(n_5916), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__u0 ( .ck(ispd_clk), .d(n_5914), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__u0 ( .ck(ispd_clk), .d(n_5912), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__u0 ( .ck(ispd_clk), .d(n_5910), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__u0 ( .ck(ispd_clk), .d(n_5908), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__u0 ( .ck(ispd_clk), .d(n_5906), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__u0 ( .ck(ispd_clk), .d(n_5852), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__u0 ( .ck(ispd_clk), .d(n_5904), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__u0 ( .ck(ispd_clk), .d(n_5902), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__u0 ( .ck(ispd_clk), .d(n_5900), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__u0 ( .ck(ispd_clk), .d(n_5898), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__u0 ( .ck(ispd_clk), .d(n_5896), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__u0 ( .ck(ispd_clk), .d(n_5894), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__u0 ( .ck(ispd_clk), .d(n_5892), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__u0 ( .ck(ispd_clk), .d(n_5890), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__u0 ( .ck(ispd_clk), .d(n_5888), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__u0 ( .ck(ispd_clk), .d(n_7374), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__Q) );
in01s03 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__37__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_7__310) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__u0 ( .ck(ispd_clk), .d(n_5886), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__u0 ( .ck(ispd_clk), .d(n_5884), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__u0 ( .ck(ispd_clk), .d(n_5882), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__u0 ( .ck(ispd_clk), .d(n_5880), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__u0 ( .ck(ispd_clk), .d(n_5878), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__u0 ( .ck(ispd_clk), .d(n_5876), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__u0 ( .ck(ispd_clk), .d(n_5874), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_7__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__u0 ( .ck(ispd_clk), .d(n_6321), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__u0 ( .ck(ispd_clk), .d(n_6318), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__u0 ( .ck(ispd_clk), .d(n_6315), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__u0 ( .ck(ispd_clk), .d(n_6313), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__u0 ( .ck(ispd_clk), .d(n_6311), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__u0 ( .ck(ispd_clk), .d(n_6308), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__u0 ( .ck(ispd_clk), .d(n_6305), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__u0 ( .ck(ispd_clk), .d(n_6303), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__u0 ( .ck(ispd_clk), .d(n_6301), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__u0 ( .ck(ispd_clk), .d(n_6298), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__18__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__330) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__u0 ( .ck(ispd_clk), .d(n_6297), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__u0 ( .ck(ispd_clk), .d(n_6295), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__u0 ( .ck(ispd_clk), .d(n_6292), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__u0 ( .ck(ispd_clk), .d(n_6289), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__u0 ( .ck(ispd_clk), .d(n_6286), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__u0 ( .ck(ispd_clk), .d(n_6284), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__u0 ( .ck(ispd_clk), .d(n_6281), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__u0 ( .ck(ispd_clk), .d(n_6278), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__u0 ( .ck(ispd_clk), .d(n_6164), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__u0 ( .ck(ispd_clk), .d(n_6276), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__u0 ( .ck(ispd_clk), .d(n_6273), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__u0 ( .ck(ispd_clk), .d(n_6271), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__u0 ( .ck(ispd_clk), .d(n_6268), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__u0 ( .ck(ispd_clk), .d(n_6266), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__30__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_8__342) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__u0 ( .ck(ispd_clk), .d(n_6264), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__u0 ( .ck(ispd_clk), .d(n_5872), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__u0 ( .ck(ispd_clk), .d(n_7371), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__u0 ( .ck(ispd_clk), .d(n_6261), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__u0 ( .ck(ispd_clk), .d(n_6259), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__u0 ( .ck(ispd_clk), .d(n_6257), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__u0 ( .ck(ispd_clk), .d(n_6254), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__u0 ( .ck(ispd_clk), .d(n_6252), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__u0 ( .ck(ispd_clk), .d(n_6249), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__u0 ( .ck(ispd_clk), .d(n_6246), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_8__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__u0 ( .ck(ispd_clk), .d(n_6243), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__u0 ( .ck(ispd_clk), .d(n_6240), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__u0 ( .ck(ispd_clk), .d(n_6238), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__u0 ( .ck(ispd_clk), .d(n_6235), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__12__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__363) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__u0 ( .ck(ispd_clk), .d(n_6234), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__u0 ( .ck(ispd_clk), .d(n_6231), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__14__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__365) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__u0 ( .ck(ispd_clk), .d(n_6230), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__u0 ( .ck(ispd_clk), .d(n_6228), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__u0 ( .ck(ispd_clk), .d(n_6226), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__u0 ( .ck(ispd_clk), .d(n_6223), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__u0 ( .ck(ispd_clk), .d(n_6221), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__u0 ( .ck(ispd_clk), .d(n_6216), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__u0 ( .ck(ispd_clk), .d(n_6213), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__u0 ( .ck(ispd_clk), .d(n_6211), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__u0 ( .ck(ispd_clk), .d(n_6208), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__u0 ( .ck(ispd_clk), .d(n_6206), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__23__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__374) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__u0 ( .ck(ispd_clk), .d(n_6204), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__u0 ( .ck(ispd_clk), .d(n_6201), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__25__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__376) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__u0 ( .ck(ispd_clk), .d(n_6200), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__26__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__377) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__u0 ( .ck(ispd_clk), .d(n_6199), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__u0 ( .ck(ispd_clk), .d(n_6196), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__28__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__379) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__u0 ( .ck(ispd_clk), .d(n_6195), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__29__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__380) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__u0 ( .ck(ispd_clk), .d(n_6193), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__u0 ( .ck(ispd_clk), .d(n_6191), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__u0 ( .ck(ispd_clk), .d(n_6189), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__u0 ( .ck(ispd_clk), .d(n_6117), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__u0 ( .ck(ispd_clk), .d(n_7368), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__37__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__u0 ( .ck(ispd_clk), .d(n_6186), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__u0 ( .ck(ispd_clk), .d(n_6184), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__u0 ( .ck(ispd_clk), .d(n_6181), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__u0 ( .ck(ispd_clk), .d(n_6179), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__u0 ( .ck(ispd_clk), .d(n_6177), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__7__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__358) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__u0 ( .ck(ispd_clk), .d(n_6175), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__Q) );
in01m40 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__8__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__359) );
ms00f80 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__u0 ( .ck(ispd_clk), .d(n_6173), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__Q) );
in01m20 wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__u1 ( .a(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_reg_9__9__Q), .o(wishbone_slave_unit_fifos_wbr_fifo_storage_mem_9__360) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus1) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_93) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_94) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_rgrey_minus1_sync_data_out_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_95) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg_0__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23552), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg_1__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23554), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_70) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg_2__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23556), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_71) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_i_synchronizer_reg_wgrey_next_sync_data_out_reg_3__u0 ( .ck(ispd_clk), .d(TIMEBOOST_net_23558), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_72) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg_0__u0 ( .ck(ispd_clk), .d(n_8765), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg_1__u0 ( .ck(ispd_clk), .d(n_8713), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg_2__u0 ( .ck(ispd_clk), .d(n_8716), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_reg_3__u0 ( .ck(ispd_clk), .d(n_8714), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_plus_one_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg_0__u0 ( .ck(ispd_clk), .d(n_8745), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg_1__u0 ( .ck(ispd_clk), .d(n_8784), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg_2__u0 ( .ck(ispd_clk), .d(n_8712), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_reg_3__u0 ( .ck(ispd_clk), .d(n_8711), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_raddr_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_70), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_71), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_sync_wgrey_next_72), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rclk_wgrey_next_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_8709), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_8708), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_8707), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_8705), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_addr_reg_3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__u0 ( .ck(ispd_clk), .d(n_8703), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__u0 ( .ck(ispd_clk), .d(n_8701), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__u0 ( .ck(ispd_clk), .d(n_8699), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__u0 ( .ck(ispd_clk), .d(n_8697), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_minus1_reg_3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_8695), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_8694), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_8693), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_reg_3__u0 ( .ck(ispd_clk), .d(n_8692), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_rgrey_next_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg_0__u0 ( .ck(ispd_clk), .d(n_9340), .o(wishbone_slave_unit_fifos_wbw_whole_waddr) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg_1__u0 ( .ck(ispd_clk), .d(n_9343), .o(wishbone_slave_unit_fifos_wbw_whole_waddr_55) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg_2__u0 ( .ck(ispd_clk), .d(n_9194), .o(wishbone_slave_unit_fifos_wbw_whole_waddr_56) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_waddr_reg_3__u0 ( .ck(ispd_clk), .d(n_9189), .o(wishbone_slave_unit_fifos_wbw_whole_waddr_57) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg_0__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus1), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg_1__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_93), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg_2__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_94), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_reg_3__u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_sync_rgrey_minus_95), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wclk_rgrey_minus1_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg_0__u0 ( .ck(ispd_clk), .d(n_9187), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg_1__u0 ( .ck(ispd_clk), .d(n_9185), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg_2__u0 ( .ck(ispd_clk), .d(n_9184), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_reg_3__u0 ( .ck(ispd_clk), .d(n_9183), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_addr_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg_0__u0 ( .ck(ispd_clk), .d(n_9342), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg_1__u0 ( .ck(ispd_clk), .d(n_9192), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg_2__u0 ( .ck(ispd_clk), .d(n_9182), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_2_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_reg_3__u0 ( .ck(ispd_clk), .d(n_9181), .o(wishbone_slave_unit_fifos_wbw_fifo_ctrl_wgrey_next_3_) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_0__u0 ( .ck(ispd_clk), .d(n_12853), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_10__u0 ( .ck(ispd_clk), .d(n_12852), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_393) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_11__u0 ( .ck(ispd_clk), .d(n_12851), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_394) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_12__u0 ( .ck(ispd_clk), .d(n_12850), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_395) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_13__u0 ( .ck(ispd_clk), .d(n_12849), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_396) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_14__u0 ( .ck(ispd_clk), .d(n_12848), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_397) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_15__u0 ( .ck(ispd_clk), .d(n_12847), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_398) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_16__u0 ( .ck(ispd_clk), .d(n_12846), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_399) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_17__u0 ( .ck(ispd_clk), .d(n_12845), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_400) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_18__u0 ( .ck(ispd_clk), .d(n_15565), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_401) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_19__u0 ( .ck(ispd_clk), .d(n_12843), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_402) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_1__u0 ( .ck(ispd_clk), .d(n_12842), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_384) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_20__u0 ( .ck(ispd_clk), .d(n_12841), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_403) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_21__u0 ( .ck(ispd_clk), .d(n_12775), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_404) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_22__u0 ( .ck(ispd_clk), .d(n_12840), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_405) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_23__u0 ( .ck(ispd_clk), .d(n_12839), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_406) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_24__u0 ( .ck(ispd_clk), .d(n_15540), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_407) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_25__u0 ( .ck(ispd_clk), .d(n_12774), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_408) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_26__u0 ( .ck(ispd_clk), .d(n_12951), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_409) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_27__u0 ( .ck(ispd_clk), .d(n_12837), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_410) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_28__u0 ( .ck(ispd_clk), .d(n_12836), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_411) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_29__u0 ( .ck(ispd_clk), .d(n_12835), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_412) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_2__u0 ( .ck(ispd_clk), .d(n_12834), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_385) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_30__u0 ( .ck(ispd_clk), .d(n_12773), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_413) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_31__u0 ( .ck(ispd_clk), .d(n_12833), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_414) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_32__u0 ( .ck(ispd_clk), .d(n_12832), .o(wishbone_slave_unit_pcim_if_wbw_cbe_in) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__u0 ( .ck(ispd_clk), .d(n_12831), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_34__u0 ( .ck(ispd_clk), .d(n_12830), .o(wishbone_slave_unit_pcim_if_wbw_cbe_in_416) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_35__u0 ( .ck(ispd_clk), .d(n_12829), .o(wishbone_slave_unit_pcim_if_wbw_cbe_in_417) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__u0 ( .ck(ispd_clk), .d(n_12828), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_3__u0 ( .ck(ispd_clk), .d(n_12827), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_386) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_4__u0 ( .ck(ispd_clk), .d(n_12826), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_387) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_5__u0 ( .ck(ispd_clk), .d(n_12825), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_388) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_6__u0 ( .ck(ispd_clk), .d(n_12824), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_389) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_7__u0 ( .ck(ispd_clk), .d(n_12823), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_390) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_8__u0 ( .ck(ispd_clk), .d(n_12822), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_391) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_do_reg_b_reg_9__u0 ( .ck(ispd_clk), .d(n_12821), .o(wishbone_slave_unit_pcim_if_wbw_addr_data_in_392) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__u0 ( .ck(ispd_clk), .d(n_11513), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__u0 ( .ck(ispd_clk), .d(n_11512), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__u0 ( .ck(ispd_clk), .d(n_11510), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__u0 ( .ck(ispd_clk), .d(n_10424), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__u0 ( .ck(ispd_clk), .d(n_11509), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__u0 ( .ck(ispd_clk), .d(n_10423), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__u0 ( .ck(ispd_clk), .d(n_11507), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__u0 ( .ck(ispd_clk), .d(n_11505), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__u0 ( .ck(ispd_clk), .d(n_11503), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__u0 ( .ck(ispd_clk), .d(n_11502), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__u0 ( .ck(ispd_clk), .d(n_11500), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__u0 ( .ck(ispd_clk), .d(n_11499), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__u0 ( .ck(ispd_clk), .d(n_11497), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__u0 ( .ck(ispd_clk), .d(n_11496), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__u0 ( .ck(ispd_clk), .d(n_10421), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__u0 ( .ck(ispd_clk), .d(n_11495), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__u0 ( .ck(ispd_clk), .d(n_11493), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__u0 ( .ck(ispd_clk), .d(n_10419), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__u0 ( .ck(ispd_clk), .d(n_11492), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__u0 ( .ck(ispd_clk), .d(n_11490), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__u0 ( .ck(ispd_clk), .d(n_11489), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__u0 ( .ck(ispd_clk), .d(n_11487), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__u0 ( .ck(ispd_clk), .d(n_10418), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__u0 ( .ck(ispd_clk), .d(n_11485), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__u0 ( .ck(ispd_clk), .d(n_11484), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__u0 ( .ck(ispd_clk), .d(n_10829), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__u0 ( .ck(ispd_clk), .d(n_10828), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__u0 ( .ck(ispd_clk), .d(n_10366), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__u0 ( .ck(ispd_clk), .d(n_11710), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__u0 ( .ck(ispd_clk), .d(n_8959), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__u0 ( .ck(ispd_clk), .d(n_11483), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__u0 ( .ck(ispd_clk), .d(n_10417), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__u0 ( .ck(ispd_clk), .d(n_10416), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__u0 ( .ck(ispd_clk), .d(n_10414), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__u0 ( .ck(ispd_clk), .d(n_11482), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__u0 ( .ck(ispd_clk), .d(n_11480), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__u0 ( .ck(ispd_clk), .d(n_11479), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_0__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__u0 ( .ck(ispd_clk), .d(n_11698), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__u0 ( .ck(ispd_clk), .d(n_11697), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__u0 ( .ck(ispd_clk), .d(n_11696), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__u0 ( .ck(ispd_clk), .d(n_10515), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__u0 ( .ck(ispd_clk), .d(n_11695), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__u0 ( .ck(ispd_clk), .d(n_10513), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__u0 ( .ck(ispd_clk), .d(n_11694), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__u0 ( .ck(ispd_clk), .d(n_11693), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__u0 ( .ck(ispd_clk), .d(n_11692), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__u0 ( .ck(ispd_clk), .d(n_11691), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__u0 ( .ck(ispd_clk), .d(n_11690), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__u0 ( .ck(ispd_clk), .d(n_11689), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__u0 ( .ck(ispd_clk), .d(n_11688), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__u0 ( .ck(ispd_clk), .d(n_11687), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__u0 ( .ck(ispd_clk), .d(n_10511), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__u0 ( .ck(ispd_clk), .d(n_11686), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__u0 ( .ck(ispd_clk), .d(n_11685), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__u0 ( .ck(ispd_clk), .d(n_10509), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__u0 ( .ck(ispd_clk), .d(n_11684), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__u0 ( .ck(ispd_clk), .d(n_11683), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__u0 ( .ck(ispd_clk), .d(n_11682), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__u0 ( .ck(ispd_clk), .d(n_11681), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__u0 ( .ck(ispd_clk), .d(n_10508), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__u0 ( .ck(ispd_clk), .d(n_11680), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__u0 ( .ck(ispd_clk), .d(n_11679), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__u0 ( .ck(ispd_clk), .d(n_10848), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__u0 ( .ck(ispd_clk), .d(n_10847), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__u0 ( .ck(ispd_clk), .d(n_10506), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__u0 ( .ck(ispd_clk), .d(n_11708), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__u0 ( .ck(ispd_clk), .d(n_8916), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__u0 ( .ck(ispd_clk), .d(n_11677), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__u0 ( .ck(ispd_clk), .d(n_10503), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__u0 ( .ck(ispd_clk), .d(n_10501), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__u0 ( .ck(ispd_clk), .d(n_10499), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__u0 ( .ck(ispd_clk), .d(n_11676), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__u0 ( .ck(ispd_clk), .d(n_11675), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__u0 ( .ck(ispd_clk), .d(n_11674), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_10__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__u0 ( .ck(ispd_clk), .d(n_11336), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__u0 ( .ck(ispd_clk), .d(n_11334), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__u0 ( .ck(ispd_clk), .d(n_11332), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__u0 ( .ck(ispd_clk), .d(n_10365), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__u0 ( .ck(ispd_clk), .d(n_11330), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__u0 ( .ck(ispd_clk), .d(n_10363), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__u0 ( .ck(ispd_clk), .d(n_11328), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__u0 ( .ck(ispd_clk), .d(n_11327), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__u0 ( .ck(ispd_clk), .d(n_11324), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__u0 ( .ck(ispd_clk), .d(n_11326), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__u0 ( .ck(ispd_clk), .d(n_11322), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__u0 ( .ck(ispd_clk), .d(n_11320), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__u0 ( .ck(ispd_clk), .d(n_11318), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__u0 ( .ck(ispd_clk), .d(n_11316), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__u0 ( .ck(ispd_clk), .d(n_10362), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__u0 ( .ck(ispd_clk), .d(n_11314), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__u0 ( .ck(ispd_clk), .d(n_11311), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__u0 ( .ck(ispd_clk), .d(n_10361), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__u0 ( .ck(ispd_clk), .d(n_11309), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__u0 ( .ck(ispd_clk), .d(n_11307), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__u0 ( .ck(ispd_clk), .d(n_11306), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__u0 ( .ck(ispd_clk), .d(n_11305), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__u0 ( .ck(ispd_clk), .d(n_10359), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__u0 ( .ck(ispd_clk), .d(n_11303), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__u0 ( .ck(ispd_clk), .d(n_11302), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__u0 ( .ck(ispd_clk), .d(n_10823), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__u0 ( .ck(ispd_clk), .d(n_10821), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__u0 ( .ck(ispd_clk), .d(n_10357), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__u0 ( .ck(ispd_clk), .d(n_11300), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__u0 ( .ck(ispd_clk), .d(n_8955), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_11__465) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__u0 ( .ck(ispd_clk), .d(n_11297), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__u0 ( .ck(ispd_clk), .d(n_10355), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__u0 ( .ck(ispd_clk), .d(n_10353), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__u0 ( .ck(ispd_clk), .d(n_10351), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__u0 ( .ck(ispd_clk), .d(n_11295), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__u0 ( .ck(ispd_clk), .d(n_11293), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__u0 ( .ck(ispd_clk), .d(n_11290), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_11__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__u0 ( .ck(ispd_clk), .d(n_11672), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__u0 ( .ck(ispd_clk), .d(n_11671), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__u0 ( .ck(ispd_clk), .d(n_11670), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__u0 ( .ck(ispd_clk), .d(n_10497), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__u0 ( .ck(ispd_clk), .d(n_11669), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__u0 ( .ck(ispd_clk), .d(n_10495), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__u0 ( .ck(ispd_clk), .d(n_11668), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__u0 ( .ck(ispd_clk), .d(n_11667), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__u0 ( .ck(ispd_clk), .d(n_11666), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__u0 ( .ck(ispd_clk), .d(n_11665), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__u0 ( .ck(ispd_clk), .d(n_11663), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__u0 ( .ck(ispd_clk), .d(n_11662), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__u0 ( .ck(ispd_clk), .d(n_11660), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__u0 ( .ck(ispd_clk), .d(n_11661), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__u0 ( .ck(ispd_clk), .d(n_10493), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__u0 ( .ck(ispd_clk), .d(n_11659), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__u0 ( .ck(ispd_clk), .d(n_11657), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__u0 ( .ck(ispd_clk), .d(n_10491), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__u0 ( .ck(ispd_clk), .d(n_11655), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__u0 ( .ck(ispd_clk), .d(n_11653), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__u0 ( .ck(ispd_clk), .d(n_11652), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__u0 ( .ck(ispd_clk), .d(n_11651), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__u0 ( .ck(ispd_clk), .d(n_10489), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__u0 ( .ck(ispd_clk), .d(n_11650), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__u0 ( .ck(ispd_clk), .d(n_11648), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__u0 ( .ck(ispd_clk), .d(n_10845), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__u0 ( .ck(ispd_clk), .d(n_10843), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__u0 ( .ck(ispd_clk), .d(n_10487), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__u0 ( .ck(ispd_clk), .d(n_11707), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__u0 ( .ck(ispd_clk), .d(n_8914), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__u0 ( .ck(ispd_clk), .d(n_11647), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__u0 ( .ck(ispd_clk), .d(n_10485), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__u0 ( .ck(ispd_clk), .d(n_10483), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__u0 ( .ck(ispd_clk), .d(n_10481), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__u0 ( .ck(ispd_clk), .d(n_11645), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__u0 ( .ck(ispd_clk), .d(n_11644), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__u0 ( .ck(ispd_clk), .d(n_11642), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_12__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__u0 ( .ck(ispd_clk), .d(n_11289), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__u0 ( .ck(ispd_clk), .d(n_11287), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__u0 ( .ck(ispd_clk), .d(n_11286), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__u0 ( .ck(ispd_clk), .d(n_10349), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__u0 ( .ck(ispd_clk), .d(n_11285), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__u0 ( .ck(ispd_clk), .d(n_10348), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__u0 ( .ck(ispd_clk), .d(n_11284), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__u0 ( .ck(ispd_clk), .d(n_11283), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__u0 ( .ck(ispd_clk), .d(n_11282), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__u0 ( .ck(ispd_clk), .d(n_11281), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__u0 ( .ck(ispd_clk), .d(n_11280), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__u0 ( .ck(ispd_clk), .d(n_11279), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__u0 ( .ck(ispd_clk), .d(n_11277), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__u0 ( .ck(ispd_clk), .d(n_11276), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__u0 ( .ck(ispd_clk), .d(n_10346), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__u0 ( .ck(ispd_clk), .d(n_11274), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__u0 ( .ck(ispd_clk), .d(n_11273), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__u0 ( .ck(ispd_clk), .d(n_10344), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__u0 ( .ck(ispd_clk), .d(n_11271), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__u0 ( .ck(ispd_clk), .d(n_11270), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__u0 ( .ck(ispd_clk), .d(n_11268), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__u0 ( .ck(ispd_clk), .d(n_11266), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__u0 ( .ck(ispd_clk), .d(n_10343), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__u0 ( .ck(ispd_clk), .d(n_11265), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__u0 ( .ck(ispd_clk), .d(n_11264), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__u0 ( .ck(ispd_clk), .d(n_10820), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__u0 ( .ck(ispd_clk), .d(n_10819), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__u0 ( .ck(ispd_clk), .d(n_10342), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__u0 ( .ck(ispd_clk), .d(n_11262), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__u0 ( .ck(ispd_clk), .d(n_8900), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_13__543) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__u0 ( .ck(ispd_clk), .d(n_11261), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__u0 ( .ck(ispd_clk), .d(n_10340), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__u0 ( .ck(ispd_clk), .d(n_10338), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__u0 ( .ck(ispd_clk), .d(n_10336), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__u0 ( .ck(ispd_clk), .d(n_11260), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__u0 ( .ck(ispd_clk), .d(n_11259), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__u0 ( .ck(ispd_clk), .d(n_11258), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_13__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__u0 ( .ck(ispd_clk), .d(n_11256), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__u0 ( .ck(ispd_clk), .d(n_11255), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__u0 ( .ck(ispd_clk), .d(n_11254), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__u0 ( .ck(ispd_clk), .d(n_10334), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__u0 ( .ck(ispd_clk), .d(n_11252), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__u0 ( .ck(ispd_clk), .d(n_10332), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__u0 ( .ck(ispd_clk), .d(n_11251), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__u0 ( .ck(ispd_clk), .d(n_11250), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__u0 ( .ck(ispd_clk), .d(n_11249), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__u0 ( .ck(ispd_clk), .d(n_11247), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__u0 ( .ck(ispd_clk), .d(n_11246), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__u0 ( .ck(ispd_clk), .d(n_11245), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__u0 ( .ck(ispd_clk), .d(n_11244), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__u0 ( .ck(ispd_clk), .d(n_11243), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__u0 ( .ck(ispd_clk), .d(n_10331), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__u0 ( .ck(ispd_clk), .d(n_11242), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__u0 ( .ck(ispd_clk), .d(n_11241), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__u0 ( .ck(ispd_clk), .d(n_10329), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__u0 ( .ck(ispd_clk), .d(n_11240), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__u0 ( .ck(ispd_clk), .d(n_11239), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__u0 ( .ck(ispd_clk), .d(n_11238), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__u0 ( .ck(ispd_clk), .d(n_11236), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__u0 ( .ck(ispd_clk), .d(n_10327), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__u0 ( .ck(ispd_clk), .d(n_11235), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__u0 ( .ck(ispd_clk), .d(n_11234), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__u0 ( .ck(ispd_clk), .d(n_10817), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__u0 ( .ck(ispd_clk), .d(n_10815), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__u0 ( .ck(ispd_clk), .d(n_10325), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__u0 ( .ck(ispd_clk), .d(n_11232), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__u0 ( .ck(ispd_clk), .d(n_8899), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_14__582) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__u0 ( .ck(ispd_clk), .d(n_11230), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__u0 ( .ck(ispd_clk), .d(n_10323), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__u0 ( .ck(ispd_clk), .d(n_10321), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__u0 ( .ck(ispd_clk), .d(n_10319), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__u0 ( .ck(ispd_clk), .d(n_11229), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__u0 ( .ck(ispd_clk), .d(n_11228), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__u0 ( .ck(ispd_clk), .d(n_11226), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_14__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__u0 ( .ck(ispd_clk), .d(n_11224), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__u0 ( .ck(ispd_clk), .d(n_11223), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__u0 ( .ck(ispd_clk), .d(n_11222), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__u0 ( .ck(ispd_clk), .d(n_10317), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__u0 ( .ck(ispd_clk), .d(n_11220), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__u0 ( .ck(ispd_clk), .d(n_10316), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__u0 ( .ck(ispd_clk), .d(n_11219), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__u0 ( .ck(ispd_clk), .d(n_11218), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__u0 ( .ck(ispd_clk), .d(n_11217), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__u0 ( .ck(ispd_clk), .d(n_11216), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__u0 ( .ck(ispd_clk), .d(n_11215), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__u0 ( .ck(ispd_clk), .d(n_11214), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__u0 ( .ck(ispd_clk), .d(n_11213), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__u0 ( .ck(ispd_clk), .d(n_11212), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__u0 ( .ck(ispd_clk), .d(n_10314), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__u0 ( .ck(ispd_clk), .d(n_11211), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__u0 ( .ck(ispd_clk), .d(n_11209), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__u0 ( .ck(ispd_clk), .d(n_10312), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__u0 ( .ck(ispd_clk), .d(n_11208), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__u0 ( .ck(ispd_clk), .d(n_11207), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__u0 ( .ck(ispd_clk), .d(n_11206), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__u0 ( .ck(ispd_clk), .d(n_11205), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__u0 ( .ck(ispd_clk), .d(n_10311), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__u0 ( .ck(ispd_clk), .d(n_11203), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__u0 ( .ck(ispd_clk), .d(n_11202), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__u0 ( .ck(ispd_clk), .d(n_10813), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__u0 ( .ck(ispd_clk), .d(n_10812), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__u0 ( .ck(ispd_clk), .d(n_10310), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__u0 ( .ck(ispd_clk), .d(n_11200), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__u0 ( .ck(ispd_clk), .d(n_8898), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_15__621) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__u0 ( .ck(ispd_clk), .d(n_11198), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__u0 ( .ck(ispd_clk), .d(n_10308), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__u0 ( .ck(ispd_clk), .d(n_10306), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__u0 ( .ck(ispd_clk), .d(n_10304), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__u0 ( .ck(ispd_clk), .d(n_11196), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__u0 ( .ck(ispd_clk), .d(n_11194), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__u0 ( .ck(ispd_clk), .d(n_11193), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_15__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__u0 ( .ck(ispd_clk), .d(n_11478), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__u0 ( .ck(ispd_clk), .d(n_11477), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__u0 ( .ck(ispd_clk), .d(n_11476), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__u0 ( .ck(ispd_clk), .d(n_10413), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__u0 ( .ck(ispd_clk), .d(n_11474), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__u0 ( .ck(ispd_clk), .d(n_10412), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__u0 ( .ck(ispd_clk), .d(n_11473), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__u0 ( .ck(ispd_clk), .d(n_11472), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__u0 ( .ck(ispd_clk), .d(n_11470), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__u0 ( .ck(ispd_clk), .d(n_11468), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__u0 ( .ck(ispd_clk), .d(n_11467), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__u0 ( .ck(ispd_clk), .d(n_11466), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__u0 ( .ck(ispd_clk), .d(n_11464), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__u0 ( .ck(ispd_clk), .d(n_11463), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__u0 ( .ck(ispd_clk), .d(n_10411), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__u0 ( .ck(ispd_clk), .d(n_11462), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__u0 ( .ck(ispd_clk), .d(n_11460), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__u0 ( .ck(ispd_clk), .d(n_10410), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__u0 ( .ck(ispd_clk), .d(n_11458), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__u0 ( .ck(ispd_clk), .d(n_11457), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__u0 ( .ck(ispd_clk), .d(n_11456), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__u0 ( .ck(ispd_clk), .d(n_11454), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__u0 ( .ck(ispd_clk), .d(n_10408), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__u0 ( .ck(ispd_clk), .d(n_11451), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__u0 ( .ck(ispd_clk), .d(n_11452), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__u0 ( .ck(ispd_clk), .d(n_10810), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__u0 ( .ck(ispd_clk), .d(n_10807), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__u0 ( .ck(ispd_clk), .d(n_10302), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__u0 ( .ck(ispd_clk), .d(n_11706), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__u0 ( .ck(ispd_clk), .d(n_8912), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__u0 ( .ck(ispd_clk), .d(n_11449), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__u0 ( .ck(ispd_clk), .d(n_10407), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__u0 ( .ck(ispd_clk), .d(n_10405), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__u0 ( .ck(ispd_clk), .d(n_10404), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__u0 ( .ck(ispd_clk), .d(n_11446), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__u0 ( .ck(ispd_clk), .d(n_11445), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__u0 ( .ck(ispd_clk), .d(n_11443), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_1__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__u0 ( .ck(ispd_clk), .d(n_11442), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__u0 ( .ck(ispd_clk), .d(n_11441), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__u0 ( .ck(ispd_clk), .d(n_11440), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__u0 ( .ck(ispd_clk), .d(n_10402), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__u0 ( .ck(ispd_clk), .d(n_11438), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__u0 ( .ck(ispd_clk), .d(n_10401), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__u0 ( .ck(ispd_clk), .d(n_11437), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__u0 ( .ck(ispd_clk), .d(n_11436), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__u0 ( .ck(ispd_clk), .d(n_11435), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__u0 ( .ck(ispd_clk), .d(n_11431), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__u0 ( .ck(ispd_clk), .d(n_11434), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__u0 ( .ck(ispd_clk), .d(n_11433), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__u0 ( .ck(ispd_clk), .d(n_11432), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__u0 ( .ck(ispd_clk), .d(n_11429), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__u0 ( .ck(ispd_clk), .d(n_10400), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__u0 ( .ck(ispd_clk), .d(n_11427), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__u0 ( .ck(ispd_clk), .d(n_11425), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__u0 ( .ck(ispd_clk), .d(n_10399), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__u0 ( .ck(ispd_clk), .d(n_11424), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__u0 ( .ck(ispd_clk), .d(n_11423), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__u0 ( .ck(ispd_clk), .d(n_11421), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__u0 ( .ck(ispd_clk), .d(n_11420), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__u0 ( .ck(ispd_clk), .d(n_10397), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__u0 ( .ck(ispd_clk), .d(n_11419), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__u0 ( .ck(ispd_clk), .d(n_11418), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__u0 ( .ck(ispd_clk), .d(n_10806), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__u0 ( .ck(ispd_clk), .d(n_10804), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__u0 ( .ck(ispd_clk), .d(n_10300), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__u0 ( .ck(ispd_clk), .d(n_11705), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__u0 ( .ck(ispd_clk), .d(n_8910), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__u0 ( .ck(ispd_clk), .d(n_11417), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__u0 ( .ck(ispd_clk), .d(n_10396), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__u0 ( .ck(ispd_clk), .d(n_10394), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__u0 ( .ck(ispd_clk), .d(n_10393), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__u0 ( .ck(ispd_clk), .d(n_11415), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__u0 ( .ck(ispd_clk), .d(n_11414), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__u0 ( .ck(ispd_clk), .d(n_11413), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_2__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__u0 ( .ck(ispd_clk), .d(n_11641), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__u0 ( .ck(ispd_clk), .d(n_11640), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__u0 ( .ck(ispd_clk), .d(n_11639), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__u0 ( .ck(ispd_clk), .d(n_10479), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__u0 ( .ck(ispd_clk), .d(n_11638), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__u0 ( .ck(ispd_clk), .d(n_10478), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__u0 ( .ck(ispd_clk), .d(n_11637), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__u0 ( .ck(ispd_clk), .d(n_11635), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__u0 ( .ck(ispd_clk), .d(n_11634), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__u0 ( .ck(ispd_clk), .d(n_11631), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__u0 ( .ck(ispd_clk), .d(n_11633), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__u0 ( .ck(ispd_clk), .d(n_11632), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__u0 ( .ck(ispd_clk), .d(n_11630), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__u0 ( .ck(ispd_clk), .d(n_11628), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__u0 ( .ck(ispd_clk), .d(n_10477), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__u0 ( .ck(ispd_clk), .d(n_11626), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__u0 ( .ck(ispd_clk), .d(n_11625), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__u0 ( .ck(ispd_clk), .d(n_10476), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__u0 ( .ck(ispd_clk), .d(n_11624), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__u0 ( .ck(ispd_clk), .d(n_11623), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__u0 ( .ck(ispd_clk), .d(n_11622), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__u0 ( .ck(ispd_clk), .d(n_11620), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__u0 ( .ck(ispd_clk), .d(n_10474), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__u0 ( .ck(ispd_clk), .d(n_11618), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__u0 ( .ck(ispd_clk), .d(n_11617), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__u0 ( .ck(ispd_clk), .d(n_10841), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__u0 ( .ck(ispd_clk), .d(n_10839), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__u0 ( .ck(ispd_clk), .d(n_10473), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__u0 ( .ck(ispd_clk), .d(n_11712), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__u0 ( .ck(ispd_clk), .d(n_8908), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__u0 ( .ck(ispd_clk), .d(n_11616), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__u0 ( .ck(ispd_clk), .d(n_10469), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__u0 ( .ck(ispd_clk), .d(n_10470), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__u0 ( .ck(ispd_clk), .d(n_10467), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__u0 ( .ck(ispd_clk), .d(n_11614), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__u0 ( .ck(ispd_clk), .d(n_11613), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__u0 ( .ck(ispd_clk), .d(n_11611), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_3__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__u0 ( .ck(ispd_clk), .d(n_11411), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__u0 ( .ck(ispd_clk), .d(n_11410), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__u0 ( .ck(ispd_clk), .d(n_11408), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__u0 ( .ck(ispd_clk), .d(n_10391), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__u0 ( .ck(ispd_clk), .d(n_11406), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__u0 ( .ck(ispd_clk), .d(n_10390), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__u0 ( .ck(ispd_clk), .d(n_11405), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__u0 ( .ck(ispd_clk), .d(n_11403), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__u0 ( .ck(ispd_clk), .d(n_11402), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__u0 ( .ck(ispd_clk), .d(n_11401), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__Q) );
in01m20 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__18__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_4__213) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__u0 ( .ck(ispd_clk), .d(n_11399), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__u0 ( .ck(ispd_clk), .d(n_11398), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__u0 ( .ck(ispd_clk), .d(n_11396), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__u0 ( .ck(ispd_clk), .d(n_11394), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__u0 ( .ck(ispd_clk), .d(n_10388), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__u0 ( .ck(ispd_clk), .d(n_11393), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__u0 ( .ck(ispd_clk), .d(n_11391), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__u0 ( .ck(ispd_clk), .d(n_10386), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__u0 ( .ck(ispd_clk), .d(n_11390), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__u0 ( .ck(ispd_clk), .d(n_11388), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__u0 ( .ck(ispd_clk), .d(n_11386), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__u0 ( .ck(ispd_clk), .d(n_11385), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__u0 ( .ck(ispd_clk), .d(n_10385), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__u0 ( .ck(ispd_clk), .d(n_11384), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__u0 ( .ck(ispd_clk), .d(n_11383), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__u0 ( .ck(ispd_clk), .d(n_10803), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__u0 ( .ck(ispd_clk), .d(n_10802), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__u0 ( .ck(ispd_clk), .d(n_10298), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__u0 ( .ck(ispd_clk), .d(n_11703), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__u0 ( .ck(ispd_clk), .d(n_8906), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__u0 ( .ck(ispd_clk), .d(n_11382), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__u0 ( .ck(ispd_clk), .d(n_10384), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__u0 ( .ck(ispd_clk), .d(n_10383), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__u0 ( .ck(ispd_clk), .d(n_10381), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__u0 ( .ck(ispd_clk), .d(n_11381), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__u0 ( .ck(ispd_clk), .d(n_11380), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__u0 ( .ck(ispd_clk), .d(n_11379), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_4__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__u0 ( .ck(ispd_clk), .d(n_11610), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__u0 ( .ck(ispd_clk), .d(n_11609), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__u0 ( .ck(ispd_clk), .d(n_11607), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__u0 ( .ck(ispd_clk), .d(n_10465), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__u0 ( .ck(ispd_clk), .d(n_11606), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__u0 ( .ck(ispd_clk), .d(n_10464), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__u0 ( .ck(ispd_clk), .d(n_11605), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__u0 ( .ck(ispd_clk), .d(n_11604), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__u0 ( .ck(ispd_clk), .d(n_11603), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__u0 ( .ck(ispd_clk), .d(n_11602), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__u0 ( .ck(ispd_clk), .d(n_11601), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__u0 ( .ck(ispd_clk), .d(n_11600), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__u0 ( .ck(ispd_clk), .d(n_11599), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__u0 ( .ck(ispd_clk), .d(n_11598), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__u0 ( .ck(ispd_clk), .d(n_10463), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__u0 ( .ck(ispd_clk), .d(n_11597), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__u0 ( .ck(ispd_clk), .d(n_11595), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__u0 ( .ck(ispd_clk), .d(n_10462), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__u0 ( .ck(ispd_clk), .d(n_11593), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__u0 ( .ck(ispd_clk), .d(n_11592), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__u0 ( .ck(ispd_clk), .d(n_11590), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__u0 ( .ck(ispd_clk), .d(n_11589), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__u0 ( .ck(ispd_clk), .d(n_10460), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__u0 ( .ck(ispd_clk), .d(n_11588), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__u0 ( .ck(ispd_clk), .d(n_11587), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__u0 ( .ck(ispd_clk), .d(n_10838), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__u0 ( .ck(ispd_clk), .d(n_10836), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__u0 ( .ck(ispd_clk), .d(n_10459), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__u0 ( .ck(ispd_clk), .d(n_11702), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__u0 ( .ck(ispd_clk), .d(n_8904), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__u0 ( .ck(ispd_clk), .d(n_11586), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__u0 ( .ck(ispd_clk), .d(n_10457), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__u0 ( .ck(ispd_clk), .d(n_10455), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__u0 ( .ck(ispd_clk), .d(n_10453), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__u0 ( .ck(ispd_clk), .d(n_11585), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__u0 ( .ck(ispd_clk), .d(n_11584), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__u0 ( .ck(ispd_clk), .d(n_11583), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_5__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__u0 ( .ck(ispd_clk), .d(n_11582), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__u0 ( .ck(ispd_clk), .d(n_11580), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__u0 ( .ck(ispd_clk), .d(n_11579), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__u0 ( .ck(ispd_clk), .d(n_10451), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__u0 ( .ck(ispd_clk), .d(n_11577), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__u0 ( .ck(ispd_clk), .d(n_10450), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__u0 ( .ck(ispd_clk), .d(n_11575), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__u0 ( .ck(ispd_clk), .d(n_11573), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__u0 ( .ck(ispd_clk), .d(n_11572), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__u0 ( .ck(ispd_clk), .d(n_11571), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__Q) );
in01s02 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__18__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_6__252) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__u0 ( .ck(ispd_clk), .d(n_11570), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__u0 ( .ck(ispd_clk), .d(n_11568), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__u0 ( .ck(ispd_clk), .d(n_11566), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__u0 ( .ck(ispd_clk), .d(n_11565), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__u0 ( .ck(ispd_clk), .d(n_10449), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__u0 ( .ck(ispd_clk), .d(n_11564), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__u0 ( .ck(ispd_clk), .d(n_11562), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__u0 ( .ck(ispd_clk), .d(n_10447), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__u0 ( .ck(ispd_clk), .d(n_11561), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__u0 ( .ck(ispd_clk), .d(n_11560), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__u0 ( .ck(ispd_clk), .d(n_11559), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__u0 ( .ck(ispd_clk), .d(n_11557), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__u0 ( .ck(ispd_clk), .d(n_10446), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__u0 ( .ck(ispd_clk), .d(n_11556), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__u0 ( .ck(ispd_clk), .d(n_11555), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__u0 ( .ck(ispd_clk), .d(n_10835), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__u0 ( .ck(ispd_clk), .d(n_10834), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__u0 ( .ck(ispd_clk), .d(n_10445), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__u0 ( .ck(ispd_clk), .d(n_11701), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__u0 ( .ck(ispd_clk), .d(n_8902), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__u0 ( .ck(ispd_clk), .d(n_11553), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__u0 ( .ck(ispd_clk), .d(n_10444), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__u0 ( .ck(ispd_clk), .d(n_10443), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__u0 ( .ck(ispd_clk), .d(n_10440), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__u0 ( .ck(ispd_clk), .d(n_11551), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__u0 ( .ck(ispd_clk), .d(n_11549), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__u0 ( .ck(ispd_clk), .d(n_11548), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_6__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__u0 ( .ck(ispd_clk), .d(n_11191), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__u0 ( .ck(ispd_clk), .d(n_11190), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__u0 ( .ck(ispd_clk), .d(n_11188), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__u0 ( .ck(ispd_clk), .d(n_10297), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__u0 ( .ck(ispd_clk), .d(n_11187), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__u0 ( .ck(ispd_clk), .d(n_10296), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__u0 ( .ck(ispd_clk), .d(n_11186), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__u0 ( .ck(ispd_clk), .d(n_11184), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__u0 ( .ck(ispd_clk), .d(n_11182), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__u0 ( .ck(ispd_clk), .d(n_11181), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__Q) );
in01s02 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__18__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__291) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__u0 ( .ck(ispd_clk), .d(n_11180), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__u0 ( .ck(ispd_clk), .d(n_11179), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__u0 ( .ck(ispd_clk), .d(n_11178), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__u0 ( .ck(ispd_clk), .d(n_11177), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__u0 ( .ck(ispd_clk), .d(n_10294), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__u0 ( .ck(ispd_clk), .d(n_11175), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__u0 ( .ck(ispd_clk), .d(n_11174), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__u0 ( .ck(ispd_clk), .d(n_10292), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__u0 ( .ck(ispd_clk), .d(n_11173), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__u0 ( .ck(ispd_clk), .d(n_11171), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__u0 ( .ck(ispd_clk), .d(n_11169), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__u0 ( .ck(ispd_clk), .d(n_11167), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__u0 ( .ck(ispd_clk), .d(n_10291), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__u0 ( .ck(ispd_clk), .d(n_11165), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__u0 ( .ck(ispd_clk), .d(n_11337), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__u0 ( .ck(ispd_clk), .d(n_10800), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__u0 ( .ck(ispd_clk), .d(n_10799), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__u0 ( .ck(ispd_clk), .d(n_10290), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__u0 ( .ck(ispd_clk), .d(n_11164), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__u0 ( .ck(ispd_clk), .d(n_9188), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__Q) );
in01s01 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__u1 ( .a(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__36__Q), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_7__309) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__u0 ( .ck(ispd_clk), .d(n_11162), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__u0 ( .ck(ispd_clk), .d(n_10289), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__u0 ( .ck(ispd_clk), .d(n_10288), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__u0 ( .ck(ispd_clk), .d(n_10286), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__u0 ( .ck(ispd_clk), .d(n_11161), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__u0 ( .ck(ispd_clk), .d(n_11159), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__u0 ( .ck(ispd_clk), .d(n_11158), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_7__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__u0 ( .ck(ispd_clk), .d(n_11377), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__u0 ( .ck(ispd_clk), .d(n_11375), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__u0 ( .ck(ispd_clk), .d(n_11373), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__u0 ( .ck(ispd_clk), .d(n_10380), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__u0 ( .ck(ispd_clk), .d(n_11372), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__u0 ( .ck(ispd_clk), .d(n_10378), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__u0 ( .ck(ispd_clk), .d(n_11370), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__u0 ( .ck(ispd_clk), .d(n_11369), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__u0 ( .ck(ispd_clk), .d(n_11367), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__u0 ( .ck(ispd_clk), .d(n_11365), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__u0 ( .ck(ispd_clk), .d(n_11363), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__u0 ( .ck(ispd_clk), .d(n_11362), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__u0 ( .ck(ispd_clk), .d(n_11361), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__u0 ( .ck(ispd_clk), .d(n_11359), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__u0 ( .ck(ispd_clk), .d(n_10377), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__u0 ( .ck(ispd_clk), .d(n_11357), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__u0 ( .ck(ispd_clk), .d(n_11355), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__u0 ( .ck(ispd_clk), .d(n_10376), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__u0 ( .ck(ispd_clk), .d(n_11353), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__u0 ( .ck(ispd_clk), .d(n_11352), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__u0 ( .ck(ispd_clk), .d(n_11350), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__u0 ( .ck(ispd_clk), .d(n_11349), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__u0 ( .ck(ispd_clk), .d(n_10374), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__u0 ( .ck(ispd_clk), .d(n_11347), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__u0 ( .ck(ispd_clk), .d(n_11345), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__u0 ( .ck(ispd_clk), .d(n_10797), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__u0 ( .ck(ispd_clk), .d(n_10795), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__u0 ( .ck(ispd_clk), .d(n_10285), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__u0 ( .ck(ispd_clk), .d(n_11700), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__u0 ( .ck(ispd_clk), .d(n_8957), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__u0 ( .ck(ispd_clk), .d(n_11344), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__u0 ( .ck(ispd_clk), .d(n_10372), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__u0 ( .ck(ispd_clk), .d(n_10370), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__u0 ( .ck(ispd_clk), .d(n_10368), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__u0 ( .ck(ispd_clk), .d(n_11342), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__u0 ( .ck(ispd_clk), .d(n_11340), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__u0 ( .ck(ispd_clk), .d(n_11338), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_8__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__u0 ( .ck(ispd_clk), .d(n_11547), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__0__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__u0 ( .ck(ispd_clk), .d(n_11546), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__10__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__u0 ( .ck(ispd_clk), .d(n_11545), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__11__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__u0 ( .ck(ispd_clk), .d(n_10439), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__12__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__u0 ( .ck(ispd_clk), .d(n_11544), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__13__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__u0 ( .ck(ispd_clk), .d(n_10438), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__14__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__u0 ( .ck(ispd_clk), .d(n_11543), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__15__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__u0 ( .ck(ispd_clk), .d(n_11542), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__16__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__u0 ( .ck(ispd_clk), .d(n_11540), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__17__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__u0 ( .ck(ispd_clk), .d(n_11538), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__18__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__u0 ( .ck(ispd_clk), .d(n_11536), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__19__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__u0 ( .ck(ispd_clk), .d(n_11535), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__1__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__u0 ( .ck(ispd_clk), .d(n_11534), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__20__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__u0 ( .ck(ispd_clk), .d(n_11533), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__21__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__u0 ( .ck(ispd_clk), .d(n_10436), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__22__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__u0 ( .ck(ispd_clk), .d(n_11532), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__23__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__u0 ( .ck(ispd_clk), .d(n_11531), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__24__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__u0 ( .ck(ispd_clk), .d(n_10434), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__25__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__u0 ( .ck(ispd_clk), .d(n_11530), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__26__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__u0 ( .ck(ispd_clk), .d(n_11528), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__27__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__u0 ( .ck(ispd_clk), .d(n_11526), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__28__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__u0 ( .ck(ispd_clk), .d(n_11524), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__29__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__u0 ( .ck(ispd_clk), .d(n_10433), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__u0 ( .ck(ispd_clk), .d(n_11521), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__30__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__u0 ( .ck(ispd_clk), .d(n_11523), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__31__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__u0 ( .ck(ispd_clk), .d(n_10833), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__32__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__u0 ( .ck(ispd_clk), .d(n_10832), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__33__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__u0 ( .ck(ispd_clk), .d(n_10432), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__34__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__u0 ( .ck(ispd_clk), .d(n_11699), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__35__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__u0 ( .ck(ispd_clk), .d(n_9191), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__36__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__u0 ( .ck(ispd_clk), .d(n_11519), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__3__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__u0 ( .ck(ispd_clk), .d(n_10430), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__4__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__u0 ( .ck(ispd_clk), .d(n_10428), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__5__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__u0 ( .ck(ispd_clk), .d(n_10426), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__6__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__u0 ( .ck(ispd_clk), .d(n_11517), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__7__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__u0 ( .ck(ispd_clk), .d(n_11516), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__8__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__u0 ( .ck(ispd_clk), .d(n_11515), .o(wishbone_slave_unit_fifos_wbw_fifo_storage_mem_reg_9__9__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__u0 ( .ck(ispd_clk), .d(n_8917), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__Q) );
in01s40 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_0__Q), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__u0 ( .ck(ispd_clk), .d(n_9146), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__Q) );
in01s40 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_1__Q), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__u0 ( .ck(ispd_clk), .d(n_8921), .o(wishbone_slave_unit_fifos_wbw_inTransactionCount_reg_2__Q) );
ms00f80 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__u0 ( .ck(ispd_clk), .d(n_8588), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__Q) );
in01f20 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__u1 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_0__Q), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_0_) );
ms00f80 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__u0 ( .ck(ispd_clk), .d(n_8669), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__Q) );
in01m40 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__u1 ( .a(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_1__Q), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_1_) );
ms00f80 wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__u0 ( .ck(ispd_clk), .d(n_8591), .o(wishbone_slave_unit_fifos_wbw_outTransactionCount_reg_2__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_bc_out_reg_0__u0 ( .ck(ispd_clk), .d(n_13499), .o(conf_wb_err_bc_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_bc_out_reg_1__u0 ( .ck(ispd_clk), .d(n_7714), .o(conf_wb_err_bc_in_846) );
ms00f80 wishbone_slave_unit_pci_initiator_if_bc_out_reg_2__u0 ( .ck(ispd_clk), .d(n_13502), .o(conf_wb_err_bc_in_847) );
ms00f80 wishbone_slave_unit_pci_initiator_if_bc_out_reg_3__u0 ( .ck(ispd_clk), .d(n_13500), .o(conf_wb_err_bc_in_848) );
ms00f80 wishbone_slave_unit_pci_initiator_if_be_out_reg_0__u0 ( .ck(ispd_clk), .d(n_13824), .o(n_1111) );
ms00f80 wishbone_slave_unit_pci_initiator_if_be_out_reg_1__u0 ( .ck(ispd_clk), .d(n_7212), .o(wishbone_slave_unit_pcim_sm_be_in_557) );
ms00f80 wishbone_slave_unit_pci_initiator_if_be_out_reg_2__u0 ( .ck(ispd_clk), .d(n_13827), .o(wishbone_slave_unit_pcim_sm_be_in_558) );
ms00f80 wishbone_slave_unit_pci_initiator_if_be_out_reg_3__u0 ( .ck(ispd_clk), .d(n_13826), .o(wishbone_slave_unit_pcim_sm_be_in_559) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_byte_address_reg_0__u0 ( .ck(ispd_clk), .d(n_13497), .o(wishbone_slave_unit_pci_initiator_if_current_byte_address) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_byte_address_reg_1__u0 ( .ck(ispd_clk), .d(n_13496), .o(wishbone_slave_unit_pci_initiator_if_current_byte_address_36) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_0__u0 ( .ck(ispd_clk), .d(n_13556), .o(conf_wb_err_addr_in_943) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_10__u0 ( .ck(ispd_clk), .d(n_13512), .o(conf_wb_err_addr_in_953) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_11__u0 ( .ck(ispd_clk), .d(n_13511), .o(conf_wb_err_addr_in_954) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_12__u0 ( .ck(ispd_clk), .d(n_13648), .o(conf_wb_err_addr_in_955) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_13__u0 ( .ck(ispd_clk), .d(n_13509), .o(conf_wb_err_addr_in_956) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_14__u0 ( .ck(ispd_clk), .d(n_13647), .o(conf_wb_err_addr_in_957) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_15__u0 ( .ck(ispd_clk), .d(n_13508), .o(conf_wb_err_addr_in_958) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_16__u0 ( .ck(ispd_clk), .d(n_13552), .o(conf_wb_err_addr_in_959) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_17__u0 ( .ck(ispd_clk), .d(n_13646), .o(conf_wb_err_addr_in_960) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_18__u0 ( .ck(ispd_clk), .d(n_13645), .o(conf_wb_err_addr_in_961) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_19__u0 ( .ck(ispd_clk), .d(n_13559), .o(conf_wb_err_addr_in_962) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_1__u0 ( .ck(ispd_clk), .d(n_13506), .o(conf_wb_err_addr_in_944) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_20__u0 ( .ck(ispd_clk), .d(n_13643), .o(conf_wb_err_addr_in_963) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_21__u0 ( .ck(ispd_clk), .d(n_13642), .o(conf_wb_err_addr_in_964) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_22__u0 ( .ck(ispd_clk), .d(n_13641), .o(conf_wb_err_addr_in_965) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_23__u0 ( .ck(ispd_clk), .d(n_13558), .o(conf_wb_err_addr_in_966) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_24__u0 ( .ck(ispd_clk), .d(n_13695), .o(conf_wb_err_addr_in_967) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_25__u0 ( .ck(ispd_clk), .d(n_13640), .o(conf_wb_err_addr_in_968) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_26__u0 ( .ck(ispd_clk), .d(n_13638), .o(conf_wb_err_addr_in_969) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_27__u0 ( .ck(ispd_clk), .d(n_13636), .o(conf_wb_err_addr_in_970) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_28__u0 ( .ck(ispd_clk), .d(n_13557), .o(conf_wb_err_addr_in_971) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__u0 ( .ck(ispd_clk), .d(n_13635), .o(wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_29__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_2__u0 ( .ck(ispd_clk), .d(n_13634), .o(conf_wb_err_addr_in_945) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_3__u0 ( .ck(ispd_clk), .d(n_13632), .o(conf_wb_err_addr_in_946) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_4__u0 ( .ck(ispd_clk), .d(n_13631), .o(conf_wb_err_addr_in_947) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_5__u0 ( .ck(ispd_clk), .d(n_13629), .o(conf_wb_err_addr_in_948) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_6__u0 ( .ck(ispd_clk), .d(n_13505), .o(conf_wb_err_addr_in_949) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_7__u0 ( .ck(ispd_clk), .d(n_13628), .o(conf_wb_err_addr_in_950) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_8__u0 ( .ck(ispd_clk), .d(n_13504), .o(conf_wb_err_addr_in_951) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_dword_address_reg_9__u0 ( .ck(ispd_clk), .d(n_13503), .o(conf_wb_err_addr_in_952) );
ms00f80 wishbone_slave_unit_pci_initiator_if_current_last_reg_u0 ( .ck(ispd_clk), .d(n_7539), .o(wishbone_slave_unit_pcim_sm_last_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_0__u0 ( .ck(ispd_clk), .d(n_7783), .o(wishbone_slave_unit_pcim_sm_data_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_10__u0 ( .ck(ispd_clk), .d(n_7782), .o(wishbone_slave_unit_pcim_sm_data_in_644) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_11__u0 ( .ck(ispd_clk), .d(n_7781), .o(wishbone_slave_unit_pcim_sm_data_in_645) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_12__u0 ( .ck(ispd_clk), .d(n_7780), .o(wishbone_slave_unit_pcim_sm_data_in_646) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_13__u0 ( .ck(ispd_clk), .d(n_7779), .o(wishbone_slave_unit_pcim_sm_data_in_647) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_14__u0 ( .ck(ispd_clk), .d(n_7777), .o(wishbone_slave_unit_pcim_sm_data_in_648) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_15__u0 ( .ck(ispd_clk), .d(n_7776), .o(wishbone_slave_unit_pcim_sm_data_in_649) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_16__u0 ( .ck(ispd_clk), .d(n_7774), .o(wishbone_slave_unit_pcim_sm_data_in_650) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_17__u0 ( .ck(ispd_clk), .d(n_7773), .o(wishbone_slave_unit_pcim_sm_data_in_651) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_18__u0 ( .ck(ispd_clk), .d(n_7771), .o(wishbone_slave_unit_pcim_sm_data_in_652) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_19__u0 ( .ck(ispd_clk), .d(n_7769), .o(wishbone_slave_unit_pcim_sm_data_in_653) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_1__u0 ( .ck(ispd_clk), .d(n_7768), .o(wishbone_slave_unit_pcim_sm_data_in_635) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_20__u0 ( .ck(ispd_clk), .d(n_7767), .o(wishbone_slave_unit_pcim_sm_data_in_654) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_21__u0 ( .ck(ispd_clk), .d(n_7766), .o(wishbone_slave_unit_pcim_sm_data_in_655) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_22__u0 ( .ck(ispd_clk), .d(n_7764), .o(wishbone_slave_unit_pcim_sm_data_in_656) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_23__u0 ( .ck(ispd_clk), .d(n_7762), .o(wishbone_slave_unit_pcim_sm_data_in_657) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_24__u0 ( .ck(ispd_clk), .d(n_7761), .o(wishbone_slave_unit_pcim_sm_data_in_658) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_25__u0 ( .ck(ispd_clk), .d(n_7760), .o(wishbone_slave_unit_pcim_sm_data_in_659) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_26__u0 ( .ck(ispd_clk), .d(n_7759), .o(wishbone_slave_unit_pcim_sm_data_in_660) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_27__u0 ( .ck(ispd_clk), .d(n_7757), .o(wishbone_slave_unit_pcim_sm_data_in_661) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_28__u0 ( .ck(ispd_clk), .d(n_7756), .o(wishbone_slave_unit_pcim_sm_data_in_662) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_29__u0 ( .ck(ispd_clk), .d(n_7755), .o(wishbone_slave_unit_pcim_sm_data_in_663) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_2__u0 ( .ck(ispd_clk), .d(n_7754), .o(wishbone_slave_unit_pcim_sm_data_in_636) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_30__u0 ( .ck(ispd_clk), .d(n_7753), .o(wishbone_slave_unit_pcim_sm_data_in_664) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_31__u0 ( .ck(ispd_clk), .d(n_7752), .o(wishbone_slave_unit_pcim_sm_data_in_665) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_3__u0 ( .ck(ispd_clk), .d(n_7751), .o(wishbone_slave_unit_pcim_sm_data_in_637) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_4__u0 ( .ck(ispd_clk), .d(n_7750), .o(wishbone_slave_unit_pcim_sm_data_in_638) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_5__u0 ( .ck(ispd_clk), .d(n_7749), .o(wishbone_slave_unit_pcim_sm_data_in_639) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_6__u0 ( .ck(ispd_clk), .d(n_7747), .o(wishbone_slave_unit_pcim_sm_data_in_640) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_7__u0 ( .ck(ispd_clk), .d(n_7746), .o(wishbone_slave_unit_pcim_sm_data_in_641) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_8__u0 ( .ck(ispd_clk), .d(n_7745), .o(wishbone_slave_unit_pcim_sm_data_in_642) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_out_reg_9__u0 ( .ck(ispd_clk), .d(n_7744), .o(wishbone_slave_unit_pcim_sm_data_in_643) );
ms00f80 wishbone_slave_unit_pci_initiator_if_data_source_reg_u0 ( .ck(ispd_clk), .d(n_4884), .o(wishbone_slave_unit_pci_initiator_if_data_source) );
ms00f80 wishbone_slave_unit_pci_initiator_if_del_read_req_reg_u0 ( .ck(ispd_clk), .d(n_8535), .o(wishbone_slave_unit_pci_initiator_if_del_read_req) );
ms00f80 wishbone_slave_unit_pci_initiator_if_del_write_req_reg_u0 ( .ck(ispd_clk), .d(n_4693), .o(wishbone_slave_unit_pci_initiator_if_del_write_req) );
ms00f80 wishbone_slave_unit_pci_initiator_if_err_recovery_reg_u0 ( .ck(ispd_clk), .d(n_7300), .o(wishbone_slave_unit_pci_initiator_if_err_recovery) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__u0 ( .ck(ispd_clk), .d(n_13550), .o(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_0__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__u0 ( .ck(ispd_clk), .d(n_7621), .o(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_1__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__u0 ( .ck(ispd_clk), .d(n_13546), .o(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_2__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__u0 ( .ck(ispd_clk), .d(n_13543), .o(wishbone_slave_unit_pci_initiator_if_intermediate_be_reg_3__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__u0 ( .ck(ispd_clk), .d(n_13540), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_0__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__u0 ( .ck(ispd_clk), .d(n_13539), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_10__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__u0 ( .ck(ispd_clk), .d(n_13538), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_11__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__u0 ( .ck(ispd_clk), .d(n_13537), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_12__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__u0 ( .ck(ispd_clk), .d(n_13536), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_13__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__u0 ( .ck(ispd_clk), .d(n_13535), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_14__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__u0 ( .ck(ispd_clk), .d(n_13534), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_15__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__u0 ( .ck(ispd_clk), .d(n_13533), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_16__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__u0 ( .ck(ispd_clk), .d(n_13532), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_17__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__u0 ( .ck(ispd_clk), .d(n_13531), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_18__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__u0 ( .ck(ispd_clk), .d(n_13530), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_19__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__u0 ( .ck(ispd_clk), .d(n_13529), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_1__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__u0 ( .ck(ispd_clk), .d(n_13528), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_20__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__u0 ( .ck(ispd_clk), .d(n_13470), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_21__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__u0 ( .ck(ispd_clk), .d(n_13527), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_22__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__u0 ( .ck(ispd_clk), .d(n_13526), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_23__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__u0 ( .ck(ispd_clk), .d(n_13525), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_24__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__u0 ( .ck(ispd_clk), .d(n_13469), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_25__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__u0 ( .ck(ispd_clk), .d(n_13627), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_26__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__u0 ( .ck(ispd_clk), .d(n_13524), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_27__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__u0 ( .ck(ispd_clk), .d(n_13523), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_28__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__u0 ( .ck(ispd_clk), .d(n_13522), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_29__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__u0 ( .ck(ispd_clk), .d(n_13521), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_2__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__u0 ( .ck(ispd_clk), .d(n_13468), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_30__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__u0 ( .ck(ispd_clk), .d(n_13520), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_31__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__u0 ( .ck(ispd_clk), .d(n_13519), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_3__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__u0 ( .ck(ispd_clk), .d(n_13518), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_4__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__u0 ( .ck(ispd_clk), .d(n_13517), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_5__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__u0 ( .ck(ispd_clk), .d(n_13516), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_6__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__u0 ( .ck(ispd_clk), .d(n_13515), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_7__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__u0 ( .ck(ispd_clk), .d(n_13514), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_8__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__u0 ( .ck(ispd_clk), .d(n_13513), .o(wishbone_slave_unit_pci_initiator_if_intermediate_data_reg_9__Q) );
ms00f80 wishbone_slave_unit_pci_initiator_if_intermediate_last_reg_u0 ( .ck(ispd_clk), .d(n_7625), .o(n_16763) );
ms00f80 wishbone_slave_unit_pci_initiator_if_last_transfered_reg_u0 ( .ck(ispd_clk), .d(n_3081), .o(wishbone_slave_unit_fifos_wbr_control_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_posted_write_req_reg_u0 ( .ck(ispd_clk), .d(n_7028), .o(wishbone_slave_unit_pci_initiator_if_posted_write_req) );
ms00f80 wishbone_slave_unit_pci_initiator_if_rdy_out_reg_u0 ( .ck(ispd_clk), .d(n_2801), .o(wishbone_slave_unit_pcim_sm_rdy_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_bound_reg_u0 ( .ck(ispd_clk), .d(n_4870), .o(wishbone_slave_unit_pci_initiator_if_read_bound) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_count_reg_0__u0 ( .ck(ispd_clk), .d(n_4861), .o(wishbone_slave_unit_pci_initiator_if_read_count_0_) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_count_reg_1__u0 ( .ck(ispd_clk), .d(n_4860), .o(wishbone_slave_unit_pci_initiator_if_read_count_1_) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_count_reg_2__u0 ( .ck(ispd_clk), .d(n_7333), .o(wishbone_slave_unit_pci_initiator_if_read_count_2_) );
ms00f80 wishbone_slave_unit_pci_initiator_if_read_count_reg_3__u0 ( .ck(ispd_clk), .d(n_7544), .o(wishbone_slave_unit_pci_initiator_if_read_count_reg_3__Q) );
in01s04 wishbone_slave_unit_pci_initiator_if_read_count_reg_3__u1 ( .a(wishbone_slave_unit_pci_initiator_if_read_count_reg_3__Q), .o(wishbone_slave_unit_pci_initiator_if_read_count_3_) );
ms00f80 wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_u0 ( .ck(ispd_clk), .d(n_3119), .o(wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_Q) );
in01s01 wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_u1 ( .a(wishbone_slave_unit_pci_initiator_if_tabort_received_out_reg_Q), .o(conf_target_abort_recv_in) );
ms00f80 wishbone_slave_unit_pci_initiator_if_write_req_int_reg_u0 ( .ck(ispd_clk), .d(n_15859), .o(wishbone_slave_unit_pci_initiator_if_write_req_int) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_cur_state_reg_0__u0 ( .ck(ispd_clk), .d(n_7617), .o(wishbone_slave_unit_pci_initiator_sm_cur_state_0_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_cur_state_reg_1__u0 ( .ck(ispd_clk), .d(n_7616), .o(wishbone_slave_unit_pci_initiator_sm_cur_state_1_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_cur_state_reg_2__u0 ( .ck(ispd_clk), .d(n_7620), .o(wishbone_slave_unit_pci_initiator_sm_cur_state_2_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_cur_state_reg_3__u0 ( .ck(ispd_clk), .d(n_7619), .o(wishbone_slave_unit_pci_initiator_sm_cur_state_3_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_decode_count_reg_0__u0 ( .ck(ispd_clk), .d(n_4537), .o(wishbone_slave_unit_pci_initiator_sm_decode_count_0_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_decode_count_reg_1__u0 ( .ck(ispd_clk), .d(n_4534), .o(wishbone_slave_unit_pci_initiator_sm_decode_count_1_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_decode_count_reg_2__u0 ( .ck(ispd_clk), .d(n_4746), .o(wishbone_slave_unit_pci_initiator_sm_decode_count_2_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_0__u0 ( .ck(ispd_clk), .d(n_6982), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_0_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_1__u0 ( .ck(ispd_clk), .d(n_6984), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_1_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_2__u0 ( .ck(ispd_clk), .d(n_6987), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_2_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_3__u0 ( .ck(ispd_clk), .d(n_5748), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_3_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_4__u0 ( .ck(ispd_clk), .d(n_5644), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_4_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_5__u0 ( .ck(ispd_clk), .d(n_6985), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_5_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_6__u0 ( .ck(ispd_clk), .d(n_5713), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_6_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_latency_timer_reg_7__u0 ( .ck(ispd_clk), .d(n_4892), .o(wishbone_slave_unit_pci_initiator_sm_latency_timer_7_) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_mabort1_reg_u0 ( .ck(ispd_clk), .d(n_2684), .o(wishbone_slave_unit_pci_initiator_sm_mabort1) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_mabort2_reg_u0 ( .ck(ispd_clk), .d(wishbone_slave_unit_pci_initiator_sm_mabort1), .o(wishbone_slave_unit_pci_initiator_sm_mabort2) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg_0__u0 ( .ck(ispd_clk), .d(n_7615), .o(wishbone_slave_unit_pci_initiator_sm_rdata_selector) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_rdata_selector_reg_1__u0 ( .ck(ispd_clk), .d(n_7614), .o(wishbone_slave_unit_pci_initiator_sm_rdata_selector_14) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_timeout_reg_u0 ( .ck(ispd_clk), .d(n_4679), .o(wishbone_slave_unit_pci_initiator_sm_timeout) );
ms00f80 wishbone_slave_unit_pci_initiator_sm_transfer_reg_u0 ( .ck(ispd_clk), .d(n_3812), .o(wishbone_slave_unit_pci_initiator_sm_transfer) );
ms00f80 wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_u0 ( .ck(ispd_clk), .d(n_14483), .o(wishbone_slave_unit_wishbone_slave_async_reset_as_wbr_flush_async_reset_data_out_reg_Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_c_state_reg_0__u0 ( .ck(ispd_clk), .d(n_14628), .o(wishbone_slave_unit_wishbone_slave_c_state) );
ms00f80 wishbone_slave_unit_wishbone_slave_c_state_reg_1__u0 ( .ck(ispd_clk), .d(n_7330), .o(wishbone_slave_unit_wishbone_slave_c_state_1) );
ms00f80 wishbone_slave_unit_wishbone_slave_c_state_reg_2__u0 ( .ck(ispd_clk), .d(n_14619), .o(wishbone_slave_unit_wishbone_slave_c_state_2) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__u0 ( .ck(ispd_clk), .d(n_8641), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_0__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__u0 ( .ck(ispd_clk), .d(n_8640), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_10__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__u0 ( .ck(ispd_clk), .d(n_8638), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_11__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__u0 ( .ck(ispd_clk), .d(n_8637), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_12__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__u0 ( .ck(ispd_clk), .d(n_8636), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_13__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__u0 ( .ck(ispd_clk), .d(n_8635), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_14__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__u0 ( .ck(ispd_clk), .d(n_8634), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_15__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__u0 ( .ck(ispd_clk), .d(n_8633), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_16__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__u0 ( .ck(ispd_clk), .d(n_8632), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_17__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__u0 ( .ck(ispd_clk), .d(n_8631), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_18__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__u0 ( .ck(ispd_clk), .d(n_8630), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_19__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__u0 ( .ck(ispd_clk), .d(n_8629), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_1__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__u0 ( .ck(ispd_clk), .d(n_8628), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_20__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__u0 ( .ck(ispd_clk), .d(n_8627), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_21__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__u0 ( .ck(ispd_clk), .d(n_8626), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_22__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__u0 ( .ck(ispd_clk), .d(n_8625), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_23__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__u0 ( .ck(ispd_clk), .d(n_8624), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_24__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__u0 ( .ck(ispd_clk), .d(n_8623), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_25__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__u0 ( .ck(ispd_clk), .d(n_8622), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_26__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__u0 ( .ck(ispd_clk), .d(n_8621), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_27__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__u0 ( .ck(ispd_clk), .d(n_8620), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_28__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__u0 ( .ck(ispd_clk), .d(n_8619), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_29__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__u0 ( .ck(ispd_clk), .d(n_8618), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_2__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__u0 ( .ck(ispd_clk), .d(n_8617), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_30__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__u0 ( .ck(ispd_clk), .d(n_8616), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_31__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__u0 ( .ck(ispd_clk), .d(n_8615), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_32__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__u0 ( .ck(ispd_clk), .d(n_8613), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_33__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__u0 ( .ck(ispd_clk), .d(n_8611), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_34__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__u0 ( .ck(ispd_clk), .d(n_8609), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_35__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__u0 ( .ck(ispd_clk), .d(n_8607), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_3__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__u0 ( .ck(ispd_clk), .d(n_8606), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_4__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__u0 ( .ck(ispd_clk), .d(n_8605), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_5__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__u0 ( .ck(ispd_clk), .d(n_8604), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_6__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__u0 ( .ck(ispd_clk), .d(n_8603), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_7__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__u0 ( .ck(ispd_clk), .d(n_8602), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_8__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__u0 ( .ck(ispd_clk), .d(n_8601), .o(wishbone_slave_unit_wishbone_slave_d_incoming_reg_9__Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_del_addr_hit_reg_u0 ( .ck(ispd_clk), .d(n_7723), .o(wishbone_slave_unit_wishbone_slave_del_addr_hit) );
ms00f80 wishbone_slave_unit_wishbone_slave_del_completion_allow_reg_u0 ( .ck(ispd_clk), .d(n_7701), .o(wishbone_slave_unit_wishbone_slave_del_completion_allow) );
ms00f80 wishbone_slave_unit_wishbone_slave_do_del_request_reg_u0 ( .ck(ispd_clk), .d(n_7722), .o(wishbone_slave_unit_wishbone_slave_do_del_request) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_0__u0 ( .ck(ispd_clk), .d(n_7541), .o(wishbone_slave_unit_wishbone_slave_img_hit_0_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_1__u0 ( .ck(ispd_clk), .d(n_7540), .o(wishbone_slave_unit_wishbone_slave_img_hit_1_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_2__u0 ( .ck(ispd_clk), .d(n_5741), .o(wishbone_slave_unit_wishbone_slave_img_hit_2_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_3__u0 ( .ck(ispd_clk), .d(n_5740), .o(wishbone_slave_unit_wishbone_slave_img_hit_3_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_hit_reg_4__u0 ( .ck(ispd_clk), .d(n_5733), .o(wishbone_slave_unit_wishbone_slave_img_hit_4_) );
ms00f80 wishbone_slave_unit_wishbone_slave_img_wallow_reg_u0 ( .ck(ispd_clk), .d(n_7721), .o(wishbone_slave_unit_wishbone_slave_img_wallow) );
ms00f80 wishbone_slave_unit_wishbone_slave_map_reg_u0 ( .ck(ispd_clk), .d(n_7542), .o(wishbone_slave_unit_wishbone_slave_map) );
ms00f80 wishbone_slave_unit_wishbone_slave_mrl_en_reg_u0 ( .ck(ispd_clk), .d(n_7719), .o(wishbone_slave_unit_wishbone_slave_mrl_en_reg_Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_pref_en_reg_u0 ( .ck(ispd_clk), .d(n_7718), .o(wishbone_slave_unit_wishbone_slave_pref_en_reg_Q) );
ms00f80 wishbone_slave_unit_wishbone_slave_wb_conf_hit_reg_u0 ( .ck(ispd_clk), .d(n_5736), .o(wishbone_slave_unit_wishbone_slave_wb_conf_hit) );
ms00f80 wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_u0 ( .ck(ispd_clk), .d(n_8525), .o(wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_Q) );
in01f80 wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_u1 ( .a(wishbone_slave_unit_wishbone_slave_wbw_data_out_sel_reg_reg_Q), .o(n_8831) );
in01f10 TIMEBOOST_cell_0 ( .a(TIMEBOOST_net_0), .o(FE_OCPN1845_n_16427) );
in01f08 TIMEBOOST_cell_1 ( .a(TIMEBOOST_net_1), .o(TIMEBOOST_net_0) );
in01f10 TIMEBOOST_cell_2 ( .a(TIMEBOOST_net_2), .o(n_3252) );
in01f08 TIMEBOOST_cell_3 ( .a(TIMEBOOST_net_3), .o(TIMEBOOST_net_2) );
in01f10 TIMEBOOST_cell_4 ( .a(TIMEBOOST_net_4), .o(FE_OFN1061_n_16720) );
in01f08 TIMEBOOST_cell_5 ( .a(TIMEBOOST_net_5), .o(TIMEBOOST_net_4) );
na03f40 TIMEBOOST_cell_6 ( .a(wishbone_slave_unit_pci_initiator_sm_cur_state_3_), .b(wishbone_slave_unit_pci_initiator_sm_cur_state_2_), .c(n_15680), .o(FE_RN_299_0) );

endmodule
